magic
tech sky130B
magscale 1 2
timestamp 1668096488
<< viali >>
rect 1869 57409 1903 57443
rect 3801 57409 3835 57443
rect 4997 57409 5031 57443
rect 6561 57409 6595 57443
rect 8125 57409 8159 57443
rect 9689 57409 9723 57443
rect 11529 57409 11563 57443
rect 12817 57409 12851 57443
rect 14381 57409 14415 57443
rect 15945 57409 15979 57443
rect 17509 57409 17543 57443
rect 19257 57409 19291 57443
rect 20637 57409 20671 57443
rect 22201 57409 22235 57443
rect 24409 57409 24443 57443
rect 25329 57409 25363 57443
rect 26985 57409 27019 57443
rect 28457 57409 28491 57443
rect 30021 57409 30055 57443
rect 32137 57409 32171 57443
rect 33149 57409 33183 57443
rect 34713 57409 34747 57443
rect 36277 57409 36311 57443
rect 37841 57409 37875 57443
rect 39865 57409 39899 57443
rect 40969 57409 41003 57443
rect 42533 57409 42567 57443
rect 44097 57409 44131 57443
rect 45661 57409 45695 57443
rect 47593 57409 47627 57443
rect 48789 57409 48823 57443
rect 50353 57409 50387 57443
rect 51917 57409 51951 57443
rect 53481 57409 53515 57443
rect 56609 57409 56643 57443
rect 57989 57409 58023 57443
rect 55321 57341 55355 57375
rect 57529 57001 57563 57035
rect 58173 56797 58207 56831
rect 58173 56321 58207 56355
rect 58173 55097 58207 55131
rect 58173 53941 58207 53975
rect 58173 52445 58207 52479
rect 58173 51357 58207 51391
rect 58173 49725 58207 49759
rect 58173 48501 58207 48535
rect 58173 47005 58207 47039
rect 58173 45917 58207 45951
rect 58173 44217 58207 44251
rect 58173 43061 58207 43095
rect 13277 42653 13311 42687
rect 15485 42585 15519 42619
rect 15669 42585 15703 42619
rect 14933 42517 14967 42551
rect 15853 42517 15887 42551
rect 13829 42245 13863 42279
rect 14657 42245 14691 42279
rect 12725 42177 12759 42211
rect 12814 42177 12848 42211
rect 12914 42177 12948 42211
rect 13093 42177 13127 42211
rect 14013 42177 14047 42211
rect 14841 42177 14875 42211
rect 15485 42177 15519 42211
rect 15669 42177 15703 42211
rect 15761 42177 15795 42211
rect 15899 42177 15933 42211
rect 15025 42109 15059 42143
rect 18613 42109 18647 42143
rect 11989 41973 12023 42007
rect 12449 41973 12483 42007
rect 14197 41973 14231 42007
rect 16129 41973 16163 42007
rect 16773 41973 16807 42007
rect 20085 41973 20119 42007
rect 11621 41769 11655 41803
rect 15485 41769 15519 41803
rect 18705 41701 18739 41735
rect 12081 41565 12115 41599
rect 12357 41565 12391 41599
rect 14381 41565 14415 41599
rect 14473 41565 14507 41599
rect 14565 41565 14599 41599
rect 14749 41565 14783 41599
rect 16598 41565 16632 41599
rect 16865 41565 16899 41599
rect 18521 41565 18555 41599
rect 19533 41565 19567 41599
rect 19625 41565 19659 41599
rect 19717 41565 19751 41599
rect 19901 41565 19935 41599
rect 20361 41565 20395 41599
rect 58173 41565 58207 41599
rect 11253 41497 11287 41531
rect 11437 41497 11471 41531
rect 18337 41497 18371 41531
rect 5181 41429 5215 41463
rect 14105 41429 14139 41463
rect 17877 41429 17911 41463
rect 19257 41429 19291 41463
rect 16773 41225 16807 41259
rect 5365 41157 5399 41191
rect 7012 41157 7046 41191
rect 8861 41157 8895 41191
rect 10793 41157 10827 41191
rect 10977 41157 11011 41191
rect 12642 41157 12676 41191
rect 14758 41157 14792 41191
rect 19818 41157 19852 41191
rect 5549 41089 5583 41123
rect 9137 41089 9171 41123
rect 9229 41089 9263 41123
rect 9321 41089 9355 41123
rect 9505 41089 9539 41123
rect 15025 41089 15059 41123
rect 15715 41089 15749 41123
rect 15853 41089 15887 41123
rect 15950 41089 15984 41123
rect 16129 41089 16163 41123
rect 17601 41089 17635 41123
rect 17785 41089 17819 41123
rect 17877 41089 17911 41123
rect 17969 41089 18003 41123
rect 27977 41089 28011 41123
rect 6745 41021 6779 41055
rect 12909 41021 12943 41055
rect 20085 41021 20119 41055
rect 27721 41021 27755 41055
rect 10057 40953 10091 40987
rect 5181 40885 5215 40919
rect 8125 40885 8159 40919
rect 10609 40885 10643 40919
rect 11529 40885 11563 40919
rect 13645 40885 13679 40919
rect 15485 40885 15519 40919
rect 18245 40885 18279 40919
rect 18705 40885 18739 40919
rect 23121 40885 23155 40919
rect 29101 40885 29135 40919
rect 8033 40681 8067 40715
rect 27813 40681 27847 40715
rect 29929 40545 29963 40579
rect 4445 40477 4479 40511
rect 4629 40477 4663 40511
rect 4724 40477 4758 40511
rect 4859 40477 4893 40511
rect 6929 40477 6963 40511
rect 8953 40477 8987 40511
rect 12909 40477 12943 40511
rect 14933 40477 14967 40511
rect 16773 40477 16807 40511
rect 19257 40477 19291 40511
rect 23857 40477 23891 40511
rect 25789 40477 25823 40511
rect 27353 40477 27387 40511
rect 28089 40477 28123 40511
rect 28181 40477 28215 40511
rect 28273 40477 28307 40511
rect 28457 40477 28491 40511
rect 58173 40477 58207 40511
rect 6684 40409 6718 40443
rect 8217 40409 8251 40443
rect 8401 40409 8435 40443
rect 9220 40409 9254 40443
rect 12642 40409 12676 40443
rect 15200 40409 15234 40443
rect 18521 40409 18555 40443
rect 19502 40409 19536 40443
rect 23590 40409 23624 40443
rect 25522 40409 25556 40443
rect 30196 40409 30230 40443
rect 5089 40341 5123 40375
rect 5549 40341 5583 40375
rect 10333 40341 10367 40375
rect 11529 40341 11563 40375
rect 16313 40341 16347 40375
rect 20637 40341 20671 40375
rect 22477 40341 22511 40375
rect 24409 40341 24443 40375
rect 29009 40341 29043 40375
rect 31309 40341 31343 40375
rect 9781 40137 9815 40171
rect 28825 40137 28859 40171
rect 30297 40137 30331 40171
rect 5457 40069 5491 40103
rect 5641 40069 5675 40103
rect 18797 40069 18831 40103
rect 30757 40069 30791 40103
rect 30941 40069 30975 40103
rect 2412 40001 2446 40035
rect 6377 40001 6411 40035
rect 6561 40001 6595 40035
rect 6653 40001 6687 40035
rect 6791 40001 6825 40035
rect 7481 40001 7515 40035
rect 8401 40001 8435 40035
rect 8668 40001 8702 40035
rect 10517 40001 10551 40035
rect 10609 40001 10643 40035
rect 10701 40001 10735 40035
rect 10885 40001 10919 40035
rect 12633 40001 12667 40035
rect 12725 40001 12759 40035
rect 12817 40001 12851 40035
rect 13001 40001 13035 40035
rect 18613 40001 18647 40035
rect 18981 40001 19015 40035
rect 19901 40001 19935 40035
rect 20168 40001 20202 40035
rect 22385 40001 22419 40035
rect 22569 40001 22603 40035
rect 22661 40001 22695 40035
rect 22753 40001 22787 40035
rect 24602 40001 24636 40035
rect 27712 40001 27746 40035
rect 29653 40001 29687 40035
rect 29837 40001 29871 40035
rect 29929 40001 29963 40035
rect 30021 40001 30055 40035
rect 31125 40001 31159 40035
rect 2145 39933 2179 39967
rect 3985 39933 4019 39967
rect 4261 39933 4295 39967
rect 5825 39933 5859 39967
rect 7021 39933 7055 39967
rect 10241 39933 10275 39967
rect 12357 39933 12391 39967
rect 23029 39933 23063 39967
rect 24869 39933 24903 39967
rect 27445 39933 27479 39967
rect 13461 39865 13495 39899
rect 3525 39797 3559 39831
rect 11621 39797 11655 39831
rect 16681 39797 16715 39831
rect 21281 39797 21315 39831
rect 23489 39797 23523 39831
rect 2605 39593 2639 39627
rect 6377 39593 6411 39627
rect 9229 39593 9263 39627
rect 10701 39593 10735 39627
rect 20085 39593 20119 39627
rect 20545 39593 20579 39627
rect 22109 39593 22143 39627
rect 23213 39593 23247 39627
rect 29561 39593 29595 39627
rect 11161 39457 11195 39491
rect 2881 39389 2915 39423
rect 2973 39389 3007 39423
rect 3065 39389 3099 39423
rect 3249 39389 3283 39423
rect 4997 39389 5031 39423
rect 5253 39389 5287 39423
rect 9505 39389 9539 39423
rect 9597 39389 9631 39423
rect 9689 39389 9723 39423
rect 9873 39389 9907 39423
rect 10333 39389 10367 39423
rect 19441 39389 19475 39423
rect 19625 39389 19659 39423
rect 19717 39389 19751 39423
rect 19809 39389 19843 39423
rect 21741 39389 21775 39423
rect 22569 39389 22603 39423
rect 22753 39389 22787 39423
rect 22845 39389 22879 39423
rect 22983 39389 23017 39423
rect 23673 39389 23707 39423
rect 26801 39389 26835 39423
rect 30389 39389 30423 39423
rect 31861 39389 31895 39423
rect 3985 39321 4019 39355
rect 4169 39321 4203 39355
rect 10517 39321 10551 39355
rect 21925 39321 21959 39355
rect 29745 39321 29779 39355
rect 29929 39321 29963 39355
rect 32128 39321 32162 39355
rect 3801 39253 3835 39287
rect 18705 39253 18739 39287
rect 28089 39253 28123 39287
rect 31401 39253 31435 39287
rect 33241 39253 33275 39287
rect 33793 39253 33827 39287
rect 4905 39049 4939 39083
rect 19533 39049 19567 39083
rect 23029 39049 23063 39083
rect 23857 39049 23891 39083
rect 27721 39049 27755 39083
rect 32137 39049 32171 39083
rect 29193 38981 29227 39015
rect 34069 38981 34103 39015
rect 35642 38981 35676 39015
rect 8953 38913 8987 38947
rect 11529 38913 11563 38947
rect 19165 38913 19199 38947
rect 19349 38913 19383 38947
rect 22385 38913 22419 38947
rect 22569 38913 22603 38947
rect 22661 38913 22695 38947
rect 22753 38913 22787 38947
rect 23489 38913 23523 38947
rect 23673 38913 23707 38947
rect 27997 38913 28031 38947
rect 28089 38913 28123 38947
rect 28181 38913 28215 38947
rect 28365 38913 28399 38947
rect 29009 38913 29043 38947
rect 30205 38913 30239 38947
rect 30472 38913 30506 38947
rect 32413 38913 32447 38947
rect 32505 38913 32539 38947
rect 32597 38913 32631 38947
rect 32781 38913 32815 38947
rect 33425 38913 33459 38947
rect 33609 38913 33643 38947
rect 33701 38913 33735 38947
rect 33793 38913 33827 38947
rect 13093 38845 13127 38879
rect 13369 38845 13403 38879
rect 28825 38845 28859 38879
rect 35909 38845 35943 38879
rect 58173 38777 58207 38811
rect 3433 38709 3467 38743
rect 10425 38709 10459 38743
rect 21925 38709 21959 38743
rect 27169 38709 27203 38743
rect 31585 38709 31619 38743
rect 34529 38709 34563 38743
rect 9873 38505 9907 38539
rect 22845 38505 22879 38539
rect 24501 38505 24535 38539
rect 30481 38505 30515 38539
rect 32413 38505 32447 38539
rect 12173 38437 12207 38471
rect 7021 38369 7055 38403
rect 7297 38369 7331 38403
rect 31953 38369 31987 38403
rect 36093 38369 36127 38403
rect 3801 38301 3835 38335
rect 9689 38301 9723 38335
rect 11989 38301 12023 38335
rect 12633 38301 12667 38335
rect 13001 38301 13035 38335
rect 15209 38301 15243 38335
rect 15485 38301 15519 38335
rect 15577 38301 15611 38335
rect 17049 38301 17083 38335
rect 17142 38301 17176 38335
rect 17325 38301 17359 38335
rect 17514 38301 17548 38335
rect 22661 38301 22695 38335
rect 27353 38301 27387 38335
rect 30757 38301 30791 38335
rect 30849 38301 30883 38335
rect 30941 38301 30975 38335
rect 31125 38301 31159 38335
rect 32597 38301 32631 38335
rect 33517 38301 33551 38335
rect 33701 38301 33735 38335
rect 33793 38301 33827 38335
rect 33931 38301 33965 38335
rect 4046 38233 4080 38267
rect 5825 38233 5859 38267
rect 6009 38233 6043 38267
rect 9505 38233 9539 38267
rect 12817 38233 12851 38267
rect 12909 38233 12943 38267
rect 15393 38233 15427 38267
rect 17417 38233 17451 38267
rect 22477 38233 22511 38267
rect 27620 38233 27654 38267
rect 31585 38233 31619 38267
rect 31769 38233 31803 38267
rect 32781 38233 32815 38267
rect 34161 38233 34195 38267
rect 35826 38233 35860 38267
rect 3157 38165 3191 38199
rect 5181 38165 5215 38199
rect 5641 38165 5675 38199
rect 13185 38165 13219 38199
rect 15761 38165 15795 38199
rect 17693 38165 17727 38199
rect 19441 38165 19475 38199
rect 28733 38165 28767 38199
rect 29929 38165 29963 38199
rect 34713 38165 34747 38199
rect 15669 37961 15703 37995
rect 20729 37961 20763 37995
rect 33793 37961 33827 37995
rect 34989 37961 35023 37995
rect 7481 37893 7515 37927
rect 8493 37893 8527 37927
rect 15393 37893 15427 37927
rect 18889 37893 18923 37927
rect 34161 37893 34195 37927
rect 34621 37893 34655 37927
rect 2605 37825 2639 37859
rect 2697 37825 2731 37859
rect 2789 37825 2823 37859
rect 2973 37825 3007 37859
rect 5181 37825 5215 37859
rect 7297 37825 7331 37859
rect 7573 37825 7607 37859
rect 7665 37825 7699 37859
rect 8309 37825 8343 37859
rect 8585 37825 8619 37859
rect 8677 37825 8711 37859
rect 12265 37825 12299 37859
rect 13369 37825 13403 37859
rect 13462 37825 13496 37859
rect 13645 37825 13679 37859
rect 13737 37825 13771 37859
rect 13834 37825 13868 37859
rect 15117 37825 15151 37859
rect 15255 37825 15289 37859
rect 15485 37825 15519 37859
rect 16937 37825 16971 37859
rect 18521 37825 18555 37859
rect 18614 37825 18648 37859
rect 18797 37825 18831 37859
rect 18986 37825 19020 37859
rect 19625 37825 19659 37859
rect 19809 37825 19843 37859
rect 19901 37825 19935 37859
rect 19993 37825 20027 37859
rect 25706 37825 25740 37859
rect 31033 37825 31067 37859
rect 32597 37825 32631 37859
rect 33977 37825 34011 37859
rect 34805 37825 34839 37859
rect 3433 37757 3467 37791
rect 12541 37757 12575 37791
rect 16681 37757 16715 37791
rect 25973 37757 26007 37791
rect 31309 37757 31343 37791
rect 20269 37689 20303 37723
rect 32781 37689 32815 37723
rect 2329 37621 2363 37655
rect 5733 37621 5767 37655
rect 7849 37621 7883 37655
rect 8861 37621 8895 37655
rect 14013 37621 14047 37655
rect 18061 37621 18095 37655
rect 19165 37621 19199 37655
rect 23581 37621 23615 37655
rect 24041 37621 24075 37655
rect 24593 37621 24627 37655
rect 29929 37621 29963 37655
rect 33333 37621 33367 37655
rect 58173 37621 58207 37655
rect 3801 37417 3835 37451
rect 15485 37417 15519 37451
rect 19625 37417 19659 37451
rect 32321 37417 32355 37451
rect 11989 37281 12023 37315
rect 14105 37281 14139 37315
rect 1869 37213 1903 37247
rect 4077 37213 4111 37247
rect 4169 37213 4203 37247
rect 4261 37213 4295 37247
rect 4445 37213 4479 37247
rect 5457 37213 5491 37247
rect 10241 37213 10275 37247
rect 12265 37213 12299 37247
rect 16773 37213 16807 37247
rect 18061 37213 18095 37247
rect 18209 37213 18243 37247
rect 18567 37213 18601 37247
rect 19257 37213 19291 37247
rect 21465 37213 21499 37247
rect 23213 37213 23247 37247
rect 23397 37213 23431 37247
rect 23489 37213 23523 37247
rect 23581 37213 23615 37247
rect 24409 37213 24443 37247
rect 27629 37213 27663 37247
rect 2136 37145 2170 37179
rect 4997 37145 5031 37179
rect 5724 37145 5758 37179
rect 10425 37145 10459 37179
rect 14350 37145 14384 37179
rect 16957 37145 16991 37179
rect 18337 37145 18371 37179
rect 18429 37145 18463 37179
rect 19441 37145 19475 37179
rect 21198 37145 21232 37179
rect 23857 37145 23891 37179
rect 24654 37145 24688 37179
rect 27896 37145 27930 37179
rect 3249 37077 3283 37111
rect 6837 37077 6871 37111
rect 10609 37077 10643 37111
rect 16589 37077 16623 37111
rect 18705 37077 18739 37111
rect 20085 37077 20119 37111
rect 22753 37077 22787 37111
rect 25789 37077 25823 37111
rect 29009 37077 29043 37111
rect 2881 36873 2915 36907
rect 6377 36873 6411 36907
rect 10333 36873 10367 36907
rect 12173 36873 12207 36907
rect 25053 36873 25087 36907
rect 27261 36873 27295 36907
rect 27721 36873 27755 36907
rect 3249 36805 3283 36839
rect 11897 36805 11931 36839
rect 13369 36805 13403 36839
rect 14657 36805 14691 36839
rect 17785 36805 17819 36839
rect 19910 36805 19944 36839
rect 23213 36805 23247 36839
rect 3065 36737 3099 36771
rect 6561 36737 6595 36771
rect 8953 36737 8987 36771
rect 9220 36737 9254 36771
rect 11621 36737 11655 36771
rect 11805 36737 11839 36771
rect 11989 36737 12023 36771
rect 13553 36737 13587 36771
rect 14841 36737 14875 36771
rect 17141 36737 17175 36771
rect 17325 36737 17359 36771
rect 17417 36737 17451 36771
rect 17509 36737 17543 36771
rect 23121 36737 23155 36771
rect 23305 36737 23339 36771
rect 23489 36737 23523 36771
rect 24409 36737 24443 36771
rect 24593 36737 24627 36771
rect 24688 36737 24722 36771
rect 24777 36737 24811 36771
rect 25513 36737 25547 36771
rect 25697 36737 25731 36771
rect 27951 36737 27985 36771
rect 28070 36737 28104 36771
rect 28186 36737 28220 36771
rect 28365 36737 28399 36771
rect 28825 36737 28859 36771
rect 33425 36737 33459 36771
rect 33609 36737 33643 36771
rect 20177 36669 20211 36703
rect 18245 36601 18279 36635
rect 34253 36601 34287 36635
rect 13185 36533 13219 36567
rect 14473 36533 14507 36567
rect 18797 36533 18831 36567
rect 22477 36533 22511 36567
rect 22937 36533 22971 36567
rect 25881 36533 25915 36567
rect 33793 36533 33827 36567
rect 34897 36533 34931 36567
rect 10149 36329 10183 36363
rect 11345 36329 11379 36363
rect 13185 36329 13219 36363
rect 14105 36329 14139 36363
rect 16681 36329 16715 36363
rect 17325 36329 17359 36363
rect 20821 36329 20855 36363
rect 24409 36329 24443 36363
rect 27629 36329 27663 36363
rect 33333 36329 33367 36363
rect 36645 36329 36679 36363
rect 7481 36261 7515 36295
rect 6101 36125 6135 36159
rect 8125 36125 8159 36159
rect 10425 36125 10459 36159
rect 10517 36125 10551 36159
rect 10609 36125 10643 36159
rect 10793 36125 10827 36159
rect 11805 36125 11839 36159
rect 14381 36125 14415 36159
rect 14473 36125 14507 36159
rect 14565 36125 14599 36159
rect 14749 36125 14783 36159
rect 16037 36125 16071 36159
rect 16221 36125 16255 36159
rect 16313 36125 16347 36159
rect 16405 36125 16439 36159
rect 17509 36125 17543 36159
rect 21649 36125 21683 36159
rect 21741 36125 21775 36159
rect 21833 36125 21867 36159
rect 22017 36125 22051 36159
rect 23121 36125 23155 36159
rect 23397 36125 23431 36159
rect 23489 36125 23523 36159
rect 24593 36125 24627 36159
rect 24777 36125 24811 36159
rect 27859 36125 27893 36159
rect 27997 36125 28031 36159
rect 28089 36125 28123 36159
rect 28273 36125 28307 36159
rect 34713 36125 34747 36159
rect 34897 36125 34931 36159
rect 34989 36125 35023 36159
rect 35081 36125 35115 36159
rect 38945 36125 38979 36159
rect 58173 36125 58207 36159
rect 6368 36057 6402 36091
rect 7941 36057 7975 36091
rect 8309 36057 8343 36091
rect 12072 36057 12106 36091
rect 17693 36057 17727 36091
rect 23305 36057 23339 36091
rect 26617 36057 26651 36091
rect 30113 36057 30147 36091
rect 30297 36057 30331 36091
rect 31033 36057 31067 36091
rect 31217 36057 31251 36091
rect 32045 36057 32079 36091
rect 37289 36057 37323 36091
rect 15301 35989 15335 36023
rect 21373 35989 21407 36023
rect 22661 35989 22695 36023
rect 23673 35989 23707 36023
rect 27169 35989 27203 36023
rect 30849 35989 30883 36023
rect 35357 35989 35391 36023
rect 6929 35785 6963 35819
rect 12449 35785 12483 35819
rect 16773 35785 16807 35819
rect 21833 35785 21867 35819
rect 29193 35785 29227 35819
rect 32873 35785 32907 35819
rect 10425 35717 10459 35751
rect 22017 35717 22051 35751
rect 3056 35649 3090 35683
rect 7205 35649 7239 35683
rect 7297 35649 7331 35683
rect 7389 35649 7423 35683
rect 7573 35649 7607 35683
rect 10609 35649 10643 35683
rect 12725 35649 12759 35683
rect 12817 35649 12851 35683
rect 12909 35649 12943 35683
rect 13093 35649 13127 35683
rect 13645 35649 13679 35683
rect 22201 35649 22235 35683
rect 27609 35649 27643 35683
rect 29377 35649 29411 35683
rect 29561 35649 29595 35683
rect 32505 35649 32539 35683
rect 32689 35649 32723 35683
rect 34457 35649 34491 35683
rect 34713 35649 34747 35683
rect 36286 35649 36320 35683
rect 36553 35649 36587 35683
rect 2789 35581 2823 35615
rect 27353 35581 27387 35615
rect 31033 35581 31067 35615
rect 31309 35581 31343 35615
rect 11897 35513 11931 35547
rect 19717 35513 19751 35547
rect 4169 35445 4203 35479
rect 6377 35445 6411 35479
rect 10793 35445 10827 35479
rect 17325 35445 17359 35479
rect 23765 35445 23799 35479
rect 24409 35445 24443 35479
rect 28733 35445 28767 35479
rect 33333 35445 33367 35479
rect 35173 35445 35207 35479
rect 11897 35241 11931 35275
rect 27445 35241 27479 35275
rect 28549 35241 28583 35275
rect 12909 35173 12943 35207
rect 10517 35105 10551 35139
rect 18061 35105 18095 35139
rect 33517 35105 33551 35139
rect 4261 35037 4295 35071
rect 6193 35037 6227 35071
rect 12357 35037 12391 35071
rect 12633 35037 12667 35071
rect 12725 35037 12759 35071
rect 16865 35037 16899 35071
rect 16957 35037 16991 35071
rect 17049 35037 17083 35071
rect 17233 35037 17267 35071
rect 17693 35037 17727 35071
rect 19349 35037 19383 35071
rect 20269 35037 20303 35071
rect 22477 35037 22511 35071
rect 27675 35037 27709 35071
rect 27813 35037 27847 35071
rect 27905 35037 27939 35071
rect 28089 35037 28123 35071
rect 28917 35037 28951 35071
rect 30067 35037 30101 35071
rect 30205 35037 30239 35071
rect 30318 35037 30352 35071
rect 30481 35037 30515 35071
rect 30941 35037 30975 35071
rect 33241 35037 33275 35071
rect 58173 35037 58207 35071
rect 4445 34969 4479 35003
rect 6377 34969 6411 35003
rect 7297 34969 7331 35003
rect 7481 34969 7515 35003
rect 10784 34969 10818 35003
rect 12541 34969 12575 35003
rect 17877 34969 17911 35003
rect 22722 34969 22756 35003
rect 28733 34969 28767 35003
rect 31186 34969 31220 35003
rect 4629 34901 4663 34935
rect 5089 34901 5123 34935
rect 6009 34901 6043 34935
rect 7665 34901 7699 34935
rect 16589 34901 16623 34935
rect 19441 34901 19475 34935
rect 21557 34901 21591 34935
rect 23857 34901 23891 34935
rect 26985 34901 27019 34935
rect 29837 34901 29871 34935
rect 32321 34901 32355 34935
rect 4353 34697 4387 34731
rect 8585 34697 8619 34731
rect 11989 34697 12023 34731
rect 18061 34697 18095 34731
rect 20085 34697 20119 34731
rect 27997 34697 28031 34731
rect 29285 34697 29319 34731
rect 33149 34697 33183 34731
rect 34253 34697 34287 34731
rect 6469 34629 6503 34663
rect 27077 34629 27111 34663
rect 28365 34629 28399 34663
rect 2513 34561 2547 34595
rect 2780 34561 2814 34595
rect 4629 34561 4663 34595
rect 4718 34561 4752 34595
rect 4813 34561 4847 34595
rect 4997 34561 5031 34595
rect 7205 34561 7239 34595
rect 7472 34561 7506 34595
rect 10333 34561 10367 34595
rect 12541 34561 12575 34595
rect 16681 34561 16715 34595
rect 16937 34561 16971 34595
rect 19165 34561 19199 34595
rect 19349 34561 19383 34595
rect 24142 34561 24176 34595
rect 24869 34561 24903 34595
rect 25053 34561 25087 34595
rect 28181 34561 28215 34595
rect 32965 34561 32999 34595
rect 33609 34561 33643 34595
rect 33793 34561 33827 34595
rect 33885 34561 33919 34595
rect 33977 34561 34011 34595
rect 10609 34493 10643 34527
rect 12725 34493 12759 34527
rect 24409 34493 24443 34527
rect 29837 34493 29871 34527
rect 30297 34493 30331 34527
rect 30573 34493 30607 34527
rect 3893 34357 3927 34391
rect 5457 34357 5491 34391
rect 19533 34357 19567 34391
rect 23029 34357 23063 34391
rect 25237 34357 25271 34391
rect 3801 34153 3835 34187
rect 5641 34153 5675 34187
rect 7021 34153 7055 34187
rect 7481 34153 7515 34187
rect 11161 34153 11195 34187
rect 35357 34153 35391 34187
rect 17969 34085 18003 34119
rect 11713 34017 11747 34051
rect 14381 34017 14415 34051
rect 20729 34017 20763 34051
rect 27537 34017 27571 34051
rect 30297 34017 30331 34051
rect 3249 33949 3283 33983
rect 4077 33949 4111 33983
rect 4169 33949 4203 33983
rect 4261 33949 4295 33983
rect 4445 33949 4479 33983
rect 5181 33949 5215 33983
rect 5917 33949 5951 33983
rect 6009 33949 6043 33983
rect 6101 33949 6135 33983
rect 6285 33949 6319 33983
rect 7757 33949 7791 33983
rect 7846 33946 7880 33980
rect 7946 33949 7980 33983
rect 8125 33949 8159 33983
rect 8953 33949 8987 33983
rect 9046 33949 9080 33983
rect 9229 33949 9263 33983
rect 9459 33949 9493 33983
rect 10517 33949 10551 33983
rect 10701 33949 10735 33983
rect 10793 33949 10827 33983
rect 10885 33949 10919 33983
rect 14105 33949 14139 33983
rect 17325 33949 17359 33983
rect 17473 33949 17507 33983
rect 17790 33949 17824 33983
rect 23397 33949 23431 33983
rect 23581 33949 23615 33983
rect 23765 33949 23799 33983
rect 25053 33949 25087 33983
rect 25216 33949 25250 33983
rect 25316 33949 25350 33983
rect 25467 33949 25501 33983
rect 35909 33949 35943 33983
rect 36093 33949 36127 33983
rect 36185 33949 36219 33983
rect 36277 33949 36311 33983
rect 9321 33881 9355 33915
rect 13369 33881 13403 33915
rect 13553 33881 13587 33915
rect 16037 33881 16071 33915
rect 16221 33881 16255 33915
rect 17601 33881 17635 33915
rect 17693 33881 17727 33915
rect 20462 33881 20496 33915
rect 23489 33881 23523 33915
rect 24501 33881 24535 33915
rect 25697 33881 25731 33915
rect 27270 33881 27304 33915
rect 30542 33881 30576 33915
rect 32137 33881 32171 33915
rect 32321 33881 32355 33915
rect 9597 33813 9631 33847
rect 19349 33813 19383 33847
rect 22201 33813 22235 33847
rect 22753 33813 22787 33847
rect 23213 33813 23247 33847
rect 26157 33813 26191 33847
rect 31677 33813 31711 33847
rect 32505 33813 32539 33847
rect 33425 33813 33459 33847
rect 36553 33813 36587 33847
rect 4813 33609 4847 33643
rect 8309 33609 8343 33643
rect 9321 33609 9355 33643
rect 14197 33609 14231 33643
rect 19717 33609 19751 33643
rect 24041 33609 24075 33643
rect 29101 33609 29135 33643
rect 29653 33609 29687 33643
rect 30987 33609 31021 33643
rect 35265 33609 35299 33643
rect 4169 33541 4203 33575
rect 4997 33541 5031 33575
rect 5181 33541 5215 33575
rect 9781 33541 9815 33575
rect 15301 33541 15335 33575
rect 15485 33541 15519 33575
rect 23397 33541 23431 33575
rect 23581 33541 23615 33575
rect 36461 33541 36495 33575
rect 38402 33541 38436 33575
rect 4353 33473 4387 33507
rect 9137 33473 9171 33507
rect 9965 33473 9999 33507
rect 10609 33473 10643 33507
rect 14013 33473 14047 33507
rect 19073 33473 19107 33507
rect 19257 33473 19291 33507
rect 19349 33473 19383 33507
rect 19441 33473 19475 33507
rect 21925 33473 21959 33507
rect 22661 33473 22695 33507
rect 24271 33473 24305 33507
rect 24409 33473 24443 33507
rect 24501 33473 24535 33507
rect 24697 33473 24731 33507
rect 25145 33473 25179 33507
rect 29929 33473 29963 33507
rect 30021 33473 30055 33507
rect 30113 33473 30147 33507
rect 30297 33473 30331 33507
rect 35817 33473 35851 33507
rect 36001 33473 36035 33507
rect 36093 33473 36127 33507
rect 36185 33473 36219 33507
rect 38669 33473 38703 33507
rect 17601 33405 17635 33439
rect 17877 33405 17911 33439
rect 23213 33405 23247 33439
rect 30757 33405 30791 33439
rect 10793 33337 10827 33371
rect 20269 33337 20303 33371
rect 58173 33337 58207 33371
rect 3985 33269 4019 33303
rect 22477 33269 22511 33303
rect 37289 33269 37323 33303
rect 7205 33065 7239 33099
rect 17785 33065 17819 33099
rect 22569 33065 22603 33099
rect 23765 33065 23799 33099
rect 29653 33065 29687 33099
rect 35449 33065 35483 33099
rect 8125 32997 8159 33031
rect 31125 32997 31159 33031
rect 37105 32997 37139 33031
rect 4997 32929 5031 32963
rect 9597 32929 9631 32963
rect 24409 32929 24443 32963
rect 38485 32929 38519 32963
rect 4077 32861 4111 32895
rect 4169 32861 4203 32895
rect 4261 32861 4295 32895
rect 4445 32861 4479 32895
rect 6377 32861 6411 32895
rect 7389 32861 7423 32895
rect 8309 32861 8343 32895
rect 9873 32861 9907 32895
rect 11713 32861 11747 32895
rect 12081 32861 12115 32895
rect 12909 32861 12943 32895
rect 14105 32861 14139 32895
rect 17601 32861 17635 32895
rect 21649 32861 21683 32895
rect 24685 32861 24719 32895
rect 28825 32861 28859 32895
rect 30941 32861 30975 32895
rect 32689 32861 32723 32895
rect 33057 32861 33091 32895
rect 35265 32861 35299 32895
rect 35909 32861 35943 32895
rect 36093 32861 36127 32895
rect 36185 32861 36219 32895
rect 36277 32861 36311 32895
rect 38218 32861 38252 32895
rect 6561 32793 6595 32827
rect 11897 32793 11931 32827
rect 11989 32793 12023 32827
rect 12725 32793 12759 32827
rect 14372 32793 14406 32827
rect 21404 32793 21438 32827
rect 28641 32793 28675 32827
rect 32781 32793 32815 32827
rect 32873 32793 32907 32827
rect 35081 32793 35115 32827
rect 3801 32725 3835 32759
rect 6745 32725 6779 32759
rect 12265 32725 12299 32759
rect 13093 32725 13127 32759
rect 15485 32725 15519 32759
rect 20269 32725 20303 32759
rect 28457 32725 28491 32759
rect 32505 32725 32539 32759
rect 36553 32725 36587 32759
rect 4629 32521 4663 32555
rect 7573 32521 7607 32555
rect 11621 32521 11655 32555
rect 30941 32521 30975 32555
rect 35265 32521 35299 32555
rect 36185 32521 36219 32555
rect 9965 32453 9999 32487
rect 14565 32453 14599 32487
rect 15025 32453 15059 32487
rect 15209 32453 15243 32487
rect 17049 32453 17083 32487
rect 21097 32453 21131 32487
rect 21833 32453 21867 32487
rect 27353 32453 27387 32487
rect 32689 32453 32723 32487
rect 35817 32453 35851 32487
rect 2780 32385 2814 32419
rect 5825 32385 5859 32419
rect 6653 32385 6687 32419
rect 6742 32385 6776 32419
rect 6837 32385 6871 32419
rect 7021 32385 7055 32419
rect 9045 32385 9079 32419
rect 9781 32385 9815 32419
rect 12734 32385 12768 32419
rect 13001 32385 13035 32419
rect 13921 32385 13955 32419
rect 14105 32385 14139 32419
rect 14200 32385 14234 32419
rect 14335 32385 14369 32419
rect 16681 32385 16715 32419
rect 16774 32385 16808 32419
rect 16957 32385 16991 32419
rect 17146 32385 17180 32419
rect 20913 32385 20947 32419
rect 22063 32385 22097 32419
rect 22201 32385 22235 32419
rect 22293 32385 22327 32419
rect 22477 32385 22511 32419
rect 22937 32385 22971 32419
rect 24133 32385 24167 32419
rect 24296 32385 24330 32419
rect 24396 32385 24430 32419
rect 24547 32385 24581 32419
rect 25237 32385 25271 32419
rect 29817 32385 29851 32419
rect 32597 32385 32631 32419
rect 32781 32385 32815 32419
rect 32965 32385 32999 32419
rect 36001 32385 36035 32419
rect 2513 32317 2547 32351
rect 8769 32317 8803 32351
rect 15393 32317 15427 32351
rect 21281 32317 21315 32351
rect 29561 32317 29595 32351
rect 3893 32249 3927 32283
rect 23121 32249 23155 32283
rect 6377 32181 6411 32215
rect 10149 32181 10183 32215
rect 17325 32181 17359 32215
rect 24777 32181 24811 32215
rect 28641 32181 28675 32215
rect 32413 32181 32447 32215
rect 58173 32181 58207 32215
rect 7021 31977 7055 32011
rect 10333 31977 10367 32011
rect 12541 31977 12575 32011
rect 17509 31977 17543 32011
rect 19993 31977 20027 32011
rect 22845 31977 22879 32011
rect 27721 31977 27755 32011
rect 28273 31977 28307 32011
rect 30113 31977 30147 32011
rect 36001 31977 36035 32011
rect 37013 31977 37047 32011
rect 26341 31909 26375 31943
rect 31217 31909 31251 31943
rect 32229 31909 32263 31943
rect 8953 31841 8987 31875
rect 16129 31841 16163 31875
rect 25789 31841 25823 31875
rect 1869 31773 1903 31807
rect 5733 31773 5767 31807
rect 8033 31773 8067 31807
rect 12817 31773 12851 31807
rect 12906 31767 12940 31801
rect 13001 31773 13035 31807
rect 13185 31773 13219 31807
rect 16396 31773 16430 31807
rect 18153 31773 18187 31807
rect 19809 31773 19843 31807
rect 20453 31773 20487 31807
rect 25522 31773 25556 31807
rect 26525 31773 26559 31807
rect 28549 31773 28583 31807
rect 28641 31773 28675 31807
rect 28733 31773 28767 31807
rect 28917 31773 28951 31807
rect 31401 31773 31435 31807
rect 31493 31773 31527 31807
rect 31769 31773 31803 31807
rect 32413 31773 32447 31807
rect 32505 31773 32539 31807
rect 32781 31773 32815 31807
rect 35817 31773 35851 31807
rect 38126 31773 38160 31807
rect 38393 31773 38427 31807
rect 2136 31705 2170 31739
rect 9220 31705 9254 31739
rect 17969 31705 18003 31739
rect 30021 31705 30055 31739
rect 31585 31705 31619 31739
rect 32597 31705 32631 31739
rect 35633 31705 35667 31739
rect 3249 31637 3283 31671
rect 14197 31637 14231 31671
rect 18337 31637 18371 31671
rect 24409 31637 24443 31671
rect 9689 31433 9723 31467
rect 13461 31433 13495 31467
rect 16681 31433 16715 31467
rect 22017 31433 22051 31467
rect 24225 31433 24259 31467
rect 26157 31433 26191 31467
rect 30665 31433 30699 31467
rect 6622 31365 6656 31399
rect 14013 31365 14047 31399
rect 24593 31365 24627 31399
rect 28733 31365 28767 31399
rect 32597 31365 32631 31399
rect 2145 31297 2179 31331
rect 2412 31297 2446 31331
rect 9919 31297 9953 31331
rect 10054 31297 10088 31331
rect 10154 31297 10188 31331
rect 10333 31297 10367 31331
rect 10885 31297 10919 31331
rect 16957 31297 16991 31331
rect 17049 31297 17083 31331
rect 17141 31297 17175 31331
rect 17325 31297 17359 31331
rect 20177 31297 20211 31331
rect 21281 31297 21315 31331
rect 21833 31297 21867 31331
rect 23029 31297 23063 31331
rect 23489 31297 23523 31331
rect 24409 31297 24443 31331
rect 28641 31297 28675 31331
rect 28825 31297 28859 31331
rect 29009 31297 29043 31331
rect 32505 31297 32539 31331
rect 32689 31297 32723 31331
rect 32873 31297 32907 31331
rect 6377 31229 6411 31263
rect 19901 31229 19935 31263
rect 25053 31229 25087 31263
rect 22845 31161 22879 31195
rect 28457 31161 28491 31195
rect 3525 31093 3559 31127
rect 4077 31093 4111 31127
rect 7757 31093 7791 31127
rect 12265 31093 12299 31127
rect 12817 31093 12851 31127
rect 17785 31093 17819 31127
rect 19349 31093 19383 31127
rect 29745 31093 29779 31127
rect 32321 31093 32355 31127
rect 2605 30889 2639 30923
rect 7573 30889 7607 30923
rect 23857 30889 23891 30923
rect 17325 30821 17359 30855
rect 15485 30753 15519 30787
rect 19257 30753 19291 30787
rect 22937 30753 22971 30787
rect 32413 30753 32447 30787
rect 2881 30685 2915 30719
rect 2970 30679 3004 30713
rect 3065 30682 3099 30716
rect 3249 30685 3283 30719
rect 3985 30685 4019 30719
rect 4169 30685 4203 30719
rect 6193 30685 6227 30719
rect 9689 30685 9723 30719
rect 9873 30685 9907 30719
rect 21281 30685 21315 30719
rect 21373 30685 21407 30719
rect 21649 30685 21683 30719
rect 22661 30685 22695 30719
rect 23673 30685 23707 30719
rect 24501 30685 24535 30719
rect 24685 30685 24719 30719
rect 24777 30685 24811 30719
rect 24869 30685 24903 30719
rect 26985 30685 27019 30719
rect 28549 30685 28583 30719
rect 28917 30685 28951 30719
rect 31033 30685 31067 30719
rect 31217 30685 31251 30719
rect 31309 30685 31343 30719
rect 31401 30685 31435 30719
rect 32137 30685 32171 30719
rect 34713 30685 34747 30719
rect 37105 30685 37139 30719
rect 58173 30685 58207 30719
rect 3801 30617 3835 30651
rect 6460 30617 6494 30651
rect 12173 30617 12207 30651
rect 13185 30617 13219 30651
rect 13369 30617 13403 30651
rect 15218 30617 15252 30651
rect 16037 30617 16071 30651
rect 19524 30617 19558 30651
rect 21465 30617 21499 30651
rect 25145 30617 25179 30651
rect 26718 30617 26752 30651
rect 28641 30617 28675 30651
rect 28733 30617 28767 30651
rect 30573 30617 30607 30651
rect 33793 30617 33827 30651
rect 33977 30617 34011 30651
rect 36838 30617 36872 30651
rect 9505 30549 9539 30583
rect 10885 30549 10919 30583
rect 12633 30549 12667 30583
rect 13553 30549 13587 30583
rect 14105 30549 14139 30583
rect 20637 30549 20671 30583
rect 21097 30549 21131 30583
rect 25605 30549 25639 30583
rect 28365 30549 28399 30583
rect 31677 30549 31711 30583
rect 34161 30549 34195 30583
rect 34897 30549 34931 30583
rect 35725 30549 35759 30583
rect 2697 30345 2731 30379
rect 6377 30345 6411 30379
rect 10793 30345 10827 30379
rect 13001 30345 13035 30379
rect 15853 30345 15887 30379
rect 28365 30345 28399 30379
rect 30757 30345 30791 30379
rect 31217 30345 31251 30379
rect 4353 30277 4387 30311
rect 11989 30277 12023 30311
rect 14197 30277 14231 30311
rect 16773 30277 16807 30311
rect 19717 30277 19751 30311
rect 22293 30277 22327 30311
rect 22385 30277 22419 30311
rect 28641 30277 28675 30311
rect 28733 30277 28767 30311
rect 31401 30277 31435 30311
rect 33701 30277 33735 30311
rect 34805 30277 34839 30311
rect 2973 30209 3007 30243
rect 3065 30209 3099 30243
rect 3157 30215 3191 30249
rect 3341 30209 3375 30243
rect 4077 30209 4111 30243
rect 4261 30209 4295 30243
rect 4445 30209 4479 30243
rect 5825 30209 5859 30243
rect 6653 30209 6687 30243
rect 6745 30209 6779 30243
rect 6837 30209 6871 30243
rect 7021 30209 7055 30243
rect 9919 30209 9953 30243
rect 10054 30209 10088 30243
rect 10154 30209 10188 30243
rect 10333 30209 10367 30243
rect 12173 30209 12207 30243
rect 12817 30209 12851 30243
rect 13001 30209 13035 30243
rect 13553 30209 13587 30243
rect 13737 30209 13771 30243
rect 13829 30209 13863 30243
rect 13921 30209 13955 30243
rect 16957 30209 16991 30243
rect 19073 30209 19107 30243
rect 19901 30209 19935 30243
rect 22109 30209 22143 30243
rect 22477 30209 22511 30243
rect 24961 30209 24995 30243
rect 28549 30209 28583 30243
rect 28917 30209 28951 30243
rect 29929 30209 29963 30243
rect 30573 30209 30607 30243
rect 30757 30209 30791 30243
rect 31585 30209 31619 30243
rect 32689 30209 32723 30243
rect 34161 30209 34195 30243
rect 34345 30209 34379 30243
rect 34437 30209 34471 30243
rect 34529 30209 34563 30243
rect 35541 30209 35575 30243
rect 37289 30209 37323 30243
rect 37473 30209 37507 30243
rect 12357 30141 12391 30175
rect 17141 30141 17175 30175
rect 24685 30141 24719 30175
rect 29745 30141 29779 30175
rect 30113 30141 30147 30175
rect 32965 30141 32999 30175
rect 35265 30141 35299 30175
rect 5089 30073 5123 30107
rect 9229 30073 9263 30107
rect 4629 30005 4663 30039
rect 7573 30005 7607 30039
rect 9689 30005 9723 30039
rect 14749 30005 14783 30039
rect 19533 30005 19567 30039
rect 22661 30005 22695 30039
rect 37657 30005 37691 30039
rect 3249 29801 3283 29835
rect 6929 29801 6963 29835
rect 13461 29801 13495 29835
rect 19901 29801 19935 29835
rect 29561 29801 29595 29835
rect 32965 29801 32999 29835
rect 20821 29733 20855 29767
rect 21925 29733 21959 29767
rect 9229 29665 9263 29699
rect 11345 29665 11379 29699
rect 18061 29665 18095 29699
rect 23857 29665 23891 29699
rect 2881 29597 2915 29631
rect 3065 29597 3099 29631
rect 4077 29597 4111 29631
rect 4353 29597 4387 29631
rect 4445 29597 4479 29631
rect 6745 29597 6779 29631
rect 7573 29597 7607 29631
rect 9496 29597 9530 29631
rect 11069 29597 11103 29631
rect 12449 29597 12483 29631
rect 12633 29597 12667 29631
rect 12817 29597 12851 29631
rect 15761 29597 15795 29631
rect 19257 29597 19291 29631
rect 19441 29597 19475 29631
rect 19533 29597 19567 29631
rect 19625 29597 19659 29631
rect 21005 29597 21039 29631
rect 21373 29597 21407 29631
rect 24777 29597 24811 29631
rect 24961 29597 24995 29631
rect 25053 29597 25087 29631
rect 25145 29597 25179 29631
rect 27261 29597 27295 29631
rect 31585 29597 31619 29631
rect 31852 29597 31886 29631
rect 35541 29597 35575 29631
rect 35725 29597 35759 29631
rect 35817 29597 35851 29631
rect 35909 29597 35943 29631
rect 38669 29597 38703 29631
rect 58173 29597 58207 29631
rect 4261 29529 4295 29563
rect 6561 29529 6595 29563
rect 12725 29529 12759 29563
rect 15945 29529 15979 29563
rect 21097 29529 21131 29563
rect 21189 29529 21223 29563
rect 22845 29529 22879 29563
rect 25421 29529 25455 29563
rect 26994 29529 27028 29563
rect 36185 29529 36219 29563
rect 38402 29529 38436 29563
rect 4629 29461 4663 29495
rect 7389 29461 7423 29495
rect 10609 29461 10643 29495
rect 13001 29461 13035 29495
rect 16129 29461 16163 29495
rect 16681 29461 16715 29495
rect 18613 29461 18647 29495
rect 22937 29461 22971 29495
rect 25881 29461 25915 29495
rect 30389 29461 30423 29495
rect 34989 29461 35023 29495
rect 37289 29461 37323 29495
rect 19165 29257 19199 29291
rect 25145 29257 25179 29291
rect 30021 29257 30055 29291
rect 34897 29257 34931 29291
rect 17325 29189 17359 29223
rect 19809 29189 19843 29223
rect 20637 29189 20671 29223
rect 33885 29189 33919 29223
rect 36093 29189 36127 29223
rect 38402 29189 38436 29223
rect 9505 29121 9539 29155
rect 11897 29121 11931 29155
rect 15025 29121 15059 29155
rect 15761 29121 15795 29155
rect 15853 29121 15887 29155
rect 15945 29121 15979 29155
rect 16129 29121 16163 29155
rect 17785 29121 17819 29155
rect 18041 29121 18075 29155
rect 19993 29121 20027 29155
rect 20453 29121 20487 29155
rect 20729 29121 20763 29155
rect 20821 29121 20855 29155
rect 24777 29121 24811 29155
rect 24961 29121 24995 29155
rect 25605 29121 25639 29155
rect 29837 29121 29871 29155
rect 30021 29121 30055 29155
rect 30481 29121 30515 29155
rect 33793 29121 33827 29155
rect 33977 29121 34011 29155
rect 34161 29121 34195 29155
rect 35449 29121 35483 29155
rect 35633 29121 35667 29155
rect 35725 29121 35759 29155
rect 35817 29121 35851 29155
rect 38669 29121 38703 29155
rect 9229 29053 9263 29087
rect 10701 29053 10735 29087
rect 10977 29053 11011 29087
rect 11621 29053 11655 29087
rect 25789 28985 25823 29019
rect 37289 28985 37323 29019
rect 14381 28917 14415 28951
rect 15485 28917 15519 28951
rect 19625 28917 19659 28951
rect 21005 28917 21039 28951
rect 33609 28917 33643 28951
rect 10149 28713 10183 28747
rect 12817 28713 12851 28747
rect 14473 28713 14507 28747
rect 17877 28713 17911 28747
rect 24685 28713 24719 28747
rect 25513 28713 25547 28747
rect 29009 28713 29043 28747
rect 30113 28713 30147 28747
rect 32505 28713 32539 28747
rect 35725 28713 35759 28747
rect 9229 28645 9263 28679
rect 17325 28645 17359 28679
rect 19901 28645 19935 28679
rect 11713 28577 11747 28611
rect 14105 28577 14139 28611
rect 23305 28577 23339 28611
rect 29745 28577 29779 28611
rect 2789 28509 2823 28543
rect 2973 28509 3007 28543
rect 4721 28509 4755 28543
rect 4905 28509 4939 28543
rect 5089 28509 5123 28543
rect 9137 28509 9171 28543
rect 9321 28509 9355 28543
rect 9781 28509 9815 28543
rect 9965 28509 9999 28543
rect 11437 28509 11471 28543
rect 14289 28509 14323 28543
rect 15209 28509 15243 28543
rect 15476 28509 15510 28543
rect 18153 28509 18187 28543
rect 18245 28509 18279 28543
rect 18337 28509 18371 28543
rect 18521 28509 18555 28543
rect 19717 28509 19751 28543
rect 20453 28509 20487 28543
rect 21649 28509 21683 28543
rect 23121 28509 23155 28543
rect 24869 28509 24903 28543
rect 29929 28509 29963 28543
rect 33609 28509 33643 28543
rect 33701 28509 33735 28543
rect 33977 28509 34011 28543
rect 35357 28509 35391 28543
rect 35541 28509 35575 28543
rect 4997 28441 5031 28475
rect 7113 28441 7147 28475
rect 7297 28441 7331 28475
rect 17141 28441 17175 28475
rect 22477 28441 22511 28475
rect 25053 28441 25087 28475
rect 30757 28441 30791 28475
rect 31217 28441 31251 28475
rect 33793 28441 33827 28475
rect 3157 28373 3191 28407
rect 5273 28373 5307 28407
rect 7481 28373 7515 28407
rect 16589 28373 16623 28407
rect 22385 28373 22419 28407
rect 33425 28373 33459 28407
rect 3709 28169 3743 28203
rect 8217 28169 8251 28203
rect 12633 28169 12667 28203
rect 14197 28169 14231 28203
rect 16957 28169 16991 28203
rect 24041 28169 24075 28203
rect 12817 28101 12851 28135
rect 15209 28101 15243 28135
rect 18613 28101 18647 28135
rect 32689 28101 32723 28135
rect 33701 28101 33735 28135
rect 2596 28033 2630 28067
rect 6837 28033 6871 28067
rect 7093 28033 7127 28067
rect 8677 28033 8711 28067
rect 8770 28033 8804 28067
rect 8953 28033 8987 28067
rect 9045 28033 9079 28067
rect 9142 28033 9176 28067
rect 11529 28033 11563 28067
rect 11692 28033 11726 28067
rect 11792 28033 11826 28067
rect 11897 28033 11931 28067
rect 13001 28033 13035 28067
rect 13461 28033 13495 28067
rect 13645 28033 13679 28067
rect 14841 28033 14875 28067
rect 14934 28033 14968 28067
rect 15117 28033 15151 28067
rect 15306 28033 15340 28067
rect 18797 28033 18831 28067
rect 20729 28033 20763 28067
rect 23949 28033 23983 28067
rect 29837 28033 29871 28067
rect 32597 28033 32631 28067
rect 32781 28033 32815 28067
rect 32965 28033 32999 28067
rect 33609 28033 33643 28067
rect 33793 28033 33827 28067
rect 33977 28033 34011 28067
rect 34529 28033 34563 28067
rect 34713 28033 34747 28067
rect 38945 28033 38979 28067
rect 2329 27965 2363 27999
rect 20453 27965 20487 27999
rect 30113 27965 30147 27999
rect 30573 27965 30607 27999
rect 30849 27965 30883 27999
rect 13553 27897 13587 27931
rect 15485 27897 15519 27931
rect 38393 27897 38427 27931
rect 58173 27897 58207 27931
rect 4261 27829 4295 27863
rect 9321 27829 9355 27863
rect 9781 27829 9815 27863
rect 12173 27829 12207 27863
rect 17693 27829 17727 27863
rect 19533 27829 19567 27863
rect 22017 27829 22051 27863
rect 23305 27829 23339 27863
rect 28733 27829 28767 27863
rect 32413 27829 32447 27863
rect 33425 27829 33459 27863
rect 34897 27829 34931 27863
rect 40233 27829 40267 27863
rect 2605 27625 2639 27659
rect 6929 27625 6963 27659
rect 9873 27625 9907 27659
rect 13093 27625 13127 27659
rect 37289 27625 37323 27659
rect 19349 27557 19383 27591
rect 28917 27557 28951 27591
rect 15025 27489 15059 27523
rect 26801 27489 26835 27523
rect 30941 27489 30975 27523
rect 31677 27489 31711 27523
rect 2881 27421 2915 27455
rect 2970 27415 3004 27449
rect 3065 27418 3099 27452
rect 3249 27421 3283 27455
rect 4169 27421 4203 27455
rect 4721 27421 4755 27455
rect 4814 27421 4848 27455
rect 4997 27421 5031 27455
rect 5089 27421 5123 27455
rect 5227 27421 5261 27455
rect 6469 27421 6503 27455
rect 7205 27421 7239 27455
rect 7297 27421 7331 27455
rect 7389 27421 7423 27455
rect 7573 27421 7607 27455
rect 9781 27421 9815 27455
rect 9965 27421 9999 27455
rect 11713 27421 11747 27455
rect 14749 27421 14783 27455
rect 21189 27421 21223 27455
rect 21373 27421 21407 27455
rect 21465 27421 21499 27455
rect 21557 27421 21591 27455
rect 22477 27421 22511 27455
rect 24961 27421 24995 27455
rect 31401 27421 31435 27455
rect 32689 27421 32723 27455
rect 32873 27421 32907 27455
rect 32984 27421 33018 27455
rect 33103 27421 33137 27455
rect 33977 27421 34011 27455
rect 34161 27421 34195 27455
rect 34713 27421 34747 27455
rect 34897 27421 34931 27455
rect 34989 27421 35023 27455
rect 35081 27421 35115 27455
rect 38669 27421 38703 27455
rect 3985 27353 4019 27387
rect 11980 27353 12014 27387
rect 16865 27353 16899 27387
rect 17049 27353 17083 27387
rect 22722 27353 22756 27387
rect 25206 27353 25240 27387
rect 27046 27353 27080 27387
rect 28733 27353 28767 27387
rect 30674 27353 30708 27387
rect 33793 27353 33827 27387
rect 35357 27353 35391 27387
rect 38402 27353 38436 27387
rect 3801 27285 3835 27319
rect 5365 27285 5399 27319
rect 8125 27285 8159 27319
rect 10425 27285 10459 27319
rect 16313 27285 16347 27319
rect 21833 27285 21867 27319
rect 23857 27285 23891 27319
rect 24409 27285 24443 27319
rect 26341 27285 26375 27319
rect 28181 27285 28215 27319
rect 29561 27285 29595 27319
rect 33333 27285 33367 27319
rect 4353 27081 4387 27115
rect 15485 27081 15519 27115
rect 17325 27081 17359 27115
rect 24869 27081 24903 27115
rect 25973 27081 26007 27115
rect 30665 27081 30699 27115
rect 32505 27081 32539 27115
rect 34529 27081 34563 27115
rect 35081 27081 35115 27115
rect 5181 27013 5215 27047
rect 7021 27013 7055 27047
rect 7113 27013 7147 27047
rect 13093 27013 13127 27047
rect 14841 27013 14875 27047
rect 22262 27013 22296 27047
rect 3433 26945 3467 26979
rect 3522 26951 3556 26985
rect 3617 26948 3651 26982
rect 3801 26945 3835 26979
rect 4813 26945 4847 26979
rect 4906 26945 4940 26979
rect 5089 26945 5123 26979
rect 5278 26945 5312 26979
rect 6745 26945 6779 26979
rect 6838 26945 6872 26979
rect 7251 26945 7285 26979
rect 10701 26945 10735 26979
rect 12081 26945 12115 26979
rect 15945 26945 15979 26979
rect 16129 26945 16163 26979
rect 17141 26945 17175 26979
rect 18981 26945 19015 26979
rect 19165 26945 19199 26979
rect 20085 26945 20119 26979
rect 24225 26945 24259 26979
rect 24409 26945 24443 26979
rect 24504 26945 24538 26979
rect 24593 26945 24627 26979
rect 25329 26945 25363 26979
rect 25513 26945 25547 26979
rect 25605 26945 25639 26979
rect 25697 26945 25731 26979
rect 26985 26945 27019 26979
rect 29653 26945 29687 26979
rect 33149 26945 33183 26979
rect 33416 26945 33450 26979
rect 10977 26877 11011 26911
rect 11805 26877 11839 26911
rect 16957 26877 16991 26911
rect 17785 26877 17819 26911
rect 19809 26877 19843 26911
rect 22017 26877 22051 26911
rect 29377 26877 29411 26911
rect 31217 26877 31251 26911
rect 2697 26741 2731 26775
rect 3157 26741 3191 26775
rect 5457 26741 5491 26775
rect 7389 26741 7423 26775
rect 16037 26741 16071 26775
rect 19349 26741 19383 26775
rect 23397 26741 23431 26775
rect 28273 26741 28307 26775
rect 28825 26741 28859 26775
rect 58173 26741 58207 26775
rect 6285 26537 6319 26571
rect 10885 26537 10919 26571
rect 12909 26537 12943 26571
rect 23765 26537 23799 26571
rect 25881 26537 25915 26571
rect 31677 26537 31711 26571
rect 32597 26537 32631 26571
rect 2881 26469 2915 26503
rect 7941 26469 7975 26503
rect 11897 26469 11931 26503
rect 20361 26469 20395 26503
rect 24777 26469 24811 26503
rect 14381 26401 14415 26435
rect 16405 26401 16439 26435
rect 18245 26401 18279 26435
rect 37841 26401 37875 26435
rect 3065 26333 3099 26367
rect 3249 26333 3283 26367
rect 4077 26333 4111 26367
rect 4166 26330 4200 26364
rect 4266 26333 4300 26367
rect 4445 26333 4479 26367
rect 5917 26333 5951 26367
rect 6101 26333 6135 26367
rect 7021 26333 7055 26367
rect 7126 26333 7160 26367
rect 7226 26327 7260 26361
rect 7389 26333 7423 26367
rect 10793 26333 10827 26367
rect 11713 26333 11747 26367
rect 14105 26333 14139 26367
rect 16129 26333 16163 26367
rect 17141 26333 17175 26367
rect 18521 26333 18555 26367
rect 19533 26333 19567 26367
rect 19625 26333 19659 26367
rect 19717 26333 19751 26367
rect 19901 26333 19935 26367
rect 23213 26333 23247 26367
rect 25237 26333 25271 26367
rect 30389 26333 30423 26367
rect 38485 26333 38519 26367
rect 3801 26265 3835 26299
rect 5365 26265 5399 26299
rect 6745 26265 6779 26299
rect 16957 26265 16991 26299
rect 21649 26265 21683 26299
rect 24409 26265 24443 26299
rect 24593 26265 24627 26299
rect 26065 26265 26099 26299
rect 26249 26265 26283 26299
rect 37574 26265 37608 26299
rect 38669 26265 38703 26299
rect 19257 26197 19291 26231
rect 29653 26197 29687 26231
rect 36461 26197 36495 26231
rect 38301 26197 38335 26231
rect 3985 25993 4019 26027
rect 5273 25993 5307 26027
rect 6377 25993 6411 26027
rect 14197 25993 14231 26027
rect 18153 25993 18187 26027
rect 21189 25993 21223 26027
rect 22477 25993 22511 26027
rect 24317 25993 24351 26027
rect 30297 25993 30331 26027
rect 37289 25993 37323 26027
rect 2872 25925 2906 25959
rect 4813 25925 4847 25959
rect 7490 25925 7524 25959
rect 13461 25925 13495 25959
rect 14657 25925 14691 25959
rect 15485 25925 15519 25959
rect 19266 25925 19300 25959
rect 23581 25925 23615 25959
rect 24501 25925 24535 25959
rect 25789 25925 25823 25959
rect 40754 25925 40788 25959
rect 2605 25857 2639 25891
rect 9505 25857 9539 25891
rect 9689 25857 9723 25891
rect 12541 25857 12575 25891
rect 13645 25857 13679 25891
rect 14841 25857 14875 25891
rect 17141 25857 17175 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22109 25857 22143 25891
rect 22201 25857 22235 25891
rect 23351 25857 23385 25891
rect 23489 25857 23523 25891
rect 23764 25857 23798 25891
rect 23857 25857 23891 25891
rect 24685 25857 24719 25891
rect 25973 25857 26007 25891
rect 28558 25857 28592 25891
rect 29653 25857 29687 25891
rect 29837 25857 29871 25891
rect 29932 25857 29966 25891
rect 30021 25857 30055 25891
rect 36645 25857 36679 25891
rect 37545 25857 37579 25891
rect 37654 25857 37688 25891
rect 37749 25857 37783 25891
rect 37933 25857 37967 25891
rect 39782 25857 39816 25891
rect 40049 25857 40083 25891
rect 40509 25857 40543 25891
rect 7757 25789 7791 25823
rect 12817 25789 12851 25823
rect 19533 25789 19567 25823
rect 25605 25789 25639 25823
rect 28825 25789 28859 25823
rect 10977 25721 11011 25755
rect 31309 25721 31343 25755
rect 9873 25653 9907 25687
rect 13277 25653 13311 25687
rect 15577 25653 15611 25687
rect 16957 25653 16991 25687
rect 23213 25653 23247 25687
rect 27445 25653 27479 25687
rect 30757 25653 30791 25687
rect 38669 25653 38703 25687
rect 41889 25653 41923 25687
rect 9045 25449 9079 25483
rect 18521 25449 18555 25483
rect 29009 25449 29043 25483
rect 36829 25449 36863 25483
rect 38577 25449 38611 25483
rect 10701 25381 10735 25415
rect 16773 25381 16807 25415
rect 12173 25313 12207 25347
rect 18613 25313 18647 25347
rect 19257 25313 19291 25347
rect 27261 25313 27295 25347
rect 7205 25245 7239 25279
rect 7665 25245 7699 25279
rect 9827 25245 9861 25279
rect 9962 25242 9996 25276
rect 10062 25245 10096 25279
rect 10241 25245 10275 25279
rect 14841 25245 14875 25279
rect 18705 25245 18739 25279
rect 23116 25245 23150 25279
rect 23213 25245 23247 25279
rect 23488 25245 23522 25279
rect 23581 25245 23615 25279
rect 24777 25245 24811 25279
rect 24961 25245 24995 25279
rect 25053 25245 25087 25279
rect 25191 25245 25225 25279
rect 28641 25245 28675 25279
rect 29837 25245 29871 25279
rect 30021 25245 30055 25279
rect 30113 25245 30147 25279
rect 30205 25245 30239 25279
rect 32321 25245 32355 25279
rect 36461 25245 36495 25279
rect 37473 25245 37507 25279
rect 37933 25245 37967 25279
rect 38112 25242 38146 25276
rect 38209 25245 38243 25279
rect 38321 25245 38355 25279
rect 58173 25245 58207 25279
rect 5549 25177 5583 25211
rect 12440 25177 12474 25211
rect 15086 25177 15120 25211
rect 19524 25177 19558 25211
rect 23305 25177 23339 25211
rect 25421 25177 25455 25211
rect 26994 25177 27028 25211
rect 28825 25177 28859 25211
rect 30481 25177 30515 25211
rect 32054 25177 32088 25211
rect 36645 25177 36679 25211
rect 9597 25109 9631 25143
rect 13553 25109 13587 25143
rect 14289 25109 14323 25143
rect 16221 25109 16255 25143
rect 18337 25109 18371 25143
rect 20637 25109 20671 25143
rect 22937 25109 22971 25143
rect 25881 25109 25915 25143
rect 30941 25109 30975 25143
rect 2605 24905 2639 24939
rect 12633 24905 12667 24939
rect 14749 24905 14783 24939
rect 19533 24905 19567 24939
rect 25329 24905 25363 24939
rect 27629 24905 27663 24939
rect 29745 24905 29779 24939
rect 39405 24905 39439 24939
rect 8760 24837 8794 24871
rect 20177 24837 20211 24871
rect 23489 24837 23523 24871
rect 25513 24837 25547 24871
rect 26433 24837 26467 24871
rect 3718 24769 3752 24803
rect 3985 24769 4019 24803
rect 10609 24769 10643 24803
rect 10698 24772 10732 24806
rect 10798 24769 10832 24803
rect 10977 24769 11011 24803
rect 12909 24769 12943 24803
rect 13001 24769 13035 24803
rect 13093 24769 13127 24803
rect 13277 24769 13311 24803
rect 15025 24769 15059 24803
rect 15117 24769 15151 24803
rect 15209 24769 15243 24803
rect 15393 24769 15427 24803
rect 16957 24769 16991 24803
rect 18889 24769 18923 24803
rect 19052 24769 19086 24803
rect 19168 24769 19202 24803
rect 19303 24769 19337 24803
rect 20361 24769 20395 24803
rect 23300 24769 23334 24803
rect 23397 24769 23431 24803
rect 23617 24769 23651 24803
rect 23765 24769 23799 24803
rect 24593 24769 24627 24803
rect 25697 24769 25731 24803
rect 27859 24769 27893 24803
rect 27994 24769 28028 24803
rect 28094 24769 28128 24803
rect 28273 24769 28307 24803
rect 29377 24769 29411 24803
rect 29561 24769 29595 24803
rect 31318 24769 31352 24803
rect 31585 24769 31619 24803
rect 34998 24769 35032 24803
rect 37933 24769 37967 24803
rect 38096 24775 38130 24809
rect 38196 24775 38230 24809
rect 38347 24769 38381 24803
rect 39037 24769 39071 24803
rect 39221 24769 39255 24803
rect 8493 24701 8527 24735
rect 35265 24701 35299 24735
rect 12081 24633 12115 24667
rect 38577 24633 38611 24667
rect 6653 24565 6687 24599
rect 9873 24565 9907 24599
rect 10333 24565 10367 24599
rect 11529 24565 11563 24599
rect 14197 24565 14231 24599
rect 16129 24565 16163 24599
rect 16773 24565 16807 24599
rect 19993 24565 20027 24599
rect 23121 24565 23155 24599
rect 27169 24565 27203 24599
rect 28825 24565 28859 24599
rect 30205 24565 30239 24599
rect 33885 24565 33919 24599
rect 37473 24565 37507 24599
rect 5825 24361 5859 24395
rect 15209 24361 15243 24395
rect 16129 24361 16163 24395
rect 21465 24361 21499 24395
rect 28089 24361 28123 24395
rect 29561 24361 29595 24395
rect 30757 24361 30791 24395
rect 31309 24361 31343 24395
rect 33609 24361 33643 24395
rect 36553 24361 36587 24395
rect 14197 24293 14231 24327
rect 19717 24293 19751 24327
rect 7021 24225 7055 24259
rect 10057 24225 10091 24259
rect 27261 24225 27295 24259
rect 32505 24225 32539 24259
rect 6469 24157 6503 24191
rect 7288 24157 7322 24191
rect 12061 24157 12095 24191
rect 12170 24151 12204 24185
rect 12265 24157 12299 24191
rect 12449 24157 12483 24191
rect 13461 24157 13495 24191
rect 15393 24157 15427 24191
rect 17417 24157 17451 24191
rect 17601 24157 17635 24191
rect 17693 24157 17727 24191
rect 22707 24157 22741 24191
rect 23065 24157 23099 24191
rect 23213 24157 23247 24191
rect 27905 24157 27939 24191
rect 30113 24157 30147 24191
rect 30297 24157 30331 24191
rect 30389 24157 30423 24191
rect 30481 24157 30515 24191
rect 32965 24157 32999 24191
rect 33149 24157 33183 24191
rect 33241 24157 33275 24191
rect 33333 24157 33367 24191
rect 38761 24157 38795 24191
rect 58173 24157 58207 24191
rect 9689 24089 9723 24123
rect 9873 24089 9907 24123
rect 10977 24089 11011 24123
rect 11161 24089 11195 24123
rect 11345 24089 11379 24123
rect 13277 24089 13311 24123
rect 15577 24089 15611 24123
rect 22845 24089 22879 24123
rect 22937 24089 22971 24123
rect 26525 24089 26559 24123
rect 27077 24089 27111 24123
rect 27721 24089 27755 24123
rect 6285 24021 6319 24055
rect 8401 24021 8435 24055
rect 11805 24021 11839 24055
rect 14749 24021 14783 24055
rect 16957 24021 16991 24055
rect 22569 24021 22603 24055
rect 37473 24021 37507 24055
rect 11529 23817 11563 23851
rect 17325 23817 17359 23851
rect 19809 23817 19843 23851
rect 25145 23817 25179 23851
rect 30021 23817 30055 23851
rect 39313 23817 39347 23851
rect 2697 23749 2731 23783
rect 3525 23749 3559 23783
rect 7757 23749 7791 23783
rect 9965 23749 9999 23783
rect 12642 23749 12676 23783
rect 13369 23749 13403 23783
rect 14381 23749 14415 23783
rect 15485 23749 15519 23783
rect 19901 23749 19935 23783
rect 21833 23749 21867 23783
rect 22017 23749 22051 23783
rect 25789 23749 25823 23783
rect 27721 23749 27755 23783
rect 29837 23749 29871 23783
rect 36553 23749 36587 23783
rect 2513 23681 2547 23715
rect 3341 23681 3375 23715
rect 5825 23681 5859 23715
rect 7205 23681 7239 23715
rect 10149 23681 10183 23715
rect 10333 23681 10367 23715
rect 12909 23681 12943 23715
rect 14289 23681 14323 23715
rect 14473 23681 14507 23715
rect 14657 23681 14691 23715
rect 15209 23681 15243 23715
rect 15393 23681 15427 23715
rect 15577 23681 15611 23715
rect 18153 23681 18187 23715
rect 20637 23681 20671 23715
rect 20821 23681 20855 23715
rect 20913 23681 20947 23715
rect 21005 23681 21039 23715
rect 22201 23681 22235 23715
rect 27537 23681 27571 23715
rect 29653 23681 29687 23715
rect 33986 23681 34020 23715
rect 36369 23681 36403 23715
rect 38200 23681 38234 23715
rect 5549 23613 5583 23647
rect 6929 23613 6963 23647
rect 10793 23613 10827 23647
rect 34253 23613 34287 23647
rect 37933 23613 37967 23647
rect 2329 23545 2363 23579
rect 16773 23545 16807 23579
rect 21281 23545 21315 23579
rect 25973 23545 26007 23579
rect 3157 23477 3191 23511
rect 14105 23477 14139 23511
rect 15761 23477 15795 23511
rect 18337 23477 18371 23511
rect 27905 23477 27939 23511
rect 32873 23477 32907 23511
rect 36737 23477 36771 23511
rect 12633 23273 12667 23307
rect 15025 23273 15059 23307
rect 24501 23273 24535 23307
rect 33517 23273 33551 23307
rect 38117 23273 38151 23307
rect 3893 23205 3927 23239
rect 32689 23205 32723 23239
rect 5641 23137 5675 23171
rect 17141 23137 17175 23171
rect 18153 23137 18187 23171
rect 19809 23137 19843 23171
rect 28733 23137 28767 23171
rect 36093 23137 36127 23171
rect 2881 23069 2915 23103
rect 2973 23069 3007 23103
rect 3065 23066 3099 23100
rect 3249 23069 3283 23103
rect 4537 23069 4571 23103
rect 4721 23069 4755 23103
rect 4813 23069 4847 23103
rect 4905 23069 4939 23103
rect 7849 23069 7883 23103
rect 11529 23069 11563 23103
rect 11621 23069 11655 23103
rect 11897 23069 11931 23103
rect 15485 23069 15519 23103
rect 15633 23069 15667 23103
rect 15761 23069 15795 23103
rect 15991 23069 16025 23103
rect 17417 23069 17451 23103
rect 17877 23069 17911 23103
rect 20085 23069 20119 23103
rect 22845 23069 22879 23103
rect 32045 23069 32079 23103
rect 32229 23069 32263 23103
rect 32321 23069 32355 23103
rect 32413 23069 32447 23103
rect 33333 23069 33367 23103
rect 37473 23069 37507 23103
rect 37657 23069 37691 23103
rect 37749 23069 37783 23103
rect 37841 23069 37875 23103
rect 5181 23001 5215 23035
rect 5886 23001 5920 23035
rect 7481 23001 7515 23035
rect 7665 23001 7699 23035
rect 11713 23001 11747 23035
rect 15853 23001 15887 23035
rect 21097 23001 21131 23035
rect 28466 23001 28500 23035
rect 33149 23001 33183 23035
rect 35826 23001 35860 23035
rect 2605 22933 2639 22967
rect 7021 22933 7055 22967
rect 11345 22933 11379 22967
rect 16129 22933 16163 22967
rect 27353 22933 27387 22967
rect 31493 22933 31527 22967
rect 34713 22933 34747 22967
rect 37013 22933 37047 22967
rect 20269 22729 20303 22763
rect 27721 22729 27755 22763
rect 29469 22729 29503 22763
rect 32137 22729 32171 22763
rect 33701 22729 33735 22763
rect 9597 22661 9631 22695
rect 9689 22661 9723 22695
rect 20545 22661 20579 22695
rect 22100 22661 22134 22695
rect 25973 22661 26007 22695
rect 30113 22661 30147 22695
rect 32321 22661 32355 22695
rect 32505 22661 32539 22695
rect 3157 22593 3191 22627
rect 3246 22593 3280 22627
rect 3341 22593 3375 22627
rect 3525 22593 3559 22627
rect 3985 22593 4019 22627
rect 4148 22593 4182 22627
rect 4264 22596 4298 22630
rect 4353 22593 4387 22627
rect 5457 22593 5491 22627
rect 5641 22593 5675 22627
rect 6377 22593 6411 22627
rect 6561 22593 6595 22627
rect 6656 22593 6690 22627
rect 6791 22593 6825 22627
rect 9413 22593 9447 22627
rect 9781 22593 9815 22627
rect 19625 22593 19659 22627
rect 20448 22593 20482 22627
rect 20637 22593 20671 22627
rect 20765 22593 20799 22627
rect 20913 22593 20947 22627
rect 21833 22593 21867 22627
rect 23857 22593 23891 22627
rect 24685 22593 24719 22627
rect 24869 22593 24903 22627
rect 24964 22593 24998 22627
rect 25053 22593 25087 22627
rect 26157 22593 26191 22627
rect 27997 22593 28031 22627
rect 28089 22593 28123 22627
rect 28181 22593 28215 22627
rect 28365 22593 28399 22627
rect 33057 22593 33091 22627
rect 33241 22593 33275 22627
rect 33333 22593 33367 22627
rect 33425 22593 33459 22627
rect 38669 22593 38703 22627
rect 38936 22593 38970 22627
rect 5825 22525 5859 22559
rect 19533 22525 19567 22559
rect 2421 22457 2455 22491
rect 25789 22457 25823 22491
rect 30297 22457 30331 22491
rect 40509 22457 40543 22491
rect 58173 22457 58207 22491
rect 2881 22389 2915 22423
rect 4629 22389 4663 22423
rect 7021 22389 7055 22423
rect 7573 22389 7607 22423
rect 9965 22389 9999 22423
rect 16037 22389 16071 22423
rect 19257 22389 19291 22423
rect 19625 22389 19659 22423
rect 23213 22389 23247 22423
rect 23765 22389 23799 22423
rect 25329 22389 25363 22423
rect 27261 22389 27295 22423
rect 40049 22389 40083 22423
rect 4169 22185 4203 22219
rect 5365 22185 5399 22219
rect 7481 22185 7515 22219
rect 15669 22185 15703 22219
rect 18521 22185 18555 22219
rect 19441 22185 19475 22219
rect 29745 22185 29779 22219
rect 39865 22185 39899 22219
rect 41337 22185 41371 22219
rect 26341 22117 26375 22151
rect 29561 22117 29595 22151
rect 14289 22049 14323 22083
rect 19533 22049 19567 22083
rect 24409 22049 24443 22083
rect 30757 22049 30791 22083
rect 32965 22049 32999 22083
rect 38209 22049 38243 22083
rect 2982 21981 3016 22015
rect 3249 21981 3283 22015
rect 6101 21981 6135 22015
rect 9229 21981 9263 22015
rect 9413 21981 9447 22015
rect 9597 21981 9631 22015
rect 17693 21981 17727 22015
rect 18613 21981 18647 22015
rect 18705 21981 18739 22015
rect 19625 21981 19659 22015
rect 24961 21981 24995 22015
rect 29745 21981 29779 22015
rect 29837 21981 29871 22015
rect 30021 21981 30055 22015
rect 30573 21981 30607 22015
rect 31217 21981 31251 22015
rect 32781 21981 32815 22015
rect 35817 21981 35851 22015
rect 36185 21981 36219 22015
rect 38945 21981 38979 22015
rect 39034 21981 39068 22015
rect 39150 21981 39184 22015
rect 39313 21981 39347 22015
rect 40141 21981 40175 22015
rect 40233 21981 40267 22015
rect 40325 21981 40359 22015
rect 40509 21981 40543 22015
rect 3801 21913 3835 21947
rect 3985 21913 4019 21947
rect 6368 21913 6402 21947
rect 9505 21913 9539 21947
rect 14556 21913 14590 21947
rect 16129 21913 16163 21947
rect 21833 21913 21867 21947
rect 22661 21913 22695 21947
rect 25228 21913 25262 21947
rect 27353 21913 27387 21947
rect 32597 21913 32631 21947
rect 35909 21913 35943 21947
rect 36001 21913 36035 21947
rect 40969 21913 41003 21947
rect 41153 21913 41187 21947
rect 1869 21845 1903 21879
rect 4721 21845 4755 21879
rect 9781 21845 9815 21879
rect 18337 21845 18371 21879
rect 19257 21845 19291 21879
rect 20085 21845 20119 21879
rect 20913 21845 20947 21879
rect 22569 21845 22603 21879
rect 23581 21845 23615 21879
rect 26801 21845 26835 21879
rect 33517 21845 33551 21879
rect 35633 21845 35667 21879
rect 37197 21845 37231 21879
rect 38669 21845 38703 21879
rect 3801 21641 3835 21675
rect 5641 21641 5675 21675
rect 14565 21641 14599 21675
rect 21189 21641 21223 21675
rect 25513 21641 25547 21675
rect 27353 21641 27387 21675
rect 29377 21641 29411 21675
rect 32137 21641 32171 21675
rect 4528 21573 4562 21607
rect 6745 21573 6779 21607
rect 7113 21573 7147 21607
rect 12725 21573 12759 21607
rect 12909 21573 12943 21607
rect 17325 21573 17359 21607
rect 25973 21573 26007 21607
rect 26341 21573 26375 21607
rect 28089 21573 28123 21607
rect 28181 21573 28215 21607
rect 29837 21573 29871 21607
rect 30849 21573 30883 21607
rect 30941 21573 30975 21607
rect 32597 21573 32631 21607
rect 35624 21573 35658 21607
rect 37289 21573 37323 21607
rect 39006 21573 39040 21607
rect 2421 21505 2455 21539
rect 2688 21505 2722 21539
rect 4261 21505 4295 21539
rect 8208 21505 8242 21539
rect 13921 21505 13955 21539
rect 14105 21505 14139 21539
rect 14197 21505 14231 21539
rect 14335 21505 14369 21539
rect 15209 21505 15243 21539
rect 15393 21505 15427 21539
rect 16037 21505 16071 21539
rect 17877 21505 17911 21539
rect 18040 21505 18074 21539
rect 18153 21505 18187 21539
rect 18245 21505 18279 21539
rect 18981 21505 19015 21539
rect 19165 21505 19199 21539
rect 22477 21505 22511 21539
rect 22569 21505 22603 21539
rect 22661 21505 22695 21539
rect 22845 21505 22879 21539
rect 24869 21505 24903 21539
rect 25053 21505 25087 21539
rect 25145 21505 25179 21539
rect 25237 21505 25271 21539
rect 26157 21505 26191 21539
rect 27261 21505 27295 21539
rect 27905 21505 27939 21539
rect 28273 21505 28307 21539
rect 29561 21505 29595 21539
rect 30665 21505 30699 21539
rect 31033 21505 31067 21539
rect 32321 21505 32355 21539
rect 37565 21505 37599 21539
rect 37657 21505 37691 21539
rect 37749 21505 37783 21539
rect 37933 21505 37967 21539
rect 7941 21437 7975 21471
rect 15025 21437 15059 21471
rect 19809 21437 19843 21471
rect 20085 21437 20119 21471
rect 23581 21437 23615 21471
rect 23857 21437 23891 21471
rect 29653 21437 29687 21471
rect 32413 21437 32447 21471
rect 35357 21437 35391 21471
rect 38761 21437 38795 21471
rect 11621 21369 11655 21403
rect 19349 21369 19383 21403
rect 31217 21369 31251 21403
rect 9321 21301 9355 21335
rect 12173 21301 12207 21335
rect 13369 21301 13403 21335
rect 15853 21301 15887 21335
rect 16773 21301 16807 21335
rect 18521 21301 18555 21335
rect 22201 21301 22235 21335
rect 28457 21301 28491 21335
rect 29561 21301 29595 21335
rect 32413 21301 32447 21335
rect 36737 21301 36771 21335
rect 40141 21301 40175 21335
rect 58173 21301 58207 21335
rect 10149 21097 10183 21131
rect 15393 21097 15427 21131
rect 17601 21097 17635 21131
rect 25145 21097 25179 21131
rect 28365 21097 28399 21131
rect 31309 21097 31343 21131
rect 32137 21097 32171 21131
rect 35633 21097 35667 21131
rect 36737 21097 36771 21131
rect 40233 21097 40267 21131
rect 24593 21029 24627 21063
rect 26985 21029 27019 21063
rect 31953 21029 31987 21063
rect 11253 20961 11287 20995
rect 14381 20961 14415 20995
rect 19257 20961 19291 20995
rect 9689 20893 9723 20927
rect 10379 20893 10413 20927
rect 10517 20893 10551 20927
rect 10609 20893 10643 20927
rect 10793 20893 10827 20927
rect 11437 20893 11471 20927
rect 14105 20893 14139 20927
rect 15577 20893 15611 20927
rect 15761 20893 15795 20927
rect 18061 20893 18095 20927
rect 18245 20893 18279 20927
rect 18337 20893 18371 20927
rect 18429 20893 18463 20927
rect 21281 20893 21315 20927
rect 21465 20893 21499 20927
rect 21557 20893 21591 20927
rect 21649 20893 21683 20927
rect 22385 20893 22419 20927
rect 22641 20893 22675 20927
rect 24409 20893 24443 20927
rect 25605 20893 25639 20927
rect 27813 20893 27847 20927
rect 28089 20893 28123 20927
rect 28181 20893 28215 20927
rect 29745 20893 29779 20927
rect 30113 20893 30147 20927
rect 30757 20893 30791 20927
rect 30941 20893 30975 20927
rect 31125 20893 31159 20927
rect 32137 20893 32171 20927
rect 32229 20893 32263 20927
rect 35817 20893 35851 20927
rect 35909 20893 35943 20927
rect 36001 20893 36035 20927
rect 36185 20893 36219 20927
rect 40049 20893 40083 20927
rect 5733 20825 5767 20859
rect 7481 20825 7515 20859
rect 12265 20825 12299 20859
rect 12817 20825 12851 20859
rect 17233 20825 17267 20859
rect 17417 20825 17451 20859
rect 18705 20825 18739 20859
rect 19502 20825 19536 20859
rect 25850 20825 25884 20859
rect 27997 20825 28031 20859
rect 29929 20825 29963 20859
rect 30021 20825 30055 20859
rect 31033 20825 31067 20859
rect 32413 20825 32447 20859
rect 36921 20825 36955 20859
rect 37105 20825 37139 20859
rect 39865 20825 39899 20859
rect 7941 20757 7975 20791
rect 12909 20757 12943 20791
rect 20637 20757 20671 20791
rect 21925 20757 21959 20791
rect 23765 20757 23799 20791
rect 30297 20757 30331 20791
rect 7665 20553 7699 20587
rect 11529 20553 11563 20587
rect 13645 20553 13679 20587
rect 17601 20553 17635 20587
rect 19533 20553 19567 20587
rect 20637 20553 20671 20587
rect 32137 20553 32171 20587
rect 6745 20485 6779 20519
rect 8576 20485 8610 20519
rect 10149 20485 10183 20519
rect 11713 20485 11747 20519
rect 12817 20485 12851 20519
rect 13001 20485 13035 20519
rect 18420 20485 18454 20519
rect 21097 20485 21131 20519
rect 22192 20485 22226 20519
rect 23765 20485 23799 20519
rect 32597 20485 32631 20519
rect 36001 20485 36035 20519
rect 7113 20417 7147 20451
rect 10379 20417 10413 20451
rect 10517 20417 10551 20451
rect 10609 20420 10643 20454
rect 10793 20417 10827 20451
rect 11897 20417 11931 20451
rect 13461 20417 13495 20451
rect 13645 20417 13679 20451
rect 14749 20417 14783 20451
rect 18153 20417 18187 20451
rect 23949 20417 23983 20451
rect 24133 20417 24167 20451
rect 29101 20417 29135 20451
rect 30389 20417 30423 20451
rect 32321 20417 32355 20451
rect 32413 20417 32447 20451
rect 35909 20417 35943 20451
rect 36093 20417 36127 20451
rect 36277 20417 36311 20451
rect 8309 20349 8343 20383
rect 14657 20349 14691 20383
rect 21925 20349 21959 20383
rect 28825 20349 28859 20383
rect 30113 20349 30147 20383
rect 35725 20281 35759 20315
rect 9689 20213 9723 20247
rect 14381 20213 14415 20247
rect 14565 20213 14599 20247
rect 15209 20213 15243 20247
rect 23305 20213 23339 20247
rect 32321 20213 32355 20247
rect 10057 20009 10091 20043
rect 11897 20009 11931 20043
rect 14197 20009 14231 20043
rect 21833 20009 21867 20043
rect 22477 20009 22511 20043
rect 35081 20009 35115 20043
rect 40233 20009 40267 20043
rect 6377 19941 6411 19975
rect 14657 19941 14691 19975
rect 5641 19873 5675 19907
rect 11345 19873 11379 19907
rect 26341 19873 26375 19907
rect 2513 19805 2547 19839
rect 9597 19805 9631 19839
rect 12725 19805 12759 19839
rect 12817 19805 12851 19839
rect 12909 19805 12943 19839
rect 13093 19805 13127 19839
rect 15439 19805 15473 19839
rect 15577 19805 15611 19839
rect 15669 19805 15703 19839
rect 15853 19805 15887 19839
rect 22661 19805 22695 19839
rect 30941 19805 30975 19839
rect 32781 19805 32815 19839
rect 35265 19805 35299 19839
rect 35449 19805 35483 19839
rect 35633 19805 35667 19839
rect 58173 19805 58207 19839
rect 4445 19737 4479 19771
rect 5457 19737 5491 19771
rect 6193 19737 6227 19771
rect 10241 19737 10275 19771
rect 10425 19737 10459 19771
rect 22845 19737 22879 19771
rect 28089 19737 28123 19771
rect 28549 19737 28583 19771
rect 31125 19737 31159 19771
rect 32597 19737 32631 19771
rect 35357 19737 35391 19771
rect 2329 19669 2363 19703
rect 6929 19669 6963 19703
rect 12449 19669 12483 19703
rect 15209 19669 15243 19703
rect 30757 19669 30791 19703
rect 32965 19669 32999 19703
rect 2421 19465 2455 19499
rect 3893 19465 3927 19499
rect 12817 19465 12851 19499
rect 18337 19465 18371 19499
rect 27169 19465 27203 19499
rect 32781 19465 32815 19499
rect 38577 19465 38611 19499
rect 41061 19465 41095 19499
rect 10609 19397 10643 19431
rect 10793 19397 10827 19431
rect 29377 19397 29411 19431
rect 31309 19397 31343 19431
rect 39712 19397 39746 19431
rect 2605 19329 2639 19363
rect 10057 19329 10091 19363
rect 11805 19329 11839 19363
rect 11897 19329 11931 19363
rect 11989 19329 12023 19363
rect 12173 19329 12207 19363
rect 13001 19329 13035 19363
rect 13185 19329 13219 19363
rect 15393 19329 15427 19363
rect 15485 19329 15519 19363
rect 15577 19329 15611 19363
rect 15761 19329 15795 19363
rect 17509 19329 17543 19363
rect 18245 19329 18279 19363
rect 18429 19329 18463 19363
rect 26985 19329 27019 19363
rect 29193 19329 29227 19363
rect 29469 19329 29503 19363
rect 29561 19329 29595 19363
rect 30665 19329 30699 19363
rect 30849 19329 30883 19363
rect 30941 19329 30975 19363
rect 31033 19329 31067 19363
rect 33894 19329 33928 19363
rect 34161 19329 34195 19363
rect 35909 19329 35943 19363
rect 39957 19329 39991 19363
rect 40417 19329 40451 19363
rect 40580 19335 40614 19369
rect 40680 19335 40714 19369
rect 40785 19329 40819 19363
rect 2789 19261 2823 19295
rect 3985 19261 4019 19295
rect 4077 19261 4111 19295
rect 9965 19261 9999 19295
rect 10977 19261 11011 19295
rect 14657 19261 14691 19295
rect 17785 19261 17819 19295
rect 18889 19261 18923 19295
rect 32137 19261 32171 19295
rect 36185 19261 36219 19295
rect 3525 19125 3559 19159
rect 5181 19125 5215 19159
rect 5733 19125 5767 19159
rect 6561 19125 6595 19159
rect 9689 19125 9723 19159
rect 9873 19125 9907 19159
rect 11529 19125 11563 19159
rect 15117 19125 15151 19159
rect 29745 19125 29779 19159
rect 3801 18921 3835 18955
rect 5733 18921 5767 18955
rect 10241 18921 10275 18955
rect 13553 18921 13587 18955
rect 16681 18921 16715 18955
rect 30849 18921 30883 18955
rect 33333 18921 33367 18955
rect 40233 18921 40267 18955
rect 3249 18853 3283 18887
rect 4261 18785 4295 18819
rect 4353 18785 4387 18819
rect 7757 18785 7791 18819
rect 19257 18785 19291 18819
rect 32229 18785 32263 18819
rect 36093 18785 36127 18819
rect 1869 18717 1903 18751
rect 2136 18717 2170 18751
rect 12173 18717 12207 18751
rect 15301 18717 15335 18751
rect 15557 18717 15591 18751
rect 17141 18717 17175 18751
rect 17408 18717 17442 18751
rect 19988 18717 20022 18751
rect 20085 18717 20119 18751
rect 20360 18717 20394 18751
rect 20453 18717 20487 18751
rect 24409 18717 24443 18751
rect 24777 18717 24811 18751
rect 29561 18717 29595 18751
rect 29745 18717 29779 18751
rect 29929 18717 29963 18751
rect 31962 18717 31996 18751
rect 32689 18717 32723 18751
rect 32873 18717 32907 18751
rect 32965 18717 32999 18751
rect 33057 18717 33091 18751
rect 36369 18717 36403 18751
rect 37013 18717 37047 18751
rect 37381 18717 37415 18751
rect 40049 18717 40083 18751
rect 58173 18717 58207 18751
rect 5825 18649 5859 18683
rect 7490 18649 7524 18683
rect 12440 18649 12474 18683
rect 20177 18649 20211 18683
rect 24593 18649 24627 18683
rect 24685 18649 24719 18683
rect 26157 18649 26191 18683
rect 26341 18649 26375 18683
rect 26985 18649 27019 18683
rect 27169 18649 27203 18683
rect 29837 18649 29871 18683
rect 37105 18649 37139 18683
rect 37197 18649 37231 18683
rect 39865 18649 39899 18683
rect 4169 18581 4203 18615
rect 6377 18581 6411 18615
rect 8309 18581 8343 18615
rect 11345 18581 11379 18615
rect 18521 18581 18555 18615
rect 19809 18581 19843 18615
rect 21465 18581 21499 18615
rect 23673 18581 23707 18615
rect 24961 18581 24995 18615
rect 25973 18581 26007 18615
rect 26801 18581 26835 18615
rect 30113 18581 30147 18615
rect 36829 18581 36863 18615
rect 4629 18377 4663 18411
rect 6837 18377 6871 18411
rect 8125 18377 8159 18411
rect 16681 18377 16715 18411
rect 18337 18377 18371 18411
rect 21925 18377 21959 18411
rect 25053 18377 25087 18411
rect 29193 18377 29227 18411
rect 32597 18377 32631 18411
rect 35265 18377 35299 18411
rect 9864 18309 9898 18343
rect 15761 18309 15795 18343
rect 19533 18309 19567 18343
rect 36553 18309 36587 18343
rect 40969 18309 41003 18343
rect 1777 18241 1811 18275
rect 2421 18241 2455 18275
rect 2677 18241 2711 18275
rect 5457 18241 5491 18275
rect 7021 18241 7055 18275
rect 7389 18241 7423 18275
rect 7573 18241 7607 18275
rect 8401 18241 8435 18275
rect 15945 18241 15979 18275
rect 16129 18241 16163 18275
rect 16865 18241 16899 18275
rect 17049 18241 17083 18275
rect 17785 18241 17819 18275
rect 17877 18241 17911 18275
rect 18705 18241 18739 18275
rect 19257 18241 19291 18275
rect 19349 18241 19383 18275
rect 20133 18241 20167 18275
rect 20269 18241 20303 18275
rect 20361 18241 20395 18275
rect 20544 18241 20578 18275
rect 20637 18241 20671 18275
rect 21833 18241 21867 18275
rect 22017 18241 22051 18275
rect 23765 18241 23799 18275
rect 23949 18241 23983 18275
rect 24041 18241 24075 18275
rect 24133 18241 24167 18275
rect 26166 18241 26200 18275
rect 26433 18241 26467 18275
rect 26985 18241 27019 18275
rect 27252 18241 27286 18275
rect 29377 18241 29411 18275
rect 29653 18241 29687 18275
rect 30113 18241 30147 18275
rect 33977 18241 34011 18275
rect 36369 18241 36403 18275
rect 36461 18241 36495 18275
rect 36737 18241 36771 18275
rect 37381 18241 37415 18275
rect 39874 18241 39908 18275
rect 40141 18241 40175 18275
rect 40785 18241 40819 18275
rect 5089 18173 5123 18207
rect 5549 18173 5583 18207
rect 7205 18173 7239 18207
rect 7297 18173 7331 18207
rect 9597 18173 9631 18207
rect 18613 18173 18647 18207
rect 22477 18173 22511 18207
rect 22753 18173 22787 18207
rect 29561 18173 29595 18207
rect 30389 18173 30423 18207
rect 1961 18105 1995 18139
rect 5733 18105 5767 18139
rect 19993 18105 20027 18139
rect 36185 18105 36219 18139
rect 37565 18105 37599 18139
rect 3801 18037 3835 18071
rect 10977 18037 11011 18071
rect 11713 18037 11747 18071
rect 17509 18037 17543 18071
rect 17693 18037 17727 18071
rect 18521 18037 18555 18071
rect 21189 18037 21223 18071
rect 24317 18037 24351 18071
rect 28365 18037 28399 18071
rect 29653 18037 29687 18071
rect 33517 18037 33551 18071
rect 38761 18037 38795 18071
rect 40601 18037 40635 18071
rect 2421 17833 2455 17867
rect 4629 17833 4663 17867
rect 9229 17833 9263 17867
rect 11253 17833 11287 17867
rect 18613 17833 18647 17867
rect 25697 17833 25731 17867
rect 27445 17833 27479 17867
rect 30297 17833 30331 17867
rect 30481 17833 30515 17867
rect 39865 17833 39899 17867
rect 29745 17765 29779 17799
rect 2789 17697 2823 17731
rect 5457 17697 5491 17731
rect 8401 17697 8435 17731
rect 13553 17697 13587 17731
rect 19809 17697 19843 17731
rect 40969 17697 41003 17731
rect 2605 17629 2639 17663
rect 5549 17629 5583 17663
rect 9321 17629 9355 17663
rect 9413 17629 9447 17663
rect 11069 17629 11103 17663
rect 11253 17629 11287 17663
rect 17785 17629 17819 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 20085 17629 20119 17663
rect 20545 17629 20579 17663
rect 20821 17629 20855 17663
rect 23581 17629 23615 17663
rect 24409 17629 24443 17663
rect 24685 17629 24719 17663
rect 25973 17629 26007 17663
rect 26065 17629 26099 17663
rect 26157 17629 26191 17663
rect 26341 17629 26375 17663
rect 26801 17629 26835 17663
rect 26985 17629 27019 17663
rect 27077 17629 27111 17663
rect 27169 17629 27203 17663
rect 29561 17629 29595 17663
rect 30481 17629 30515 17663
rect 30573 17629 30607 17663
rect 30757 17629 30791 17663
rect 35081 17629 35115 17663
rect 35173 17629 35207 17663
rect 35449 17629 35483 17663
rect 36093 17629 36127 17663
rect 36461 17629 36495 17663
rect 37105 17629 37139 17663
rect 37289 17629 37323 17663
rect 37473 17629 37507 17663
rect 38761 17629 38795 17663
rect 40141 17629 40175 17663
rect 40230 17623 40264 17657
rect 40325 17626 40359 17660
rect 40509 17629 40543 17663
rect 5733 17561 5767 17595
rect 8134 17561 8168 17595
rect 11805 17561 11839 17595
rect 35265 17561 35299 17595
rect 36185 17561 36219 17595
rect 36277 17561 36311 17595
rect 37197 17561 37231 17595
rect 38577 17561 38611 17595
rect 5089 17493 5123 17527
rect 6469 17493 6503 17527
rect 7021 17493 7055 17527
rect 9045 17493 9079 17527
rect 9965 17493 9999 17527
rect 10517 17493 10551 17527
rect 17601 17493 17635 17527
rect 22109 17493 22143 17527
rect 34897 17493 34931 17527
rect 35909 17493 35943 17527
rect 36921 17493 36955 17527
rect 38945 17493 38979 17527
rect 3893 17289 3927 17323
rect 5457 17289 5491 17323
rect 7205 17289 7239 17323
rect 9321 17289 9355 17323
rect 12909 17289 12943 17323
rect 20637 17289 20671 17323
rect 21925 17289 21959 17323
rect 24501 17289 24535 17323
rect 27077 17289 27111 17323
rect 34023 17289 34057 17323
rect 39037 17289 39071 17323
rect 10241 17221 10275 17255
rect 11621 17221 11655 17255
rect 13277 17221 13311 17255
rect 39589 17221 39623 17255
rect 3709 17153 3743 17187
rect 4445 17153 4479 17187
rect 5733 17153 5767 17187
rect 7389 17153 7423 17187
rect 7757 17153 7791 17187
rect 7941 17153 7975 17187
rect 9873 17153 9907 17187
rect 10021 17153 10055 17187
rect 10149 17153 10183 17187
rect 10338 17153 10372 17187
rect 11529 17153 11563 17187
rect 11713 17153 11747 17187
rect 13049 17153 13083 17187
rect 13185 17153 13219 17187
rect 13405 17153 13439 17187
rect 13553 17153 13587 17187
rect 20545 17153 20579 17187
rect 20729 17153 20763 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 22477 17153 22511 17187
rect 22661 17153 22695 17187
rect 23765 17153 23799 17187
rect 24685 17153 24719 17187
rect 24961 17153 24995 17187
rect 37565 17153 37599 17187
rect 3249 17085 3283 17119
rect 7573 17085 7607 17119
rect 7665 17085 7699 17119
rect 21189 17085 21223 17119
rect 24041 17085 24075 17119
rect 24777 17085 24811 17119
rect 25605 17085 25639 17119
rect 33793 17085 33827 17119
rect 35081 17085 35115 17119
rect 35357 17085 35391 17119
rect 37289 17085 37323 17119
rect 4629 17017 4663 17051
rect 19993 17017 20027 17051
rect 22661 17017 22695 17051
rect 58173 17017 58207 17051
rect 6653 16949 6687 16983
rect 10517 16949 10551 16983
rect 12449 16949 12483 16983
rect 14105 16949 14139 16983
rect 18153 16949 18187 16983
rect 19533 16949 19567 16983
rect 24961 16949 24995 16983
rect 40877 16949 40911 16983
rect 5273 16745 5307 16779
rect 12725 16745 12759 16779
rect 13553 16745 13587 16779
rect 16405 16745 16439 16779
rect 17509 16745 17543 16779
rect 18245 16745 18279 16779
rect 19717 16745 19751 16779
rect 20361 16745 20395 16779
rect 21925 16745 21959 16779
rect 22661 16745 22695 16779
rect 24593 16745 24627 16779
rect 25329 16745 25363 16779
rect 26709 16745 26743 16779
rect 35909 16745 35943 16779
rect 11897 16677 11931 16711
rect 27813 16677 27847 16711
rect 37933 16677 37967 16711
rect 15301 16609 15335 16643
rect 16957 16609 16991 16643
rect 21373 16609 21407 16643
rect 23213 16609 23247 16643
rect 23765 16609 23799 16643
rect 26157 16609 26191 16643
rect 27077 16609 27111 16643
rect 29561 16609 29595 16643
rect 30389 16609 30423 16643
rect 32045 16609 32079 16643
rect 32873 16609 32907 16643
rect 33333 16609 33367 16643
rect 33609 16609 33643 16643
rect 37289 16609 37323 16643
rect 39313 16609 39347 16643
rect 4445 16541 4479 16575
rect 9965 16541 9999 16575
rect 10113 16541 10147 16575
rect 10241 16541 10275 16575
rect 10430 16541 10464 16575
rect 11253 16541 11287 16575
rect 11346 16541 11380 16575
rect 11759 16541 11793 16575
rect 12725 16541 12759 16575
rect 12909 16541 12943 16575
rect 13369 16541 13403 16575
rect 13553 16541 13587 16575
rect 14749 16541 14783 16575
rect 18061 16541 18095 16575
rect 18245 16541 18279 16575
rect 19809 16541 19843 16575
rect 20361 16541 20395 16575
rect 20545 16541 20579 16575
rect 22477 16541 22511 16575
rect 22661 16541 22695 16575
rect 23121 16541 23155 16575
rect 23305 16541 23339 16575
rect 24593 16541 24627 16575
rect 24685 16541 24719 16575
rect 24869 16541 24903 16575
rect 26893 16541 26927 16575
rect 30205 16541 30239 16575
rect 34805 16541 34839 16575
rect 34989 16541 35023 16575
rect 35081 16541 35115 16575
rect 35173 16541 35207 16575
rect 10333 16473 10367 16507
rect 11529 16473 11563 16507
rect 11621 16473 11655 16507
rect 14565 16473 14599 16507
rect 27629 16473 27663 16507
rect 35449 16473 35483 16507
rect 37022 16473 37056 16507
rect 39046 16473 39080 16507
rect 4261 16405 4295 16439
rect 10609 16405 10643 16439
rect 24409 16405 24443 16439
rect 5457 16201 5491 16235
rect 10517 16201 10551 16235
rect 19349 16201 19383 16235
rect 20821 16201 20855 16235
rect 21833 16201 21867 16235
rect 22753 16201 22787 16235
rect 35173 16201 35207 16235
rect 37473 16201 37507 16235
rect 3157 16133 3191 16167
rect 12173 16133 12207 16167
rect 18429 16133 18463 16167
rect 31585 16133 31619 16167
rect 35357 16133 35391 16167
rect 38209 16133 38243 16167
rect 2421 16065 2455 16099
rect 7665 16065 7699 16099
rect 7757 16065 7791 16099
rect 10425 16065 10459 16099
rect 10609 16065 10643 16099
rect 12081 16065 12115 16099
rect 12265 16065 12299 16099
rect 13277 16065 13311 16099
rect 13553 16065 13587 16099
rect 14657 16065 14691 16099
rect 14749 16065 14783 16099
rect 14841 16065 14875 16099
rect 15025 16065 15059 16099
rect 15485 16065 15519 16099
rect 15669 16065 15703 16099
rect 15761 16065 15795 16099
rect 15853 16065 15887 16099
rect 16957 16065 16991 16099
rect 17141 16065 17175 16099
rect 17233 16065 17267 16099
rect 17325 16065 17359 16099
rect 18061 16065 18095 16099
rect 18245 16065 18279 16099
rect 19257 16065 19291 16099
rect 19441 16065 19475 16099
rect 26249 16065 26283 16099
rect 27813 16065 27847 16099
rect 31217 16065 31251 16099
rect 31401 16065 31435 16099
rect 32137 16065 32171 16099
rect 32321 16065 32355 16099
rect 32413 16065 32447 16099
rect 32505 16065 32539 16099
rect 34621 16065 34655 16099
rect 35541 16065 35575 16099
rect 37289 16065 37323 16099
rect 38925 16065 38959 16099
rect 39037 16065 39071 16099
rect 39129 16065 39163 16099
rect 39313 16065 39347 16099
rect 25053 15997 25087 16031
rect 27537 15997 27571 16031
rect 34345 15997 34379 16031
rect 38669 15997 38703 16031
rect 20177 15929 20211 15963
rect 2237 15861 2271 15895
rect 4629 15861 4663 15895
rect 7389 15861 7423 15895
rect 7573 15861 7607 15895
rect 9965 15861 9999 15895
rect 11621 15861 11655 15895
rect 14381 15861 14415 15895
rect 16129 15861 16163 15895
rect 17601 15861 17635 15895
rect 23857 15861 23891 15895
rect 26433 15861 26467 15895
rect 32781 15861 32815 15895
rect 58173 15861 58207 15895
rect 2513 15657 2547 15691
rect 4077 15657 4111 15691
rect 4721 15657 4755 15691
rect 7205 15657 7239 15691
rect 10425 15657 10459 15691
rect 12909 15657 12943 15691
rect 23213 15657 23247 15691
rect 23489 15657 23523 15691
rect 25145 15657 25179 15691
rect 25697 15657 25731 15691
rect 26525 15657 26559 15691
rect 29837 15657 29871 15691
rect 34069 15657 34103 15691
rect 7297 15521 7331 15555
rect 10517 15521 10551 15555
rect 14105 15521 14139 15555
rect 18705 15521 18739 15555
rect 23581 15521 23615 15555
rect 27169 15521 27203 15555
rect 35081 15521 35115 15555
rect 2145 15453 2179 15487
rect 2329 15453 2363 15487
rect 3065 15453 3099 15487
rect 3893 15453 3927 15487
rect 5549 15453 5583 15487
rect 5641 15453 5675 15487
rect 7389 15453 7423 15487
rect 8953 15453 8987 15487
rect 9229 15453 9263 15487
rect 10609 15453 10643 15487
rect 12725 15453 12759 15487
rect 14372 15453 14406 15487
rect 16681 15453 16715 15487
rect 20453 15453 20487 15487
rect 22109 15453 22143 15487
rect 23397 15453 23431 15487
rect 23673 15453 23707 15487
rect 24409 15453 24443 15487
rect 26433 15453 26467 15487
rect 26617 15453 26651 15487
rect 28273 15453 28307 15487
rect 30389 15453 30423 15487
rect 30573 15453 30607 15487
rect 30665 15453 30699 15487
rect 30757 15453 30791 15487
rect 32873 15453 32907 15487
rect 34713 15453 34747 15487
rect 34897 15453 34931 15487
rect 35541 15453 35575 15487
rect 35725 15453 35759 15487
rect 36829 15453 36863 15487
rect 37657 15453 37691 15487
rect 37841 15453 37875 15487
rect 16926 15385 16960 15419
rect 20637 15385 20671 15419
rect 28089 15385 28123 15419
rect 31033 15385 31067 15419
rect 32606 15385 32640 15419
rect 36185 15385 36219 15419
rect 37013 15385 37047 15419
rect 3249 15317 3283 15351
rect 5181 15317 5215 15351
rect 5825 15317 5859 15351
rect 7021 15317 7055 15351
rect 10241 15317 10275 15351
rect 12173 15317 12207 15351
rect 15485 15317 15519 15351
rect 18061 15317 18095 15351
rect 19809 15317 19843 15351
rect 20269 15317 20303 15351
rect 28457 15317 28491 15351
rect 31493 15317 31527 15351
rect 35725 15317 35759 15351
rect 37197 15317 37231 15351
rect 38025 15317 38059 15351
rect 2973 15113 3007 15147
rect 14197 15113 14231 15147
rect 15117 15113 15151 15147
rect 16681 15113 16715 15147
rect 22845 15113 22879 15147
rect 29837 15113 29871 15147
rect 31217 15113 31251 15147
rect 34069 15113 34103 15147
rect 34989 15113 35023 15147
rect 38669 15113 38703 15147
rect 16865 15045 16899 15079
rect 20922 15045 20956 15079
rect 22477 15045 22511 15079
rect 22569 15045 22603 15079
rect 23581 15045 23615 15079
rect 25789 15045 25823 15079
rect 31585 15045 31619 15079
rect 36737 15045 36771 15079
rect 38117 15045 38151 15079
rect 39782 15045 39816 15079
rect 1593 14977 1627 15011
rect 1860 14977 1894 15011
rect 3433 14977 3467 15011
rect 3689 14977 3723 15011
rect 6377 14977 6411 15011
rect 6644 14977 6678 15011
rect 15301 14977 15335 15011
rect 15485 14977 15519 15011
rect 17049 14977 17083 15011
rect 17969 14977 18003 15011
rect 18225 14977 18259 15011
rect 22293 14977 22327 15011
rect 22661 14977 22695 15011
rect 23305 14977 23339 15011
rect 23489 14977 23523 15011
rect 23673 14977 23707 15011
rect 24501 14977 24535 15011
rect 24777 14977 24811 15011
rect 25605 14977 25639 15011
rect 28713 14977 28747 15011
rect 31401 14977 31435 15011
rect 33250 14977 33284 15011
rect 33517 14977 33551 15011
rect 34805 14977 34839 15011
rect 37473 14977 37507 15011
rect 37657 14977 37691 15011
rect 37749 14977 37783 15011
rect 37841 14977 37875 15011
rect 40049 14977 40083 15011
rect 21189 14909 21223 14943
rect 24593 14909 24627 14943
rect 28457 14909 28491 14943
rect 34621 14909 34655 14943
rect 19349 14841 19383 14875
rect 24317 14841 24351 14875
rect 4813 14773 4847 14807
rect 7757 14773 7791 14807
rect 12449 14773 12483 14807
rect 19809 14773 19843 14807
rect 23857 14773 23891 14807
rect 24501 14773 24535 14807
rect 25973 14773 26007 14807
rect 32137 14773 32171 14807
rect 2513 14569 2547 14603
rect 3801 14569 3835 14603
rect 6929 14569 6963 14603
rect 7481 14569 7515 14603
rect 11621 14569 11655 14603
rect 20913 14569 20947 14603
rect 24593 14569 24627 14603
rect 28549 14569 28583 14603
rect 34161 14569 34195 14603
rect 23581 14501 23615 14535
rect 2973 14433 3007 14467
rect 3157 14433 3191 14467
rect 4169 14433 4203 14467
rect 5457 14433 5491 14467
rect 6469 14433 6503 14467
rect 6561 14433 6595 14467
rect 10977 14433 11011 14467
rect 36553 14433 36587 14467
rect 38761 14433 38795 14467
rect 2881 14365 2915 14399
rect 3985 14365 4019 14399
rect 5549 14365 5583 14399
rect 6193 14365 6227 14399
rect 6377 14365 6411 14399
rect 6745 14365 6779 14399
rect 20269 14365 20303 14399
rect 20453 14362 20487 14396
rect 20545 14365 20579 14399
rect 20683 14365 20717 14399
rect 23029 14365 23063 14399
rect 23397 14365 23431 14399
rect 24593 14365 24627 14399
rect 24685 14365 24719 14399
rect 24869 14365 24903 14399
rect 27893 14365 27927 14399
rect 28089 14365 28123 14399
rect 28181 14365 28215 14399
rect 28273 14365 28307 14399
rect 29745 14365 29779 14399
rect 34897 14365 34931 14399
rect 35081 14365 35115 14399
rect 36277 14365 36311 14399
rect 37197 14365 37231 14399
rect 38485 14365 38519 14399
rect 39865 14365 39899 14399
rect 40141 14365 40175 14399
rect 58173 14365 58207 14399
rect 5089 14297 5123 14331
rect 10710 14297 10744 14331
rect 11529 14297 11563 14331
rect 21465 14297 21499 14331
rect 23213 14297 23247 14331
rect 23305 14297 23339 14331
rect 25881 14297 25915 14331
rect 26065 14297 26099 14331
rect 26249 14297 26283 14331
rect 29561 14297 29595 14331
rect 5733 14229 5767 14263
rect 9597 14229 9631 14263
rect 24409 14229 24443 14263
rect 25329 14229 25363 14263
rect 26709 14229 26743 14263
rect 27353 14229 27387 14263
rect 29929 14229 29963 14263
rect 35081 14229 35115 14263
rect 37105 14229 37139 14263
rect 3433 14025 3467 14059
rect 5089 14025 5123 14059
rect 10149 14025 10183 14059
rect 23489 14025 23523 14059
rect 37841 14025 37875 14059
rect 38761 14025 38795 14059
rect 5549 13957 5583 13991
rect 17233 13957 17267 13991
rect 21097 13957 21131 13991
rect 27445 13957 27479 13991
rect 32965 13957 32999 13991
rect 33149 13957 33183 13991
rect 35173 13957 35207 13991
rect 5457 13889 5491 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 9965 13889 9999 13923
rect 13205 13889 13239 13923
rect 17417 13889 17451 13923
rect 24613 13889 24647 13923
rect 26019 13889 26053 13923
rect 26157 13889 26191 13923
rect 26249 13889 26283 13923
rect 26433 13889 26467 13923
rect 29909 13889 29943 13923
rect 34989 13889 35023 13923
rect 37749 13889 37783 13923
rect 39874 13889 39908 13923
rect 40141 13889 40175 13923
rect 5733 13821 5767 13855
rect 6469 13821 6503 13855
rect 9689 13821 9723 13855
rect 9781 13821 9815 13855
rect 13461 13821 13495 13855
rect 17601 13821 17635 13855
rect 24869 13821 24903 13855
rect 29653 13821 29687 13855
rect 35357 13821 35391 13855
rect 12081 13753 12115 13787
rect 31033 13753 31067 13787
rect 14933 13685 14967 13719
rect 19993 13685 20027 13719
rect 25789 13685 25823 13719
rect 28733 13685 28767 13719
rect 17877 13481 17911 13515
rect 19257 13481 19291 13515
rect 22845 13481 22879 13515
rect 26985 13481 27019 13515
rect 28733 13481 28767 13515
rect 29561 13481 29595 13515
rect 32045 13481 32079 13515
rect 36093 13481 36127 13515
rect 38853 13481 38887 13515
rect 16037 13413 16071 13447
rect 24961 13413 24995 13447
rect 39865 13413 39899 13447
rect 21465 13345 21499 13379
rect 33057 13345 33091 13379
rect 9965 13277 9999 13311
rect 13369 13277 13403 13311
rect 14427 13277 14461 13311
rect 14565 13277 14599 13311
rect 14678 13274 14712 13308
rect 14841 13277 14875 13311
rect 16589 13277 16623 13311
rect 19441 13277 19475 13311
rect 20177 13277 20211 13311
rect 20361 13277 20395 13311
rect 21732 13277 21766 13311
rect 26065 13277 26099 13311
rect 26157 13277 26191 13311
rect 26254 13277 26288 13311
rect 26445 13277 26479 13311
rect 27261 13277 27295 13311
rect 27353 13277 27387 13311
rect 27445 13274 27479 13308
rect 27629 13277 27663 13311
rect 28089 13277 28123 13311
rect 28252 13271 28286 13305
rect 28365 13277 28399 13311
rect 28503 13277 28537 13311
rect 32781 13277 32815 13311
rect 34713 13277 34747 13311
rect 37381 13277 37415 13311
rect 37473 13277 37507 13311
rect 37565 13277 37599 13311
rect 37749 13277 37783 13311
rect 38209 13277 38243 13311
rect 38393 13277 38427 13311
rect 38485 13277 38519 13311
rect 38577 13277 38611 13311
rect 40049 13277 40083 13311
rect 58173 13277 58207 13311
rect 10232 13209 10266 13243
rect 13185 13209 13219 13243
rect 13553 13209 13587 13243
rect 25145 13209 25179 13243
rect 25329 13209 25363 13243
rect 34958 13209 34992 13243
rect 36645 13209 36679 13243
rect 11345 13141 11379 13175
rect 14197 13141 14231 13175
rect 15393 13141 15427 13175
rect 20545 13141 20579 13175
rect 25789 13141 25823 13175
rect 37105 13141 37139 13175
rect 3341 12937 3375 12971
rect 4261 12937 4295 12971
rect 11805 12937 11839 12971
rect 21281 12937 21315 12971
rect 24961 12937 24995 12971
rect 27997 12937 28031 12971
rect 31585 12937 31619 12971
rect 33241 12937 33275 12971
rect 37657 12937 37691 12971
rect 12940 12869 12974 12903
rect 15485 12869 15519 12903
rect 15669 12869 15703 12903
rect 26074 12869 26108 12903
rect 29009 12869 29043 12903
rect 31309 12869 31343 12903
rect 39690 12869 39724 12903
rect 2145 12801 2179 12835
rect 2329 12801 2363 12835
rect 7858 12801 7892 12835
rect 8852 12801 8886 12835
rect 14427 12801 14461 12835
rect 14565 12801 14599 12835
rect 14657 12807 14691 12841
rect 14841 12801 14875 12835
rect 17794 12801 17828 12835
rect 18061 12801 18095 12835
rect 20315 12801 20349 12835
rect 20453 12801 20487 12835
rect 20545 12801 20579 12835
rect 20729 12801 20763 12835
rect 26341 12801 26375 12835
rect 29745 12801 29779 12835
rect 29837 12801 29871 12835
rect 29929 12801 29963 12835
rect 30113 12801 30147 12835
rect 31033 12801 31067 12835
rect 31217 12801 31251 12835
rect 31401 12801 31435 12835
rect 32413 12801 32447 12835
rect 32505 12801 32539 12835
rect 32597 12801 32631 12835
rect 32781 12801 32815 12835
rect 35817 12801 35851 12835
rect 37289 12801 37323 12835
rect 37473 12801 37507 12835
rect 39957 12801 39991 12835
rect 3433 12733 3467 12767
rect 3617 12733 3651 12767
rect 8125 12733 8159 12767
rect 8585 12733 8619 12767
rect 13185 12733 13219 12767
rect 19165 12733 19199 12767
rect 19441 12733 19475 12767
rect 35541 12733 35575 12767
rect 2973 12665 3007 12699
rect 6745 12665 6779 12699
rect 14197 12665 14231 12699
rect 16681 12665 16715 12699
rect 38577 12665 38611 12699
rect 2513 12597 2547 12631
rect 9965 12597 9999 12631
rect 15301 12597 15335 12631
rect 20085 12597 20119 12631
rect 27077 12597 27111 12631
rect 29469 12597 29503 12631
rect 32137 12597 32171 12631
rect 10517 12393 10551 12427
rect 15485 12393 15519 12427
rect 17509 12393 17543 12427
rect 21189 12393 21223 12427
rect 29929 12393 29963 12427
rect 36369 12393 36403 12427
rect 3249 12325 3283 12359
rect 7941 12325 7975 12359
rect 22753 12325 22787 12359
rect 31401 12325 31435 12359
rect 5733 12257 5767 12291
rect 10149 12257 10183 12291
rect 11069 12257 11103 12291
rect 19809 12257 19843 12291
rect 33241 12257 33275 12291
rect 1869 12189 1903 12223
rect 5825 12189 5859 12223
rect 9781 12189 9815 12223
rect 9965 12189 9999 12223
rect 10057 12189 10091 12223
rect 10333 12189 10367 12223
rect 13185 12189 13219 12223
rect 14105 12189 14139 12223
rect 17785 12189 17819 12223
rect 17877 12189 17911 12223
rect 17969 12189 18003 12223
rect 18153 12189 18187 12223
rect 20076 12189 20110 12223
rect 29745 12189 29779 12223
rect 30849 12189 30883 12223
rect 31217 12189 31251 12223
rect 32974 12189 33008 12223
rect 34161 12189 34195 12223
rect 34989 12189 35023 12223
rect 35081 12189 35115 12223
rect 35173 12189 35207 12223
rect 35357 12189 35391 12223
rect 2136 12121 2170 12155
rect 6653 12121 6687 12155
rect 13369 12121 13403 12155
rect 13553 12121 13587 12155
rect 14372 12121 14406 12155
rect 16681 12121 16715 12155
rect 16865 12121 16899 12155
rect 19349 12121 19383 12155
rect 22017 12121 22051 12155
rect 22569 12121 22603 12155
rect 29561 12121 29595 12155
rect 31033 12121 31067 12155
rect 31125 12121 31159 12155
rect 34713 12121 34747 12155
rect 36277 12121 36311 12155
rect 5365 12053 5399 12087
rect 6009 12053 6043 12087
rect 8953 12053 8987 12087
rect 17049 12053 17083 12087
rect 18705 12053 18739 12087
rect 25697 12053 25731 12087
rect 31861 12053 31895 12087
rect 38025 12053 38059 12087
rect 2237 11849 2271 11883
rect 7205 11849 7239 11883
rect 9137 11849 9171 11883
rect 11713 11849 11747 11883
rect 14657 11849 14691 11883
rect 16681 11849 16715 11883
rect 19625 11849 19659 11883
rect 27261 11849 27295 11883
rect 31585 11849 31619 11883
rect 25973 11781 26007 11815
rect 28396 11781 28430 11815
rect 31309 11781 31343 11815
rect 2421 11713 2455 11747
rect 3413 11713 3447 11747
rect 5733 11713 5767 11747
rect 6469 11713 6503 11747
rect 6653 11713 6687 11747
rect 7021 11713 7055 11747
rect 8401 11713 8435 11747
rect 8585 11713 8619 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 11529 11713 11563 11747
rect 14887 11713 14921 11747
rect 15006 11713 15040 11747
rect 15106 11713 15140 11747
rect 15301 11713 15335 11747
rect 17794 11713 17828 11747
rect 18061 11713 18095 11747
rect 19533 11713 19567 11747
rect 22569 11713 22603 11747
rect 22753 11713 22787 11747
rect 24961 11713 24995 11747
rect 25789 11713 25823 11747
rect 28641 11713 28675 11747
rect 31033 11713 31067 11747
rect 31217 11713 31251 11747
rect 31401 11713 31435 11747
rect 32781 11713 32815 11747
rect 36093 11713 36127 11747
rect 38485 11713 38519 11747
rect 3157 11645 3191 11679
rect 6745 11645 6779 11679
rect 6837 11645 6871 11679
rect 8677 11645 8711 11679
rect 9689 11645 9723 11679
rect 32505 11645 32539 11679
rect 33793 11645 33827 11679
rect 38209 11645 38243 11679
rect 5549 11577 5583 11611
rect 24777 11577 24811 11611
rect 58173 11577 58207 11611
rect 4537 11509 4571 11543
rect 7757 11509 7791 11543
rect 15761 11509 15795 11543
rect 18889 11509 18923 11543
rect 22385 11509 22419 11543
rect 36277 11509 36311 11543
rect 39037 11509 39071 11543
rect 3249 11305 3283 11339
rect 7021 11305 7055 11339
rect 17509 11305 17543 11339
rect 18705 11305 18739 11339
rect 24409 11305 24443 11339
rect 26801 11305 26835 11339
rect 29561 11305 29595 11339
rect 32045 11305 32079 11339
rect 35909 11305 35943 11339
rect 11161 11237 11195 11271
rect 28457 11237 28491 11271
rect 37749 11237 37783 11271
rect 4629 11169 4663 11203
rect 5641 11169 5675 11203
rect 5825 11169 5859 11203
rect 6377 11169 6411 11203
rect 7481 11169 7515 11203
rect 32781 11169 32815 11203
rect 33057 11169 33091 11203
rect 3065 11101 3099 11135
rect 4353 11101 4387 11135
rect 6745 11101 6779 11135
rect 6837 11101 6871 11135
rect 12449 11101 12483 11135
rect 12633 11101 12667 11135
rect 17785 11101 17819 11135
rect 17877 11101 17911 11135
rect 17969 11101 18003 11135
rect 18153 11101 18187 11135
rect 22109 11101 22143 11135
rect 22845 11101 22879 11135
rect 22934 11101 22968 11135
rect 23034 11101 23068 11135
rect 23225 11101 23259 11135
rect 26893 11101 26927 11135
rect 29009 11101 29043 11135
rect 29745 11101 29779 11135
rect 30113 11101 30147 11135
rect 31861 11101 31895 11135
rect 35081 11101 35115 11135
rect 36461 11101 36495 11135
rect 38669 11101 38703 11135
rect 38832 11101 38866 11135
rect 38945 11101 38979 11135
rect 39083 11101 39117 11135
rect 5549 11033 5583 11067
rect 10977 11033 11011 11067
rect 29837 11033 29871 11067
rect 29929 11033 29963 11067
rect 31677 11033 31711 11067
rect 35265 11033 35299 11067
rect 5181 10965 5215 10999
rect 12265 10965 12299 10999
rect 22569 10965 22603 10999
rect 34897 10965 34931 10999
rect 39313 10965 39347 10999
rect 4077 10761 4111 10795
rect 12357 10761 12391 10795
rect 22385 10761 22419 10795
rect 23581 10761 23615 10795
rect 28181 10761 28215 10795
rect 30113 10761 30147 10795
rect 37657 10761 37691 10795
rect 12817 10693 12851 10727
rect 20453 10693 20487 10727
rect 22109 10693 22143 10727
rect 27905 10693 27939 10727
rect 28641 10693 28675 10727
rect 31217 10693 31251 10727
rect 4261 10625 4295 10659
rect 6653 10625 6687 10659
rect 7849 10625 7883 10659
rect 11621 10625 11655 10659
rect 12725 10625 12759 10659
rect 13553 10625 13587 10659
rect 18889 10625 18923 10659
rect 19717 10625 19751 10659
rect 20269 10625 20303 10659
rect 21833 10625 21867 10659
rect 22017 10625 22051 10659
rect 22201 10625 22235 10659
rect 23765 10625 23799 10659
rect 24409 10625 24443 10659
rect 27629 10625 27663 10659
rect 27813 10625 27847 10659
rect 27997 10625 28031 10659
rect 31033 10625 31067 10659
rect 31125 10625 31159 10659
rect 31401 10625 31435 10659
rect 32137 10625 32171 10659
rect 32321 10625 32355 10659
rect 32416 10631 32450 10665
rect 32505 10625 32539 10659
rect 34529 10625 34563 10659
rect 34796 10625 34830 10659
rect 37289 10625 37323 10659
rect 37473 10625 37507 10659
rect 39598 10625 39632 10659
rect 39865 10625 39899 10659
rect 4445 10557 4479 10591
rect 6377 10557 6411 10591
rect 7665 10557 7699 10591
rect 12909 10557 12943 10591
rect 23029 10557 23063 10591
rect 23949 10557 23983 10591
rect 24685 10557 24719 10591
rect 11805 10489 11839 10523
rect 19073 10489 19107 10523
rect 30849 10489 30883 10523
rect 38485 10489 38519 10523
rect 8861 10421 8895 10455
rect 18337 10421 18371 10455
rect 32781 10421 32815 10455
rect 35909 10421 35943 10455
rect 58173 10421 58207 10455
rect 10885 10217 10919 10251
rect 22201 10217 22235 10251
rect 25053 10217 25087 10251
rect 31953 10217 31987 10251
rect 32505 10217 32539 10251
rect 34713 10217 34747 10251
rect 35817 10217 35851 10251
rect 8953 10149 8987 10183
rect 17233 10149 17267 10183
rect 6101 10081 6135 10115
rect 9597 10081 9631 10115
rect 13093 10081 13127 10115
rect 16497 10081 16531 10115
rect 24501 10081 24535 10115
rect 28181 10081 28215 10115
rect 28457 10081 28491 10115
rect 29837 10081 29871 10115
rect 2605 10013 2639 10047
rect 6377 10013 6411 10047
rect 7205 10013 7239 10047
rect 7941 10013 7975 10047
rect 8033 10013 8067 10047
rect 13277 10013 13311 10047
rect 20821 10013 20855 10047
rect 21088 10013 21122 10047
rect 23489 10013 23523 10047
rect 23581 10013 23615 10047
rect 23673 10013 23707 10047
rect 23857 10013 23891 10047
rect 24409 10013 24443 10047
rect 24593 10013 24627 10047
rect 29561 10013 29595 10047
rect 34069 10013 34103 10047
rect 34989 10013 35023 10047
rect 35081 10013 35115 10047
rect 35194 10013 35228 10047
rect 35357 10013 35391 10047
rect 36645 10013 36679 10047
rect 36829 10013 36863 10047
rect 12173 9945 12207 9979
rect 16313 9945 16347 9979
rect 17049 9945 17083 9979
rect 27353 9945 27387 9979
rect 27537 9945 27571 9979
rect 31585 9945 31619 9979
rect 31769 9945 31803 9979
rect 38025 9945 38059 9979
rect 38209 9945 38243 9979
rect 2421 9877 2455 9911
rect 7297 9877 7331 9911
rect 8217 9877 8251 9911
rect 9321 9877 9355 9911
rect 9413 9877 9447 9911
rect 13461 9877 13495 9911
rect 18705 9877 18739 9911
rect 19625 9877 19659 9911
rect 22661 9877 22695 9911
rect 23213 9877 23247 9911
rect 27721 9877 27755 9911
rect 36461 9877 36495 9911
rect 37289 9877 37323 9911
rect 37841 9877 37875 9911
rect 9689 9673 9723 9707
rect 11713 9673 11747 9707
rect 24501 9673 24535 9707
rect 39957 9673 39991 9707
rect 2412 9605 2446 9639
rect 10149 9605 10183 9639
rect 19165 9605 19199 9639
rect 33250 9605 33284 9639
rect 34621 9605 34655 9639
rect 38117 9605 38151 9639
rect 38822 9605 38856 9639
rect 4353 9537 4387 9571
rect 6561 9537 6595 9571
rect 8309 9537 8343 9571
rect 8576 9537 8610 9571
rect 10425 9537 10459 9571
rect 12173 9537 12207 9571
rect 12440 9537 12474 9571
rect 15209 9537 15243 9571
rect 18337 9537 18371 9571
rect 19809 9537 19843 9571
rect 19993 9537 20027 9571
rect 22661 9537 22695 9571
rect 22928 9537 22962 9571
rect 24685 9537 24719 9571
rect 24869 9537 24903 9571
rect 25329 9537 25363 9571
rect 25513 9537 25547 9571
rect 27169 9537 27203 9571
rect 27629 9537 27663 9571
rect 27905 9537 27939 9571
rect 29837 9537 29871 9571
rect 34529 9537 34563 9571
rect 34713 9537 34747 9571
rect 34897 9537 34931 9571
rect 36093 9537 36127 9571
rect 36277 9537 36311 9571
rect 36369 9537 36403 9571
rect 36461 9537 36495 9571
rect 37461 9537 37495 9571
rect 37636 9543 37670 9577
rect 37736 9543 37770 9577
rect 37887 9537 37921 9571
rect 38577 9537 38611 9571
rect 2145 9469 2179 9503
rect 4445 9469 4479 9503
rect 4629 9469 4663 9503
rect 6837 9469 6871 9503
rect 10333 9469 10367 9503
rect 10793 9469 10827 9503
rect 17325 9469 17359 9503
rect 19901 9469 19935 9503
rect 20453 9469 20487 9503
rect 20729 9469 20763 9503
rect 29561 9469 29595 9503
rect 33517 9469 33551 9503
rect 3525 9401 3559 9435
rect 19349 9401 19383 9435
rect 34345 9401 34379 9435
rect 35541 9401 35575 9435
rect 3985 9333 4019 9367
rect 5273 9333 5307 9367
rect 13553 9333 13587 9367
rect 14565 9333 14599 9367
rect 15301 9333 15335 9367
rect 17877 9333 17911 9367
rect 18521 9333 18555 9367
rect 24041 9333 24075 9367
rect 25697 9333 25731 9367
rect 26985 9333 27019 9367
rect 32137 9333 32171 9367
rect 36737 9333 36771 9367
rect 2697 9129 2731 9163
rect 8953 9129 8987 9163
rect 12817 9129 12851 9163
rect 18613 9129 18647 9163
rect 23489 9129 23523 9163
rect 28917 9129 28951 9163
rect 31217 9129 31251 9163
rect 37749 9129 37783 9163
rect 4169 9061 4203 9095
rect 10057 8993 10091 9027
rect 10793 8993 10827 9027
rect 11161 8993 11195 9027
rect 12265 8993 12299 9027
rect 12357 8993 12391 9027
rect 17233 8993 17267 9027
rect 19901 8993 19935 9027
rect 20821 8993 20855 9027
rect 21097 8993 21131 9027
rect 25605 8993 25639 9027
rect 27629 8993 27663 9027
rect 36369 8993 36403 9027
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 4353 8925 4387 8959
rect 6377 8925 6411 8959
rect 6653 8925 6687 8959
rect 7665 8925 7699 8959
rect 9137 8925 9171 8959
rect 10149 8925 10183 8959
rect 11253 8925 11287 8959
rect 13369 8925 13403 8959
rect 15393 8925 15427 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 22937 8925 22971 8959
rect 23213 8925 23247 8959
rect 23305 8925 23339 8959
rect 27905 8925 27939 8959
rect 29837 8925 29871 8959
rect 36636 8925 36670 8959
rect 58173 8925 58207 8959
rect 9689 8857 9723 8891
rect 10333 8857 10367 8891
rect 15638 8857 15672 8891
rect 17500 8857 17534 8891
rect 23121 8857 23155 8891
rect 25872 8857 25906 8891
rect 30082 8857 30116 8891
rect 5181 8789 5215 8823
rect 7849 8789 7883 8823
rect 11437 8789 11471 8823
rect 12449 8789 12483 8823
rect 13553 8789 13587 8823
rect 16773 8789 16807 8823
rect 19349 8789 19383 8823
rect 26985 8789 27019 8823
rect 11713 8585 11747 8619
rect 13553 8585 13587 8619
rect 15577 8585 15611 8619
rect 18061 8585 18095 8619
rect 23029 8585 23063 8619
rect 25881 8585 25915 8619
rect 29009 8585 29043 8619
rect 30021 8585 30055 8619
rect 4629 8517 4663 8551
rect 5181 8517 5215 8551
rect 8217 8517 8251 8551
rect 22753 8517 22787 8551
rect 29653 8517 29687 8551
rect 29745 8517 29779 8551
rect 3157 8449 3191 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 6653 8449 6687 8483
rect 10977 8449 11011 8483
rect 11897 8449 11931 8483
rect 14666 8449 14700 8483
rect 15393 8449 15427 8483
rect 17141 8449 17175 8483
rect 18337 8449 18371 8483
rect 18429 8449 18463 8483
rect 18521 8449 18555 8483
rect 18705 8449 18739 8483
rect 19717 8449 19751 8483
rect 22477 8449 22511 8483
rect 22661 8449 22695 8483
rect 22845 8449 22879 8483
rect 25237 8449 25271 8483
rect 25421 8449 25455 8483
rect 25513 8449 25547 8483
rect 25605 8449 25639 8483
rect 27537 8449 27571 8483
rect 27629 8449 27663 8483
rect 27721 8449 27755 8483
rect 27905 8449 27939 8483
rect 28365 8449 28399 8483
rect 28549 8449 28583 8483
rect 28641 8449 28675 8483
rect 28733 8449 28767 8483
rect 29469 8449 29503 8483
rect 29837 8449 29871 8483
rect 34529 8449 34563 8483
rect 34621 8449 34655 8483
rect 34713 8449 34747 8483
rect 34897 8449 34931 8483
rect 3249 8381 3283 8415
rect 3433 8381 3467 8415
rect 6377 8381 6411 8415
rect 11529 8381 11563 8415
rect 12541 8381 12575 8415
rect 14933 8381 14967 8415
rect 19441 8381 19475 8415
rect 20729 8381 20763 8415
rect 1501 8313 1535 8347
rect 1961 8313 1995 8347
rect 3985 8313 4019 8347
rect 8401 8313 8435 8347
rect 10333 8313 10367 8347
rect 17325 8313 17359 8347
rect 24685 8313 24719 8347
rect 27261 8313 27295 8347
rect 33701 8313 33735 8347
rect 2789 8245 2823 8279
rect 5825 8245 5859 8279
rect 11897 8245 11931 8279
rect 26341 8245 26375 8279
rect 34253 8245 34287 8279
rect 3893 8041 3927 8075
rect 13277 8041 13311 8075
rect 16037 8041 16071 8075
rect 17877 8041 17911 8075
rect 18337 8041 18371 8075
rect 22937 8041 22971 8075
rect 28825 8041 28859 8075
rect 34713 8041 34747 8075
rect 14565 7973 14599 8007
rect 34161 7973 34195 8007
rect 2421 7905 2455 7939
rect 5365 7905 5399 7939
rect 5825 7905 5859 7939
rect 6561 7905 6595 7939
rect 11161 7905 11195 7939
rect 12357 7905 12391 7939
rect 12449 7905 12483 7939
rect 32781 7905 32815 7939
rect 2605 7837 2639 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 6101 7837 6135 7871
rect 6929 7837 6963 7871
rect 7021 7837 7055 7871
rect 10793 7837 10827 7871
rect 10977 7837 11011 7871
rect 11069 7837 11103 7871
rect 11345 7837 11379 7871
rect 12173 7837 12207 7871
rect 12541 7837 12575 7871
rect 12725 7837 12759 7871
rect 14749 7837 14783 7871
rect 15301 7837 15335 7871
rect 18521 7837 18555 7871
rect 19441 7837 19475 7871
rect 19533 7837 19567 7871
rect 20085 7837 20119 7871
rect 22385 7837 22419 7871
rect 22569 7837 22603 7871
rect 22753 7837 22787 7871
rect 27445 7837 27479 7871
rect 33048 7837 33082 7871
rect 34897 7837 34931 7871
rect 35081 7837 35115 7871
rect 37197 7837 37231 7871
rect 37360 7837 37394 7871
rect 37473 7837 37507 7871
rect 37611 7837 37645 7871
rect 58173 7837 58207 7871
rect 1961 7769 1995 7803
rect 8309 7769 8343 7803
rect 18705 7769 18739 7803
rect 22661 7769 22695 7803
rect 27712 7769 27746 7803
rect 36737 7769 36771 7803
rect 2789 7701 2823 7735
rect 4445 7701 4479 7735
rect 7205 7701 7239 7735
rect 7757 7701 7791 7735
rect 8953 7701 8987 7735
rect 11529 7701 11563 7735
rect 11989 7701 12023 7735
rect 15485 7701 15519 7735
rect 17233 7701 17267 7735
rect 19257 7701 19291 7735
rect 23489 7701 23523 7735
rect 37841 7701 37875 7735
rect 3801 7497 3835 7531
rect 5825 7497 5859 7531
rect 12173 7497 12207 7531
rect 21281 7497 21315 7531
rect 22753 7497 22787 7531
rect 28365 7497 28399 7531
rect 34437 7497 34471 7531
rect 38761 7497 38795 7531
rect 6469 7429 6503 7463
rect 11621 7429 11655 7463
rect 12725 7429 12759 7463
rect 22385 7429 22419 7463
rect 25513 7429 25547 7463
rect 25697 7429 25731 7463
rect 27077 7429 27111 7463
rect 31033 7429 31067 7463
rect 31493 7429 31527 7463
rect 35725 7429 35759 7463
rect 2421 7361 2455 7395
rect 2688 7361 2722 7395
rect 8318 7361 8352 7395
rect 14473 7361 14507 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 19165 7361 19199 7395
rect 19901 7361 19935 7395
rect 20157 7361 20191 7395
rect 22201 7361 22235 7395
rect 22477 7361 22511 7395
rect 22569 7361 22603 7395
rect 23489 7361 23523 7395
rect 23578 7361 23612 7395
rect 23673 7361 23707 7395
rect 23857 7361 23891 7395
rect 24547 7361 24581 7395
rect 24682 7364 24716 7398
rect 24782 7361 24816 7395
rect 24961 7361 24995 7395
rect 25881 7361 25915 7395
rect 27997 7361 28031 7395
rect 28181 7361 28215 7395
rect 34621 7361 34655 7395
rect 34713 7361 34747 7395
rect 34805 7361 34839 7395
rect 34989 7361 35023 7395
rect 35633 7361 35667 7395
rect 35817 7361 35851 7395
rect 36001 7361 36035 7395
rect 36737 7361 36771 7395
rect 37289 7361 37323 7395
rect 37468 7361 37502 7395
rect 37584 7361 37618 7395
rect 37703 7361 37737 7395
rect 38393 7361 38427 7395
rect 38577 7361 38611 7395
rect 8585 7293 8619 7327
rect 19441 7293 19475 7327
rect 35449 7225 35483 7259
rect 1961 7157 1995 7191
rect 4813 7157 4847 7191
rect 7205 7157 7239 7191
rect 9413 7157 9447 7191
rect 9873 7157 9907 7191
rect 15117 7157 15151 7191
rect 16681 7157 16715 7191
rect 23213 7157 23247 7191
rect 24317 7157 24351 7191
rect 29745 7157 29779 7191
rect 37933 7157 37967 7191
rect 1593 6953 1627 6987
rect 2605 6953 2639 6987
rect 20913 6953 20947 6987
rect 24501 6953 24535 6987
rect 7389 6817 7423 6851
rect 7481 6817 7515 6851
rect 7849 6817 7883 6851
rect 9873 6817 9907 6851
rect 15393 6817 15427 6851
rect 34069 6817 34103 6851
rect 2789 6749 2823 6783
rect 5365 6749 5399 6783
rect 7113 6749 7147 6783
rect 7297 6749 7331 6783
rect 7665 6749 7699 6783
rect 9597 6749 9631 6783
rect 11253 6749 11287 6783
rect 15623 6749 15657 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 16037 6749 16071 6783
rect 18705 6749 18739 6783
rect 22477 6749 22511 6783
rect 22753 6749 22787 6783
rect 26801 6749 26835 6783
rect 27905 6749 27939 6783
rect 30205 6749 30239 6783
rect 35173 6749 35207 6783
rect 36921 6749 36955 6783
rect 37933 6749 37967 6783
rect 38189 6749 38223 6783
rect 8953 6681 8987 6715
rect 11520 6681 11554 6715
rect 14841 6681 14875 6715
rect 16681 6681 16715 6715
rect 16865 6681 16899 6715
rect 18061 6681 18095 6715
rect 19625 6681 19659 6715
rect 28089 6681 28123 6715
rect 30472 6681 30506 6715
rect 2145 6613 2179 6647
rect 3985 6613 4019 6647
rect 4537 6613 4571 6647
rect 6009 6613 6043 6647
rect 6561 6613 6595 6647
rect 8401 6613 8435 6647
rect 12633 6613 12667 6647
rect 16497 6613 16531 6647
rect 18521 6613 18555 6647
rect 25513 6613 25547 6647
rect 27721 6613 27755 6647
rect 31585 6613 31619 6647
rect 39313 6613 39347 6647
rect 3525 6409 3559 6443
rect 4445 6409 4479 6443
rect 8309 6409 8343 6443
rect 16681 6409 16715 6443
rect 19809 6409 19843 6443
rect 24685 6409 24719 6443
rect 28457 6409 28491 6443
rect 30757 6409 30791 6443
rect 33793 6409 33827 6443
rect 39129 6409 39163 6443
rect 1869 6341 1903 6375
rect 12826 6341 12860 6375
rect 17049 6341 17083 6375
rect 22017 6341 22051 6375
rect 22201 6341 22235 6375
rect 29285 6341 29319 6375
rect 29469 6341 29503 6375
rect 37994 6341 38028 6375
rect 2421 6273 2455 6307
rect 2513 6273 2547 6307
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7481 6273 7515 6307
rect 8125 6273 8159 6307
rect 8769 6273 8803 6307
rect 13093 6273 13127 6307
rect 15209 6273 15243 6307
rect 15372 6273 15406 6307
rect 15488 6273 15522 6307
rect 15577 6273 15611 6307
rect 16865 6273 16899 6307
rect 20085 6273 20119 6307
rect 20177 6273 20211 6307
rect 20269 6273 20303 6307
rect 20453 6273 20487 6307
rect 23305 6273 23339 6307
rect 23572 6273 23606 6307
rect 27077 6273 27111 6307
rect 27333 6273 27367 6307
rect 30113 6273 30147 6307
rect 30297 6273 30331 6307
rect 30389 6273 30423 6307
rect 30481 6273 30515 6307
rect 31217 6273 31251 6307
rect 34621 6273 34655 6307
rect 34713 6273 34747 6307
rect 34805 6273 34839 6307
rect 34989 6273 35023 6307
rect 35725 6273 35759 6307
rect 35909 6273 35943 6307
rect 36001 6273 36035 6307
rect 36093 6273 36127 6307
rect 37749 6273 37783 6307
rect 3617 6205 3651 6239
rect 3801 6205 3835 6239
rect 5549 6205 5583 6239
rect 9413 6205 9447 6239
rect 19073 6205 19107 6239
rect 19349 6205 19383 6239
rect 21833 6205 21867 6239
rect 25605 6205 25639 6239
rect 25881 6205 25915 6239
rect 29653 6205 29687 6239
rect 3157 6137 3191 6171
rect 7665 6137 7699 6171
rect 58173 6137 58207 6171
rect 2697 6069 2731 6103
rect 5089 6069 5123 6103
rect 6377 6069 6411 6103
rect 8953 6069 8987 6103
rect 10149 6069 10183 6103
rect 10609 6069 10643 6103
rect 11713 6069 11747 6103
rect 14657 6069 14691 6103
rect 15853 6069 15887 6103
rect 20913 6069 20947 6103
rect 34345 6069 34379 6103
rect 36369 6069 36403 6103
rect 5733 5865 5767 5899
rect 6745 5865 6779 5899
rect 12817 5865 12851 5899
rect 13369 5865 13403 5899
rect 17049 5865 17083 5899
rect 20269 5865 20303 5899
rect 24409 5865 24443 5899
rect 26985 5865 27019 5899
rect 30665 5865 30699 5899
rect 34713 5865 34747 5899
rect 36001 5865 36035 5899
rect 37381 5865 37415 5899
rect 3249 5797 3283 5831
rect 6837 5797 6871 5831
rect 8217 5797 8251 5831
rect 10149 5797 10183 5831
rect 10517 5797 10551 5831
rect 17877 5797 17911 5831
rect 1869 5729 1903 5763
rect 5457 5729 5491 5763
rect 10241 5729 10275 5763
rect 18705 5729 18739 5763
rect 32045 5729 32079 5763
rect 5549 5661 5583 5695
rect 6929 5661 6963 5695
rect 7665 5661 7699 5695
rect 8401 5661 8435 5695
rect 9413 5661 9447 5695
rect 10020 5661 10054 5695
rect 11437 5661 11471 5695
rect 12081 5661 12115 5695
rect 13369 5661 13403 5695
rect 13553 5661 13587 5695
rect 14841 5661 14875 5695
rect 14930 5661 14964 5695
rect 15025 5658 15059 5692
rect 15209 5661 15243 5695
rect 15669 5661 15703 5695
rect 15925 5661 15959 5695
rect 24593 5661 24627 5695
rect 24777 5661 24811 5695
rect 26525 5661 26559 5695
rect 27261 5661 27295 5695
rect 27353 5661 27387 5695
rect 27445 5661 27479 5695
rect 27629 5661 27663 5695
rect 29837 5661 29871 5695
rect 30021 5661 30055 5695
rect 34897 5661 34931 5695
rect 35817 5661 35851 5695
rect 37197 5661 37231 5695
rect 2136 5593 2170 5627
rect 4077 5593 4111 5627
rect 6653 5593 6687 5627
rect 9873 5593 9907 5627
rect 18337 5593 18371 5627
rect 18521 5593 18555 5627
rect 19349 5593 19383 5627
rect 19533 5593 19567 5627
rect 31778 5593 31812 5627
rect 35081 5593 35115 5627
rect 35633 5593 35667 5627
rect 37013 5593 37047 5627
rect 4629 5525 4663 5559
rect 5089 5525 5123 5559
rect 7481 5525 7515 5559
rect 14565 5525 14599 5559
rect 19717 5525 19751 5559
rect 30205 5525 30239 5559
rect 6561 5321 6595 5355
rect 8677 5321 8711 5355
rect 14289 5321 14323 5355
rect 16129 5321 16163 5355
rect 23121 5321 23155 5355
rect 30849 5321 30883 5355
rect 35633 5321 35667 5355
rect 2789 5253 2823 5287
rect 4353 5253 4387 5287
rect 7113 5253 7147 5287
rect 7665 5253 7699 5287
rect 10977 5253 11011 5287
rect 14994 5253 15028 5287
rect 1961 5185 1995 5219
rect 2053 5185 2087 5219
rect 4905 5185 4939 5219
rect 5549 5185 5583 5219
rect 6377 5185 6411 5219
rect 7849 5185 7883 5219
rect 8033 5185 8067 5219
rect 8493 5185 8527 5219
rect 9597 5185 9631 5219
rect 14749 5185 14783 5219
rect 17693 5185 17727 5219
rect 18521 5185 18555 5219
rect 18705 5185 18739 5219
rect 18797 5185 18831 5219
rect 18889 5185 18923 5219
rect 19625 5185 19659 5219
rect 19809 5185 19843 5219
rect 19901 5185 19935 5219
rect 19993 5185 20027 5219
rect 20729 5185 20763 5219
rect 24234 5185 24268 5219
rect 24501 5185 24535 5219
rect 30205 5185 30239 5219
rect 30389 5191 30423 5225
rect 30481 5185 30515 5219
rect 30573 5185 30607 5219
rect 6653 5117 6687 5151
rect 10609 5117 10643 5151
rect 12633 5117 12667 5151
rect 17969 5117 18003 5151
rect 24961 5117 24995 5151
rect 25237 5117 25271 5151
rect 54401 5117 54435 5151
rect 7113 5049 7147 5083
rect 10057 5049 10091 5083
rect 10517 5049 10551 5083
rect 13277 5049 13311 5083
rect 29653 5049 29687 5083
rect 55045 5049 55079 5083
rect 1777 4981 1811 5015
rect 5089 4981 5123 5015
rect 5733 4981 5767 5015
rect 10425 4981 10459 5015
rect 11989 4981 12023 5015
rect 19165 4981 19199 5015
rect 20269 4981 20303 5015
rect 53757 4981 53791 5015
rect 58173 4981 58207 5015
rect 3985 4777 4019 4811
rect 5365 4777 5399 4811
rect 6469 4777 6503 4811
rect 8217 4777 8251 4811
rect 9229 4777 9263 4811
rect 10241 4777 10275 4811
rect 10701 4777 10735 4811
rect 12081 4777 12115 4811
rect 12265 4777 12299 4811
rect 35909 4777 35943 4811
rect 3249 4709 3283 4743
rect 7297 4709 7331 4743
rect 10609 4709 10643 4743
rect 16957 4709 16991 4743
rect 18337 4709 18371 4743
rect 21281 4709 21315 4743
rect 30665 4709 30699 4743
rect 52837 4709 52871 4743
rect 55321 4709 55355 4743
rect 8125 4641 8159 4675
rect 9100 4641 9134 4675
rect 9321 4641 9355 4675
rect 9413 4641 9447 4675
rect 10517 4641 10551 4675
rect 31493 4641 31527 4675
rect 37289 4641 37323 4675
rect 54125 4641 54159 4675
rect 55965 4641 55999 4675
rect 2605 4573 2639 4607
rect 3057 4573 3091 4607
rect 3801 4573 3835 4607
rect 4445 4573 4479 4607
rect 5457 4573 5491 4607
rect 6009 4573 6043 4607
rect 6377 4573 6411 4607
rect 6653 4573 6687 4607
rect 7113 4573 7147 4607
rect 7757 4573 7791 4607
rect 8217 4573 8251 4607
rect 11069 4573 11103 4607
rect 11621 4573 11655 4607
rect 11713 4573 11747 4607
rect 12081 4573 12115 4607
rect 12817 4573 12851 4607
rect 14197 4573 14231 4607
rect 19901 4573 19935 4607
rect 24869 4573 24903 4607
rect 26065 4573 26099 4607
rect 26755 4573 26789 4607
rect 26893 4573 26927 4607
rect 26985 4573 27019 4607
rect 27169 4573 27203 4607
rect 27813 4573 27847 4607
rect 27997 4573 28031 4607
rect 30021 4573 30055 4607
rect 30205 4573 30239 4607
rect 30297 4573 30331 4607
rect 30389 4573 30423 4607
rect 31309 4573 31343 4607
rect 37022 4573 37056 4607
rect 52193 4573 52227 4607
rect 53481 4573 53515 4607
rect 1961 4505 1995 4539
rect 8953 4505 8987 4539
rect 20146 4505 20180 4539
rect 27629 4505 27663 4539
rect 31125 4505 31159 4539
rect 2421 4437 2455 4471
rect 4629 4437 4663 4471
rect 6193 4437 6227 4471
rect 8401 4437 8435 4471
rect 13461 4437 13495 4471
rect 26525 4437 26559 4471
rect 29009 4437 29043 4471
rect 6587 4233 6621 4267
rect 7573 4233 7607 4267
rect 31585 4233 31619 4267
rect 4997 4165 5031 4199
rect 6377 4165 6411 4199
rect 19616 4165 19650 4199
rect 30472 4165 30506 4199
rect 1685 4097 1719 4131
rect 2329 4097 2363 4131
rect 2421 4097 2455 4131
rect 3157 4097 3191 4131
rect 4353 4097 4387 4131
rect 5825 4097 5859 4131
rect 7757 4097 7791 4131
rect 7941 4097 7975 4131
rect 8585 4097 8619 4131
rect 8953 4097 8987 4131
rect 9965 4097 9999 4131
rect 15025 4097 15059 4131
rect 15485 4097 15519 4131
rect 19349 4097 19383 4131
rect 30205 4097 30239 4131
rect 33517 4097 33551 4131
rect 33784 4097 33818 4131
rect 54677 4097 54711 4131
rect 4813 4029 4847 4063
rect 8493 4029 8527 4063
rect 52745 4029 52779 4063
rect 55965 4029 55999 4063
rect 2973 3961 3007 3995
rect 4169 3961 4203 3995
rect 6745 3961 6779 3995
rect 9137 3961 9171 3995
rect 34897 3961 34931 3995
rect 1869 3893 1903 3927
rect 5641 3893 5675 3927
rect 6561 3893 6595 3927
rect 7941 3893 7975 3927
rect 8953 3893 8987 3927
rect 9781 3893 9815 3927
rect 10977 3893 11011 3927
rect 11805 3893 11839 3927
rect 12449 3893 12483 3927
rect 13093 3893 13127 3927
rect 13737 3893 13771 3927
rect 14381 3893 14415 3927
rect 14841 3893 14875 3927
rect 20729 3893 20763 3927
rect 51181 3893 51215 3927
rect 51825 3893 51859 3927
rect 53389 3893 53423 3927
rect 54033 3893 54067 3927
rect 55321 3893 55355 3927
rect 58173 3893 58207 3927
rect 5181 3689 5215 3723
rect 5917 3689 5951 3723
rect 6101 3689 6135 3723
rect 9321 3689 9355 3723
rect 9781 3689 9815 3723
rect 10517 3689 10551 3723
rect 27445 3689 27479 3723
rect 8953 3621 8987 3655
rect 9413 3621 9447 3655
rect 14105 3621 14139 3655
rect 14841 3621 14875 3655
rect 46949 3621 46983 3655
rect 52837 3621 52871 3655
rect 55321 3621 55355 3655
rect 1869 3553 1903 3587
rect 3801 3553 3835 3587
rect 6837 3553 6871 3587
rect 9505 3553 9539 3587
rect 12909 3553 12943 3587
rect 26065 3553 26099 3587
rect 51549 3553 51583 3587
rect 53481 3553 53515 3587
rect 56609 3553 56643 3587
rect 2125 3485 2159 3519
rect 4068 3485 4102 3519
rect 6561 3485 6595 3519
rect 8309 3485 8343 3519
rect 10333 3485 10367 3519
rect 11069 3485 11103 3519
rect 12265 3485 12299 3519
rect 13369 3485 13403 3519
rect 15393 3485 15427 3519
rect 16037 3485 16071 3519
rect 16865 3485 16899 3519
rect 17693 3485 17727 3519
rect 18521 3485 18555 3519
rect 19625 3485 19659 3519
rect 20453 3485 20487 3519
rect 21281 3485 21315 3519
rect 22201 3485 22235 3519
rect 22661 3485 22695 3519
rect 23489 3485 23523 3519
rect 24593 3485 24627 3519
rect 25605 3485 25639 3519
rect 26332 3485 26366 3519
rect 27905 3485 27939 3519
rect 28733 3485 28767 3519
rect 34805 3485 34839 3519
rect 35449 3485 35483 3519
rect 36093 3485 36127 3519
rect 36737 3485 36771 3519
rect 37565 3485 37599 3519
rect 38669 3485 38703 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 41337 3485 41371 3519
rect 42533 3485 42567 3519
rect 43177 3485 43211 3519
rect 45017 3485 45051 3519
rect 45661 3485 45695 3519
rect 46305 3485 46339 3519
rect 47777 3485 47811 3519
rect 48421 3485 48455 3519
rect 50261 3485 50295 3519
rect 50905 3485 50939 3519
rect 52193 3485 52227 3519
rect 54125 3485 54159 3519
rect 55965 3485 55999 3519
rect 57529 3485 57563 3519
rect 58173 3485 58207 3519
rect 5733 3417 5767 3451
rect 5949 3417 5983 3451
rect 14381 3417 14415 3451
rect 14841 3417 14875 3451
rect 3249 3349 3283 3383
rect 8217 3349 8251 3383
rect 11253 3349 11287 3383
rect 13553 3349 13587 3383
rect 14289 3349 14323 3383
rect 1869 3145 1903 3179
rect 12909 3145 12943 3179
rect 3332 3077 3366 3111
rect 9597 3077 9631 3111
rect 10425 3077 10459 3111
rect 10793 3077 10827 3111
rect 1685 3009 1719 3043
rect 2605 3009 2639 3043
rect 4905 3009 4939 3043
rect 5825 3009 5859 3043
rect 7665 3009 7699 3043
rect 8125 3009 8159 3043
rect 9045 3009 9079 3043
rect 9965 3009 9999 3043
rect 11805 3009 11839 3043
rect 12725 3009 12759 3043
rect 54033 3009 54067 3043
rect 54677 3009 54711 3043
rect 55321 3009 55355 3043
rect 3065 2941 3099 2975
rect 7389 2941 7423 2975
rect 8677 2941 8711 2975
rect 16681 2941 16715 2975
rect 18061 2941 18095 2975
rect 19349 2941 19383 2975
rect 25789 2941 25823 2975
rect 33425 2941 33459 2975
rect 39221 2941 39255 2975
rect 43085 2941 43119 2975
rect 55965 2941 55999 2975
rect 56609 2941 56643 2975
rect 8493 2873 8527 2907
rect 11621 2873 11655 2907
rect 14197 2873 14231 2907
rect 34713 2873 34747 2907
rect 37933 2873 37967 2907
rect 39865 2873 39899 2907
rect 41153 2873 41187 2907
rect 43729 2873 43763 2907
rect 45017 2873 45051 2907
rect 45661 2873 45695 2907
rect 48237 2873 48271 2907
rect 49525 2873 49559 2907
rect 50813 2873 50847 2907
rect 52745 2873 52779 2907
rect 57897 2873 57931 2907
rect 2421 2805 2455 2839
rect 4445 2805 4479 2839
rect 5089 2805 5123 2839
rect 5641 2805 5675 2839
rect 8585 2805 8619 2839
rect 13553 2805 13587 2839
rect 14841 2805 14875 2839
rect 15485 2805 15519 2839
rect 16129 2805 16163 2839
rect 17417 2805 17451 2839
rect 18705 2805 18739 2839
rect 19993 2805 20027 2839
rect 20637 2805 20671 2839
rect 21281 2805 21315 2839
rect 22569 2805 22603 2839
rect 23213 2805 23247 2839
rect 23857 2805 23891 2839
rect 24501 2805 24535 2839
rect 25145 2805 25179 2839
rect 26433 2805 26467 2839
rect 27629 2805 27663 2839
rect 28089 2805 28123 2839
rect 28917 2805 28951 2839
rect 29561 2805 29595 2839
rect 30021 2805 30055 2839
rect 30665 2805 30699 2839
rect 32137 2805 32171 2839
rect 32781 2805 32815 2839
rect 34069 2805 34103 2839
rect 35357 2805 35391 2839
rect 36001 2805 36035 2839
rect 37289 2805 37323 2839
rect 38577 2805 38611 2839
rect 40509 2805 40543 2839
rect 42441 2805 42475 2839
rect 44373 2805 44407 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48881 2805 48915 2839
rect 50169 2805 50203 2839
rect 51457 2805 51491 2839
rect 53389 2805 53423 2839
rect 1777 2601 1811 2635
rect 5595 2601 5629 2635
rect 6653 2601 6687 2635
rect 12449 2601 12483 2635
rect 13553 2601 13587 2635
rect 19993 2601 20027 2635
rect 55321 2601 55355 2635
rect 2329 2533 2363 2567
rect 10793 2533 10827 2567
rect 11621 2533 11655 2567
rect 14841 2533 14875 2567
rect 27721 2533 27755 2567
rect 36001 2533 36035 2567
rect 39865 2533 39899 2567
rect 43729 2533 43763 2567
rect 47593 2533 47627 2567
rect 51457 2533 51491 2567
rect 54033 2533 54067 2567
rect 7573 2465 7607 2499
rect 15485 2465 15519 2499
rect 17417 2465 17451 2499
rect 18705 2465 18739 2499
rect 20637 2465 20671 2499
rect 23857 2465 23891 2499
rect 25789 2465 25823 2499
rect 32781 2465 32815 2499
rect 34713 2465 34747 2499
rect 37289 2465 37323 2499
rect 40509 2465 40543 2499
rect 42441 2465 42475 2499
rect 45017 2465 45051 2499
rect 48237 2465 48271 2499
rect 50169 2465 50203 2499
rect 52745 2465 52779 2499
rect 57897 2465 57931 2499
rect 1593 2397 1627 2431
rect 2513 2397 2547 2431
rect 2973 2397 3007 2431
rect 4537 2397 4571 2431
rect 5825 2397 5859 2431
rect 7297 2397 7331 2431
rect 8953 2397 8987 2431
rect 10609 2397 10643 2431
rect 11805 2397 11839 2431
rect 12265 2397 12299 2431
rect 13369 2397 13403 2431
rect 16129 2397 16163 2431
rect 18061 2397 18095 2431
rect 21281 2397 21315 2431
rect 22569 2397 22603 2431
rect 23213 2397 23247 2431
rect 25145 2397 25179 2431
rect 26433 2397 26467 2431
rect 28365 2397 28399 2431
rect 29009 2397 29043 2431
rect 30113 2397 30147 2431
rect 30757 2397 30791 2431
rect 31217 2397 31251 2431
rect 32137 2397 32171 2431
rect 33425 2397 33459 2431
rect 35357 2397 35391 2431
rect 37933 2397 37967 2431
rect 38577 2397 38611 2431
rect 41153 2397 41187 2431
rect 43085 2397 43119 2431
rect 45661 2397 45695 2431
rect 46305 2397 46339 2431
rect 48881 2397 48915 2431
rect 50813 2397 50847 2431
rect 53389 2397 53423 2431
rect 55965 2397 55999 2431
rect 56609 2397 56643 2431
rect 6745 2329 6779 2363
rect 9781 2329 9815 2363
rect 3157 2261 3191 2295
rect 4353 2261 4387 2295
rect 9137 2261 9171 2295
rect 9873 2261 9907 2295
rect 14197 2261 14231 2295
rect 16681 2261 16715 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 1762 57400 1768 57452
rect 1820 57440 1826 57452
rect 1857 57443 1915 57449
rect 1857 57440 1869 57443
rect 1820 57412 1869 57440
rect 1820 57400 1826 57412
rect 1857 57409 1869 57412
rect 1903 57409 1915 57443
rect 1857 57403 1915 57409
rect 3326 57400 3332 57452
rect 3384 57440 3390 57452
rect 3789 57443 3847 57449
rect 3789 57440 3801 57443
rect 3384 57412 3801 57440
rect 3384 57400 3390 57412
rect 3789 57409 3801 57412
rect 3835 57409 3847 57443
rect 3789 57403 3847 57409
rect 4890 57400 4896 57452
rect 4948 57440 4954 57452
rect 4985 57443 5043 57449
rect 4985 57440 4997 57443
rect 4948 57412 4997 57440
rect 4948 57400 4954 57412
rect 4985 57409 4997 57412
rect 5031 57409 5043 57443
rect 4985 57403 5043 57409
rect 6454 57400 6460 57452
rect 6512 57440 6518 57452
rect 6549 57443 6607 57449
rect 6549 57440 6561 57443
rect 6512 57412 6561 57440
rect 6512 57400 6518 57412
rect 6549 57409 6561 57412
rect 6595 57409 6607 57443
rect 6549 57403 6607 57409
rect 8018 57400 8024 57452
rect 8076 57440 8082 57452
rect 8113 57443 8171 57449
rect 8113 57440 8125 57443
rect 8076 57412 8125 57440
rect 8076 57400 8082 57412
rect 8113 57409 8125 57412
rect 8159 57409 8171 57443
rect 9674 57440 9680 57452
rect 9635 57412 9680 57440
rect 8113 57403 8171 57409
rect 9674 57400 9680 57412
rect 9732 57400 9738 57452
rect 11146 57400 11152 57452
rect 11204 57440 11210 57452
rect 11517 57443 11575 57449
rect 11517 57440 11529 57443
rect 11204 57412 11529 57440
rect 11204 57400 11210 57412
rect 11517 57409 11529 57412
rect 11563 57409 11575 57443
rect 11517 57403 11575 57409
rect 12710 57400 12716 57452
rect 12768 57440 12774 57452
rect 12805 57443 12863 57449
rect 12805 57440 12817 57443
rect 12768 57412 12817 57440
rect 12768 57400 12774 57412
rect 12805 57409 12817 57412
rect 12851 57409 12863 57443
rect 12805 57403 12863 57409
rect 14274 57400 14280 57452
rect 14332 57440 14338 57452
rect 14369 57443 14427 57449
rect 14369 57440 14381 57443
rect 14332 57412 14381 57440
rect 14332 57400 14338 57412
rect 14369 57409 14381 57412
rect 14415 57409 14427 57443
rect 14369 57403 14427 57409
rect 15838 57400 15844 57452
rect 15896 57440 15902 57452
rect 15933 57443 15991 57449
rect 15933 57440 15945 57443
rect 15896 57412 15945 57440
rect 15896 57400 15902 57412
rect 15933 57409 15945 57412
rect 15979 57409 15991 57443
rect 15933 57403 15991 57409
rect 17402 57400 17408 57452
rect 17460 57440 17466 57452
rect 17497 57443 17555 57449
rect 17497 57440 17509 57443
rect 17460 57412 17509 57440
rect 17460 57400 17466 57412
rect 17497 57409 17509 57412
rect 17543 57409 17555 57443
rect 17497 57403 17555 57409
rect 18966 57400 18972 57452
rect 19024 57440 19030 57452
rect 19245 57443 19303 57449
rect 19245 57440 19257 57443
rect 19024 57412 19257 57440
rect 19024 57400 19030 57412
rect 19245 57409 19257 57412
rect 19291 57409 19303 57443
rect 19245 57403 19303 57409
rect 20530 57400 20536 57452
rect 20588 57440 20594 57452
rect 20625 57443 20683 57449
rect 20625 57440 20637 57443
rect 20588 57412 20637 57440
rect 20588 57400 20594 57412
rect 20625 57409 20637 57412
rect 20671 57409 20683 57443
rect 20625 57403 20683 57409
rect 22094 57400 22100 57452
rect 22152 57440 22158 57452
rect 22189 57443 22247 57449
rect 22189 57440 22201 57443
rect 22152 57412 22201 57440
rect 22152 57400 22158 57412
rect 22189 57409 22201 57412
rect 22235 57409 22247 57443
rect 22189 57403 22247 57409
rect 23658 57400 23664 57452
rect 23716 57440 23722 57452
rect 24397 57443 24455 57449
rect 24397 57440 24409 57443
rect 23716 57412 24409 57440
rect 23716 57400 23722 57412
rect 24397 57409 24409 57412
rect 24443 57409 24455 57443
rect 24397 57403 24455 57409
rect 25222 57400 25228 57452
rect 25280 57440 25286 57452
rect 25317 57443 25375 57449
rect 25317 57440 25329 57443
rect 25280 57412 25329 57440
rect 25280 57400 25286 57412
rect 25317 57409 25329 57412
rect 25363 57409 25375 57443
rect 25317 57403 25375 57409
rect 26786 57400 26792 57452
rect 26844 57440 26850 57452
rect 26973 57443 27031 57449
rect 26973 57440 26985 57443
rect 26844 57412 26985 57440
rect 26844 57400 26850 57412
rect 26973 57409 26985 57412
rect 27019 57409 27031 57443
rect 26973 57403 27031 57409
rect 28350 57400 28356 57452
rect 28408 57440 28414 57452
rect 28445 57443 28503 57449
rect 28445 57440 28457 57443
rect 28408 57412 28457 57440
rect 28408 57400 28414 57412
rect 28445 57409 28457 57412
rect 28491 57409 28503 57443
rect 28445 57403 28503 57409
rect 29914 57400 29920 57452
rect 29972 57440 29978 57452
rect 30009 57443 30067 57449
rect 30009 57440 30021 57443
rect 29972 57412 30021 57440
rect 29972 57400 29978 57412
rect 30009 57409 30021 57412
rect 30055 57409 30067 57443
rect 30009 57403 30067 57409
rect 31478 57400 31484 57452
rect 31536 57440 31542 57452
rect 32125 57443 32183 57449
rect 32125 57440 32137 57443
rect 31536 57412 32137 57440
rect 31536 57400 31542 57412
rect 32125 57409 32137 57412
rect 32171 57409 32183 57443
rect 33134 57440 33140 57452
rect 33095 57412 33140 57440
rect 32125 57403 32183 57409
rect 33134 57400 33140 57412
rect 33192 57400 33198 57452
rect 34606 57400 34612 57452
rect 34664 57440 34670 57452
rect 34701 57443 34759 57449
rect 34701 57440 34713 57443
rect 34664 57412 34713 57440
rect 34664 57400 34670 57412
rect 34701 57409 34713 57412
rect 34747 57409 34759 57443
rect 34701 57403 34759 57409
rect 36170 57400 36176 57452
rect 36228 57440 36234 57452
rect 36265 57443 36323 57449
rect 36265 57440 36277 57443
rect 36228 57412 36277 57440
rect 36228 57400 36234 57412
rect 36265 57409 36277 57412
rect 36311 57409 36323 57443
rect 36265 57403 36323 57409
rect 37734 57400 37740 57452
rect 37792 57440 37798 57452
rect 37829 57443 37887 57449
rect 37829 57440 37841 57443
rect 37792 57412 37841 57440
rect 37792 57400 37798 57412
rect 37829 57409 37841 57412
rect 37875 57409 37887 57443
rect 37829 57403 37887 57409
rect 39298 57400 39304 57452
rect 39356 57440 39362 57452
rect 39853 57443 39911 57449
rect 39853 57440 39865 57443
rect 39356 57412 39865 57440
rect 39356 57400 39362 57412
rect 39853 57409 39865 57412
rect 39899 57409 39911 57443
rect 39853 57403 39911 57409
rect 40862 57400 40868 57452
rect 40920 57440 40926 57452
rect 40957 57443 41015 57449
rect 40957 57440 40969 57443
rect 40920 57412 40969 57440
rect 40920 57400 40926 57412
rect 40957 57409 40969 57412
rect 41003 57409 41015 57443
rect 40957 57403 41015 57409
rect 42426 57400 42432 57452
rect 42484 57440 42490 57452
rect 42521 57443 42579 57449
rect 42521 57440 42533 57443
rect 42484 57412 42533 57440
rect 42484 57400 42490 57412
rect 42521 57409 42533 57412
rect 42567 57409 42579 57443
rect 42521 57403 42579 57409
rect 43990 57400 43996 57452
rect 44048 57440 44054 57452
rect 44085 57443 44143 57449
rect 44085 57440 44097 57443
rect 44048 57412 44097 57440
rect 44048 57400 44054 57412
rect 44085 57409 44097 57412
rect 44131 57409 44143 57443
rect 44085 57403 44143 57409
rect 45554 57400 45560 57452
rect 45612 57440 45618 57452
rect 45649 57443 45707 57449
rect 45649 57440 45661 57443
rect 45612 57412 45661 57440
rect 45612 57400 45618 57412
rect 45649 57409 45661 57412
rect 45695 57409 45707 57443
rect 45649 57403 45707 57409
rect 47118 57400 47124 57452
rect 47176 57440 47182 57452
rect 47581 57443 47639 57449
rect 47581 57440 47593 57443
rect 47176 57412 47593 57440
rect 47176 57400 47182 57412
rect 47581 57409 47593 57412
rect 47627 57409 47639 57443
rect 47581 57403 47639 57409
rect 48682 57400 48688 57452
rect 48740 57440 48746 57452
rect 48777 57443 48835 57449
rect 48777 57440 48789 57443
rect 48740 57412 48789 57440
rect 48740 57400 48746 57412
rect 48777 57409 48789 57412
rect 48823 57409 48835 57443
rect 48777 57403 48835 57409
rect 50154 57400 50160 57452
rect 50212 57440 50218 57452
rect 50341 57443 50399 57449
rect 50341 57440 50353 57443
rect 50212 57412 50353 57440
rect 50212 57400 50218 57412
rect 50341 57409 50353 57412
rect 50387 57409 50399 57443
rect 50341 57403 50399 57409
rect 51810 57400 51816 57452
rect 51868 57440 51874 57452
rect 51905 57443 51963 57449
rect 51905 57440 51917 57443
rect 51868 57412 51917 57440
rect 51868 57400 51874 57412
rect 51905 57409 51917 57412
rect 51951 57409 51963 57443
rect 51905 57403 51963 57409
rect 53374 57400 53380 57452
rect 53432 57440 53438 57452
rect 53469 57443 53527 57449
rect 53469 57440 53481 57443
rect 53432 57412 53481 57440
rect 53432 57400 53438 57412
rect 53469 57409 53481 57412
rect 53515 57409 53527 57443
rect 56594 57440 56600 57452
rect 56555 57412 56600 57440
rect 53469 57403 53527 57409
rect 56594 57400 56600 57412
rect 56652 57400 56658 57452
rect 57977 57443 58035 57449
rect 57977 57409 57989 57443
rect 58023 57440 58035 57443
rect 58066 57440 58072 57452
rect 58023 57412 58072 57440
rect 58023 57409 58035 57412
rect 57977 57403 58035 57409
rect 58066 57400 58072 57412
rect 58124 57400 58130 57452
rect 54938 57332 54944 57384
rect 54996 57372 55002 57384
rect 55309 57375 55367 57381
rect 55309 57372 55321 57375
rect 54996 57344 55321 57372
rect 54996 57332 55002 57344
rect 55309 57341 55321 57344
rect 55355 57341 55367 57375
rect 55309 57335 55367 57341
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 57514 57032 57520 57044
rect 57475 57004 57520 57032
rect 57514 56992 57520 57004
rect 57572 56992 57578 57044
rect 57882 56788 57888 56840
rect 57940 56828 57946 56840
rect 58161 56831 58219 56837
rect 58161 56828 58173 56831
rect 57940 56800 58173 56828
rect 57940 56788 57946 56800
rect 58161 56797 58173 56800
rect 58207 56797 58219 56831
rect 58161 56791 58219 56797
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 58161 56355 58219 56361
rect 58161 56321 58173 56355
rect 58207 56352 58219 56355
rect 58434 56352 58440 56364
rect 58207 56324 58440 56352
rect 58207 56321 58219 56324
rect 58161 56315 58219 56321
rect 58434 56312 58440 56324
rect 58492 56312 58498 56364
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 58158 55128 58164 55140
rect 58119 55100 58164 55128
rect 58158 55088 58164 55100
rect 58216 55088 58222 55140
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 57882 53932 57888 53984
rect 57940 53972 57946 53984
rect 58161 53975 58219 53981
rect 58161 53972 58173 53975
rect 57940 53944 58173 53972
rect 57940 53932 57946 53944
rect 58161 53941 58173 53944
rect 58207 53941 58219 53975
rect 58161 53935 58219 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 57882 52436 57888 52488
rect 57940 52476 57946 52488
rect 58161 52479 58219 52485
rect 58161 52476 58173 52479
rect 57940 52448 58173 52476
rect 57940 52436 57946 52448
rect 58161 52445 58173 52448
rect 58207 52445 58219 52479
rect 58161 52439 58219 52445
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 58158 51388 58164 51400
rect 58119 51360 58164 51388
rect 58158 51348 58164 51360
rect 58216 51348 58222 51400
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 58158 49756 58164 49768
rect 58119 49728 58164 49756
rect 58158 49716 58164 49728
rect 58216 49716 58222 49768
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 58158 48532 58164 48544
rect 58119 48504 58164 48532
rect 58158 48492 58164 48504
rect 58216 48492 58222 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58158 47036 58164 47048
rect 58119 47008 58164 47036
rect 58158 46996 58164 47008
rect 58216 46996 58222 47048
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 58158 45948 58164 45960
rect 58119 45920 58164 45948
rect 58158 45908 58164 45920
rect 58216 45908 58222 45960
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 58158 44248 58164 44260
rect 58119 44220 58164 44248
rect 58158 44208 58164 44220
rect 58216 44208 58222 44260
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 58158 43092 58164 43104
rect 58119 43064 58164 43092
rect 58158 43052 58164 43064
rect 58216 43052 58222 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 12710 42644 12716 42696
rect 12768 42684 12774 42696
rect 13265 42687 13323 42693
rect 13265 42684 13277 42687
rect 12768 42656 13277 42684
rect 12768 42644 12774 42656
rect 13265 42653 13277 42656
rect 13311 42684 13323 42687
rect 20438 42684 20444 42696
rect 13311 42656 20444 42684
rect 13311 42653 13323 42656
rect 13265 42647 13323 42653
rect 20438 42644 20444 42656
rect 20496 42644 20502 42696
rect 14642 42576 14648 42628
rect 14700 42616 14706 42628
rect 15473 42619 15531 42625
rect 15473 42616 15485 42619
rect 14700 42588 15485 42616
rect 14700 42576 14706 42588
rect 15473 42585 15485 42588
rect 15519 42585 15531 42619
rect 15473 42579 15531 42585
rect 15657 42619 15715 42625
rect 15657 42585 15669 42619
rect 15703 42616 15715 42619
rect 16298 42616 16304 42628
rect 15703 42588 16304 42616
rect 15703 42585 15715 42588
rect 15657 42579 15715 42585
rect 16298 42576 16304 42588
rect 16356 42576 16362 42628
rect 14918 42548 14924 42560
rect 14879 42520 14924 42548
rect 14918 42508 14924 42520
rect 14976 42508 14982 42560
rect 15841 42551 15899 42557
rect 15841 42517 15853 42551
rect 15887 42548 15899 42551
rect 15930 42548 15936 42560
rect 15887 42520 15936 42548
rect 15887 42517 15899 42520
rect 15841 42511 15899 42517
rect 15930 42508 15936 42520
rect 15988 42508 15994 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 12158 42304 12164 42356
rect 12216 42344 12222 42356
rect 12216 42316 13860 42344
rect 12216 42304 12222 42316
rect 13832 42285 13860 42316
rect 13817 42279 13875 42285
rect 13817 42245 13829 42279
rect 13863 42276 13875 42279
rect 14642 42276 14648 42288
rect 13863 42248 14648 42276
rect 13863 42245 13875 42248
rect 13817 42239 13875 42245
rect 14642 42236 14648 42248
rect 14700 42236 14706 42288
rect 12710 42208 12716 42220
rect 12671 42180 12716 42208
rect 12710 42168 12716 42180
rect 12768 42168 12774 42220
rect 12802 42211 12860 42217
rect 12802 42177 12814 42211
rect 12848 42177 12860 42211
rect 12802 42171 12860 42177
rect 12820 42140 12848 42171
rect 12894 42168 12900 42220
rect 12952 42217 12958 42220
rect 12952 42208 12960 42217
rect 13081 42211 13139 42217
rect 12952 42180 12997 42208
rect 12952 42171 12960 42180
rect 13081 42177 13093 42211
rect 13127 42177 13139 42211
rect 13081 42171 13139 42177
rect 12952 42168 12958 42171
rect 12728 42112 12848 42140
rect 12728 42084 12756 42112
rect 12710 42032 12716 42084
rect 12768 42032 12774 42084
rect 12986 42032 12992 42084
rect 13044 42072 13050 42084
rect 13096 42072 13124 42171
rect 13906 42168 13912 42220
rect 13964 42208 13970 42220
rect 14001 42211 14059 42217
rect 14001 42208 14013 42211
rect 13964 42180 14013 42208
rect 13964 42168 13970 42180
rect 14001 42177 14013 42180
rect 14047 42177 14059 42211
rect 14001 42171 14059 42177
rect 14829 42211 14887 42217
rect 14829 42177 14841 42211
rect 14875 42208 14887 42211
rect 15378 42208 15384 42220
rect 14875 42180 15384 42208
rect 14875 42177 14887 42180
rect 14829 42171 14887 42177
rect 15378 42168 15384 42180
rect 15436 42168 15442 42220
rect 15470 42168 15476 42220
rect 15528 42208 15534 42220
rect 15657 42211 15715 42217
rect 15528 42180 15573 42208
rect 15528 42168 15534 42180
rect 15657 42177 15669 42211
rect 15703 42177 15715 42211
rect 15657 42171 15715 42177
rect 15013 42143 15071 42149
rect 15013 42109 15025 42143
rect 15059 42140 15071 42143
rect 15672 42140 15700 42171
rect 15746 42168 15752 42220
rect 15804 42208 15810 42220
rect 15887 42211 15945 42217
rect 15804 42180 15849 42208
rect 15804 42168 15810 42180
rect 15887 42177 15899 42211
rect 15933 42208 15945 42211
rect 15933 42180 16574 42208
rect 15933 42177 15945 42180
rect 15887 42171 15945 42177
rect 15059 42112 15700 42140
rect 15059 42109 15071 42112
rect 15013 42103 15071 42109
rect 15470 42072 15476 42084
rect 13044 42044 15476 42072
rect 13044 42032 13050 42044
rect 15470 42032 15476 42044
rect 15528 42032 15534 42084
rect 11977 42007 12035 42013
rect 11977 41973 11989 42007
rect 12023 42004 12035 42007
rect 12066 42004 12072 42016
rect 12023 41976 12072 42004
rect 12023 41973 12035 41976
rect 11977 41967 12035 41973
rect 12066 41964 12072 41976
rect 12124 41964 12130 42016
rect 12434 41964 12440 42016
rect 12492 42004 12498 42016
rect 14185 42007 14243 42013
rect 12492 41976 12537 42004
rect 12492 41964 12498 41976
rect 14185 41973 14197 42007
rect 14231 42004 14243 42007
rect 14550 42004 14556 42016
rect 14231 41976 14556 42004
rect 14231 41973 14243 41976
rect 14185 41967 14243 41973
rect 14550 41964 14556 41976
rect 14608 41964 14614 42016
rect 16114 42004 16120 42016
rect 16075 41976 16120 42004
rect 16114 41964 16120 41976
rect 16172 41964 16178 42016
rect 16546 42004 16574 42180
rect 18601 42143 18659 42149
rect 18601 42109 18613 42143
rect 18647 42140 18659 42143
rect 19886 42140 19892 42152
rect 18647 42112 19892 42140
rect 18647 42109 18659 42112
rect 18601 42103 18659 42109
rect 19886 42100 19892 42112
rect 19944 42100 19950 42152
rect 16761 42007 16819 42013
rect 16761 42004 16773 42007
rect 16546 41976 16773 42004
rect 16761 41973 16773 41976
rect 16807 42004 16819 42007
rect 19518 42004 19524 42016
rect 16807 41976 19524 42004
rect 16807 41973 16819 41976
rect 16761 41967 16819 41973
rect 19518 41964 19524 41976
rect 19576 42004 19582 42016
rect 20073 42007 20131 42013
rect 20073 42004 20085 42007
rect 19576 41976 20085 42004
rect 19576 41964 19582 41976
rect 20073 41973 20085 41976
rect 20119 42004 20131 42007
rect 24762 42004 24768 42016
rect 20119 41976 24768 42004
rect 20119 41973 20131 41976
rect 20073 41967 20131 41973
rect 24762 41964 24768 41976
rect 24820 41964 24826 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 11609 41803 11667 41809
rect 11609 41769 11621 41803
rect 11655 41800 11667 41803
rect 12894 41800 12900 41812
rect 11655 41772 12900 41800
rect 11655 41769 11667 41772
rect 11609 41763 11667 41769
rect 12894 41760 12900 41772
rect 12952 41760 12958 41812
rect 15378 41760 15384 41812
rect 15436 41800 15442 41812
rect 15473 41803 15531 41809
rect 15473 41800 15485 41803
rect 15436 41772 15485 41800
rect 15436 41760 15442 41772
rect 15473 41769 15485 41772
rect 15519 41769 15531 41803
rect 20346 41800 20352 41812
rect 15473 41763 15531 41769
rect 16960 41772 20352 41800
rect 12710 41624 12716 41676
rect 12768 41664 12774 41676
rect 15746 41664 15752 41676
rect 12768 41636 15752 41664
rect 12768 41624 12774 41636
rect 12066 41596 12072 41608
rect 12027 41568 12072 41596
rect 12066 41556 12072 41568
rect 12124 41556 12130 41608
rect 12345 41599 12403 41605
rect 12345 41565 12357 41599
rect 12391 41596 12403 41599
rect 12986 41596 12992 41608
rect 12391 41568 12992 41596
rect 12391 41565 12403 41568
rect 12345 41559 12403 41565
rect 12986 41556 12992 41568
rect 13044 41556 13050 41608
rect 14476 41605 14504 41636
rect 15746 41624 15752 41636
rect 15804 41624 15810 41676
rect 14369 41599 14427 41605
rect 14369 41565 14381 41599
rect 14415 41565 14427 41599
rect 14369 41559 14427 41565
rect 14461 41599 14519 41605
rect 14461 41565 14473 41599
rect 14507 41565 14519 41599
rect 14461 41559 14519 41565
rect 11238 41528 11244 41540
rect 11199 41500 11244 41528
rect 11238 41488 11244 41500
rect 11296 41488 11302 41540
rect 11422 41528 11428 41540
rect 11383 41500 11428 41528
rect 11422 41488 11428 41500
rect 11480 41488 11486 41540
rect 14384 41528 14412 41559
rect 14550 41556 14556 41608
rect 14608 41596 14614 41608
rect 14737 41599 14795 41605
rect 14608 41568 14653 41596
rect 14608 41556 14614 41568
rect 14737 41565 14749 41599
rect 14783 41596 14795 41599
rect 15470 41596 15476 41608
rect 14783 41568 15476 41596
rect 14783 41565 14795 41568
rect 14737 41559 14795 41565
rect 15470 41556 15476 41568
rect 15528 41556 15534 41608
rect 16114 41556 16120 41608
rect 16172 41596 16178 41608
rect 16586 41599 16644 41605
rect 16586 41596 16598 41599
rect 16172 41568 16598 41596
rect 16172 41556 16178 41568
rect 16586 41565 16598 41568
rect 16632 41565 16644 41599
rect 16850 41596 16856 41608
rect 16811 41568 16856 41596
rect 16586 41559 16644 41565
rect 16850 41556 16856 41568
rect 16908 41556 16914 41608
rect 14918 41528 14924 41540
rect 14384 41500 14924 41528
rect 14918 41488 14924 41500
rect 14976 41528 14982 41540
rect 16960 41528 16988 41772
rect 20346 41760 20352 41772
rect 20404 41760 20410 41812
rect 18693 41735 18751 41741
rect 18693 41701 18705 41735
rect 18739 41701 18751 41735
rect 18693 41695 18751 41701
rect 18708 41664 18736 41695
rect 18708 41636 19748 41664
rect 18509 41599 18567 41605
rect 18509 41565 18521 41599
rect 18555 41596 18567 41599
rect 18690 41596 18696 41608
rect 18555 41568 18696 41596
rect 18555 41565 18567 41568
rect 18509 41559 18567 41565
rect 18690 41556 18696 41568
rect 18748 41556 18754 41608
rect 19518 41596 19524 41608
rect 19479 41568 19524 41596
rect 19518 41556 19524 41568
rect 19576 41556 19582 41608
rect 19720 41605 19748 41636
rect 19613 41599 19671 41605
rect 19613 41565 19625 41599
rect 19659 41565 19671 41599
rect 19613 41559 19671 41565
rect 19705 41599 19763 41605
rect 19705 41565 19717 41599
rect 19751 41565 19763 41599
rect 19886 41596 19892 41608
rect 19847 41568 19892 41596
rect 19705 41559 19763 41565
rect 14976 41500 16988 41528
rect 18325 41531 18383 41537
rect 14976 41488 14982 41500
rect 18325 41497 18337 41531
rect 18371 41528 18383 41531
rect 18966 41528 18972 41540
rect 18371 41500 18972 41528
rect 18371 41497 18383 41500
rect 18325 41491 18383 41497
rect 18966 41488 18972 41500
rect 19024 41488 19030 41540
rect 19334 41488 19340 41540
rect 19392 41528 19398 41540
rect 19628 41528 19656 41559
rect 19886 41556 19892 41568
rect 19944 41596 19950 41608
rect 20349 41599 20407 41605
rect 20349 41596 20361 41599
rect 19944 41568 20361 41596
rect 19944 41556 19950 41568
rect 20349 41565 20361 41568
rect 20395 41565 20407 41599
rect 58158 41596 58164 41608
rect 58119 41568 58164 41596
rect 20349 41559 20407 41565
rect 58158 41556 58164 41568
rect 58216 41556 58222 41608
rect 19392 41500 19656 41528
rect 19392 41488 19398 41500
rect 5166 41460 5172 41472
rect 5127 41432 5172 41460
rect 5166 41420 5172 41432
rect 5224 41420 5230 41472
rect 14090 41460 14096 41472
rect 14051 41432 14096 41460
rect 14090 41420 14096 41432
rect 14148 41420 14154 41472
rect 17865 41463 17923 41469
rect 17865 41429 17877 41463
rect 17911 41460 17923 41463
rect 17954 41460 17960 41472
rect 17911 41432 17960 41460
rect 17911 41429 17923 41432
rect 17865 41423 17923 41429
rect 17954 41420 17960 41432
rect 18012 41420 18018 41472
rect 19245 41463 19303 41469
rect 19245 41429 19257 41463
rect 19291 41460 19303 41463
rect 19426 41460 19432 41472
rect 19291 41432 19432 41460
rect 19291 41429 19303 41432
rect 19245 41423 19303 41429
rect 19426 41420 19432 41432
rect 19484 41420 19490 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 12526 41256 12532 41268
rect 10796 41228 12532 41256
rect 5353 41191 5411 41197
rect 5353 41157 5365 41191
rect 5399 41188 5411 41191
rect 6362 41188 6368 41200
rect 5399 41160 6368 41188
rect 5399 41157 5411 41160
rect 5353 41151 5411 41157
rect 6362 41148 6368 41160
rect 6420 41148 6426 41200
rect 10796 41197 10824 41228
rect 12526 41216 12532 41228
rect 12584 41216 12590 41268
rect 15746 41216 15752 41268
rect 15804 41256 15810 41268
rect 16761 41259 16819 41265
rect 15804 41228 15884 41256
rect 15804 41216 15810 41228
rect 7000 41191 7058 41197
rect 7000 41157 7012 41191
rect 7046 41188 7058 41191
rect 8849 41191 8907 41197
rect 8849 41188 8861 41191
rect 7046 41160 8861 41188
rect 7046 41157 7058 41160
rect 7000 41151 7058 41157
rect 8849 41157 8861 41160
rect 8895 41157 8907 41191
rect 8849 41151 8907 41157
rect 10781 41191 10839 41197
rect 10781 41157 10793 41191
rect 10827 41157 10839 41191
rect 10781 41151 10839 41157
rect 10965 41191 11023 41197
rect 10965 41157 10977 41191
rect 11011 41188 11023 41191
rect 11238 41188 11244 41200
rect 11011 41160 11244 41188
rect 11011 41157 11023 41160
rect 10965 41151 11023 41157
rect 11238 41148 11244 41160
rect 11296 41188 11302 41200
rect 12158 41188 12164 41200
rect 11296 41160 12164 41188
rect 11296 41148 11302 41160
rect 12158 41148 12164 41160
rect 12216 41148 12222 41200
rect 12434 41148 12440 41200
rect 12492 41188 12498 41200
rect 12630 41191 12688 41197
rect 12630 41188 12642 41191
rect 12492 41160 12642 41188
rect 12492 41148 12498 41160
rect 12630 41157 12642 41160
rect 12676 41157 12688 41191
rect 12630 41151 12688 41157
rect 14090 41148 14096 41200
rect 14148 41188 14154 41200
rect 14746 41191 14804 41197
rect 14746 41188 14758 41191
rect 14148 41160 14758 41188
rect 14148 41148 14154 41160
rect 14746 41157 14758 41160
rect 14792 41157 14804 41191
rect 14746 41151 14804 41157
rect 5537 41123 5595 41129
rect 5537 41089 5549 41123
rect 5583 41120 5595 41123
rect 5994 41120 6000 41132
rect 5583 41092 6000 41120
rect 5583 41089 5595 41092
rect 5537 41083 5595 41089
rect 5994 41080 6000 41092
rect 6052 41080 6058 41132
rect 9125 41123 9183 41129
rect 9125 41089 9137 41123
rect 9171 41089 9183 41123
rect 9125 41083 9183 41089
rect 9217 41123 9275 41129
rect 9217 41089 9229 41123
rect 9263 41089 9275 41123
rect 9217 41083 9275 41089
rect 6733 41055 6791 41061
rect 6733 41021 6745 41055
rect 6779 41021 6791 41055
rect 6733 41015 6791 41021
rect 4614 40876 4620 40928
rect 4672 40916 4678 40928
rect 5169 40919 5227 40925
rect 5169 40916 5181 40919
rect 4672 40888 5181 40916
rect 4672 40876 4678 40888
rect 5169 40885 5181 40888
rect 5215 40885 5227 40919
rect 6748 40916 6776 41015
rect 9140 40984 9168 41083
rect 9232 41052 9260 41083
rect 9306 41080 9312 41132
rect 9364 41120 9370 41132
rect 9493 41123 9551 41129
rect 9364 41092 9409 41120
rect 9364 41080 9370 41092
rect 9493 41089 9505 41123
rect 9539 41120 9551 41123
rect 10134 41120 10140 41132
rect 9539 41092 10140 41120
rect 9539 41089 9551 41092
rect 9493 41083 9551 41089
rect 10134 41080 10140 41092
rect 10192 41080 10198 41132
rect 14918 41080 14924 41132
rect 14976 41120 14982 41132
rect 15856 41129 15884 41228
rect 16761 41225 16773 41259
rect 16807 41256 16819 41259
rect 17954 41256 17960 41268
rect 16807 41228 17960 41256
rect 16807 41225 16819 41228
rect 16761 41219 16819 41225
rect 15013 41123 15071 41129
rect 15013 41120 15025 41123
rect 14976 41092 15025 41120
rect 14976 41080 14982 41092
rect 15013 41089 15025 41092
rect 15059 41089 15071 41123
rect 15013 41083 15071 41089
rect 15703 41123 15761 41129
rect 15703 41089 15715 41123
rect 15749 41120 15761 41123
rect 15841 41123 15899 41129
rect 15749 41089 15779 41120
rect 15703 41083 15779 41089
rect 15841 41089 15853 41123
rect 15887 41089 15899 41123
rect 15841 41083 15899 41089
rect 9950 41052 9956 41064
rect 9232 41024 9956 41052
rect 9950 41012 9956 41024
rect 10008 41012 10014 41064
rect 12894 41052 12900 41064
rect 12855 41024 12900 41052
rect 12894 41012 12900 41024
rect 12952 41012 12958 41064
rect 15470 41012 15476 41064
rect 15528 41012 15534 41064
rect 15751 41052 15779 41083
rect 15930 41080 15936 41132
rect 15988 41129 15994 41132
rect 15988 41120 15996 41129
rect 15988 41092 16033 41120
rect 15988 41083 15996 41092
rect 15988 41080 15994 41083
rect 16114 41080 16120 41132
rect 16172 41120 16178 41132
rect 16172 41092 16217 41120
rect 16172 41080 16178 41092
rect 16776 41052 16804 41219
rect 17954 41216 17960 41228
rect 18012 41216 18018 41268
rect 19334 41188 19340 41200
rect 17880 41160 19340 41188
rect 17880 41129 17908 41160
rect 19334 41148 19340 41160
rect 19392 41148 19398 41200
rect 19426 41148 19432 41200
rect 19484 41188 19490 41200
rect 19806 41191 19864 41197
rect 19806 41188 19818 41191
rect 19484 41160 19818 41188
rect 19484 41148 19490 41160
rect 19806 41157 19818 41160
rect 19852 41157 19864 41191
rect 19806 41151 19864 41157
rect 17589 41123 17647 41129
rect 17589 41089 17601 41123
rect 17635 41120 17647 41123
rect 17773 41123 17831 41129
rect 17635 41092 17724 41120
rect 17635 41089 17647 41092
rect 17589 41083 17647 41089
rect 15751 41024 16804 41052
rect 10045 40987 10103 40993
rect 10045 40984 10057 40987
rect 9140 40956 10057 40984
rect 10045 40953 10057 40956
rect 10091 40984 10103 40987
rect 10962 40984 10968 40996
rect 10091 40956 10968 40984
rect 10091 40953 10103 40956
rect 10045 40947 10103 40953
rect 10962 40944 10968 40956
rect 11020 40944 11026 40996
rect 15488 40984 15516 41012
rect 16114 40984 16120 40996
rect 15488 40956 16120 40984
rect 16114 40944 16120 40956
rect 16172 40944 16178 40996
rect 17696 40984 17724 41092
rect 17773 41089 17785 41123
rect 17819 41089 17831 41123
rect 17773 41083 17831 41089
rect 17865 41123 17923 41129
rect 17865 41089 17877 41123
rect 17911 41089 17923 41123
rect 17865 41083 17923 41089
rect 17788 41052 17816 41083
rect 17954 41080 17960 41132
rect 18012 41120 18018 41132
rect 23934 41120 23940 41132
rect 18012 41092 23940 41120
rect 18012 41080 18018 41092
rect 23934 41080 23940 41092
rect 23992 41080 23998 41132
rect 27798 41080 27804 41132
rect 27856 41120 27862 41132
rect 27965 41123 28023 41129
rect 27965 41120 27977 41123
rect 27856 41092 27977 41120
rect 27856 41080 27862 41092
rect 27965 41089 27977 41092
rect 28011 41089 28023 41123
rect 27965 41083 28023 41089
rect 18414 41052 18420 41064
rect 17788 41024 18420 41052
rect 18414 41012 18420 41024
rect 18472 41012 18478 41064
rect 20073 41055 20131 41061
rect 20073 41021 20085 41055
rect 20119 41021 20131 41055
rect 27706 41052 27712 41064
rect 27667 41024 27712 41052
rect 20073 41015 20131 41021
rect 17954 40984 17960 40996
rect 17696 40956 17960 40984
rect 17954 40944 17960 40956
rect 18012 40944 18018 40996
rect 6914 40916 6920 40928
rect 6748 40888 6920 40916
rect 5169 40879 5227 40885
rect 6914 40876 6920 40888
rect 6972 40876 6978 40928
rect 8110 40916 8116 40928
rect 8071 40888 8116 40916
rect 8110 40876 8116 40888
rect 8168 40876 8174 40928
rect 10597 40919 10655 40925
rect 10597 40885 10609 40919
rect 10643 40916 10655 40919
rect 11422 40916 11428 40928
rect 10643 40888 11428 40916
rect 10643 40885 10655 40888
rect 10597 40879 10655 40885
rect 11422 40876 11428 40888
rect 11480 40876 11486 40928
rect 11514 40876 11520 40928
rect 11572 40916 11578 40928
rect 11698 40916 11704 40928
rect 11572 40888 11704 40916
rect 11572 40876 11578 40888
rect 11698 40876 11704 40888
rect 11756 40876 11762 40928
rect 13633 40919 13691 40925
rect 13633 40885 13645 40919
rect 13679 40916 13691 40919
rect 13814 40916 13820 40928
rect 13679 40888 13820 40916
rect 13679 40885 13691 40888
rect 13633 40879 13691 40885
rect 13814 40876 13820 40888
rect 13872 40876 13878 40928
rect 15470 40916 15476 40928
rect 15431 40888 15476 40916
rect 15470 40876 15476 40888
rect 15528 40876 15534 40928
rect 18233 40919 18291 40925
rect 18233 40885 18245 40919
rect 18279 40916 18291 40919
rect 18598 40916 18604 40928
rect 18279 40888 18604 40916
rect 18279 40885 18291 40888
rect 18233 40879 18291 40885
rect 18598 40876 18604 40888
rect 18656 40876 18662 40928
rect 18690 40876 18696 40928
rect 18748 40916 18754 40928
rect 18748 40888 18793 40916
rect 18748 40876 18754 40888
rect 19334 40876 19340 40928
rect 19392 40916 19398 40928
rect 20088 40916 20116 41015
rect 27706 41012 27712 41024
rect 27764 41012 27770 41064
rect 23106 40916 23112 40928
rect 19392 40888 20116 40916
rect 23067 40888 23112 40916
rect 19392 40876 19398 40888
rect 23106 40876 23112 40888
rect 23164 40876 23170 40928
rect 29089 40919 29147 40925
rect 29089 40885 29101 40919
rect 29135 40916 29147 40919
rect 29270 40916 29276 40928
rect 29135 40888 29276 40916
rect 29135 40885 29147 40888
rect 29089 40879 29147 40885
rect 29270 40876 29276 40888
rect 29328 40876 29334 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 8021 40715 8079 40721
rect 8021 40681 8033 40715
rect 8067 40712 8079 40715
rect 9306 40712 9312 40724
rect 8067 40684 9312 40712
rect 8067 40681 8079 40684
rect 8021 40675 8079 40681
rect 9306 40672 9312 40684
rect 9364 40672 9370 40724
rect 27798 40712 27804 40724
rect 27759 40684 27804 40712
rect 27798 40672 27804 40684
rect 27856 40672 27862 40724
rect 27706 40536 27712 40588
rect 27764 40576 27770 40588
rect 29914 40576 29920 40588
rect 27764 40548 29920 40576
rect 27764 40536 27770 40548
rect 29914 40536 29920 40548
rect 29972 40536 29978 40588
rect 4430 40508 4436 40520
rect 4391 40480 4436 40508
rect 4430 40468 4436 40480
rect 4488 40468 4494 40520
rect 4614 40508 4620 40520
rect 4575 40480 4620 40508
rect 4614 40468 4620 40480
rect 4672 40468 4678 40520
rect 4706 40468 4712 40520
rect 4764 40508 4770 40520
rect 4847 40511 4905 40517
rect 4764 40480 4809 40508
rect 4764 40468 4770 40480
rect 4847 40477 4859 40511
rect 4893 40508 4905 40511
rect 5166 40508 5172 40520
rect 4893 40480 5172 40508
rect 4893 40477 4905 40480
rect 4847 40471 4905 40477
rect 5166 40468 5172 40480
rect 5224 40468 5230 40520
rect 6914 40508 6920 40520
rect 6827 40480 6920 40508
rect 6914 40468 6920 40480
rect 6972 40508 6978 40520
rect 8478 40508 8484 40520
rect 6972 40480 8484 40508
rect 6972 40468 6978 40480
rect 8478 40468 8484 40480
rect 8536 40508 8542 40520
rect 8941 40511 8999 40517
rect 8941 40508 8953 40511
rect 8536 40480 8953 40508
rect 8536 40468 8542 40480
rect 8941 40477 8953 40480
rect 8987 40508 8999 40511
rect 10502 40508 10508 40520
rect 8987 40480 10508 40508
rect 8987 40477 8999 40480
rect 8941 40471 8999 40477
rect 10502 40468 10508 40480
rect 10560 40468 10566 40520
rect 12894 40508 12900 40520
rect 12807 40480 12900 40508
rect 12894 40468 12900 40480
rect 12952 40508 12958 40520
rect 14918 40508 14924 40520
rect 12952 40480 14924 40508
rect 12952 40468 12958 40480
rect 14918 40468 14924 40480
rect 14976 40508 14982 40520
rect 16761 40511 16819 40517
rect 16761 40508 16773 40511
rect 14976 40480 16773 40508
rect 14976 40468 14982 40480
rect 16761 40477 16773 40480
rect 16807 40508 16819 40511
rect 16850 40508 16856 40520
rect 16807 40480 16856 40508
rect 16807 40477 16819 40480
rect 16761 40471 16819 40477
rect 16850 40468 16856 40480
rect 16908 40508 16914 40520
rect 19245 40511 19303 40517
rect 19245 40508 19257 40511
rect 16908 40480 19257 40508
rect 16908 40468 16914 40480
rect 19245 40477 19257 40480
rect 19291 40508 19303 40511
rect 19334 40508 19340 40520
rect 19291 40480 19340 40508
rect 19291 40477 19303 40480
rect 19245 40471 19303 40477
rect 19334 40468 19340 40480
rect 19392 40468 19398 40520
rect 23845 40511 23903 40517
rect 23845 40477 23857 40511
rect 23891 40508 23903 40511
rect 25777 40511 25835 40517
rect 25777 40508 25789 40511
rect 23891 40480 25789 40508
rect 23891 40477 23903 40480
rect 23845 40471 23903 40477
rect 25777 40477 25789 40480
rect 25823 40508 25835 40511
rect 25958 40508 25964 40520
rect 25823 40480 25964 40508
rect 25823 40477 25835 40480
rect 25777 40471 25835 40477
rect 25958 40468 25964 40480
rect 26016 40468 26022 40520
rect 27246 40468 27252 40520
rect 27304 40508 27310 40520
rect 27341 40511 27399 40517
rect 27341 40508 27353 40511
rect 27304 40480 27353 40508
rect 27304 40468 27310 40480
rect 27341 40477 27353 40480
rect 27387 40508 27399 40511
rect 28077 40511 28135 40517
rect 28077 40508 28089 40511
rect 27387 40480 28089 40508
rect 27387 40477 27399 40480
rect 27341 40471 27399 40477
rect 28077 40477 28089 40480
rect 28123 40477 28135 40511
rect 28077 40471 28135 40477
rect 28169 40511 28227 40517
rect 28169 40477 28181 40511
rect 28215 40477 28227 40511
rect 28169 40471 28227 40477
rect 28261 40511 28319 40517
rect 28261 40477 28273 40511
rect 28307 40477 28319 40511
rect 28442 40508 28448 40520
rect 28403 40480 28448 40508
rect 28261 40471 28319 40477
rect 6672 40443 6730 40449
rect 6672 40409 6684 40443
rect 6718 40440 6730 40443
rect 7006 40440 7012 40452
rect 6718 40412 7012 40440
rect 6718 40409 6730 40412
rect 6672 40403 6730 40409
rect 7006 40400 7012 40412
rect 7064 40400 7070 40452
rect 8110 40400 8116 40452
rect 8168 40440 8174 40452
rect 8205 40443 8263 40449
rect 8205 40440 8217 40443
rect 8168 40412 8217 40440
rect 8168 40400 8174 40412
rect 8205 40409 8217 40412
rect 8251 40409 8263 40443
rect 8205 40403 8263 40409
rect 8389 40443 8447 40449
rect 8389 40409 8401 40443
rect 8435 40440 8447 40443
rect 9030 40440 9036 40452
rect 8435 40412 9036 40440
rect 8435 40409 8447 40412
rect 8389 40403 8447 40409
rect 5074 40372 5080 40384
rect 5035 40344 5080 40372
rect 5074 40332 5080 40344
rect 5132 40332 5138 40384
rect 5534 40372 5540 40384
rect 5495 40344 5540 40372
rect 5534 40332 5540 40344
rect 5592 40332 5598 40384
rect 8220 40372 8248 40403
rect 9030 40400 9036 40412
rect 9088 40400 9094 40452
rect 9208 40443 9266 40449
rect 9208 40409 9220 40443
rect 9254 40440 9266 40443
rect 10226 40440 10232 40452
rect 9254 40412 10232 40440
rect 9254 40409 9266 40412
rect 9208 40403 9266 40409
rect 10226 40400 10232 40412
rect 10284 40400 10290 40452
rect 12526 40400 12532 40452
rect 12584 40440 12590 40452
rect 12630 40443 12688 40449
rect 12630 40440 12642 40443
rect 12584 40412 12642 40440
rect 12584 40400 12590 40412
rect 12630 40409 12642 40412
rect 12676 40409 12688 40443
rect 12630 40403 12688 40409
rect 15188 40443 15246 40449
rect 15188 40409 15200 40443
rect 15234 40440 15246 40443
rect 15470 40440 15476 40452
rect 15234 40412 15476 40440
rect 15234 40409 15246 40412
rect 15188 40403 15246 40409
rect 15470 40400 15476 40412
rect 15528 40400 15534 40452
rect 18506 40440 18512 40452
rect 18467 40412 18512 40440
rect 18506 40400 18512 40412
rect 18564 40400 18570 40452
rect 18598 40400 18604 40452
rect 18656 40440 18662 40452
rect 19490 40443 19548 40449
rect 19490 40440 19502 40443
rect 18656 40412 19502 40440
rect 18656 40400 18662 40412
rect 19490 40409 19502 40412
rect 19536 40409 19548 40443
rect 19490 40403 19548 40409
rect 23474 40400 23480 40452
rect 23532 40440 23538 40452
rect 23578 40443 23636 40449
rect 23578 40440 23590 40443
rect 23532 40412 23590 40440
rect 23532 40400 23538 40412
rect 23578 40409 23590 40412
rect 23624 40409 23636 40443
rect 23578 40403 23636 40409
rect 23750 40400 23756 40452
rect 23808 40440 23814 40452
rect 25510 40443 25568 40449
rect 25510 40440 25522 40443
rect 23808 40412 25522 40440
rect 23808 40400 23814 40412
rect 25510 40409 25522 40412
rect 25556 40409 25568 40443
rect 25510 40403 25568 40409
rect 9858 40372 9864 40384
rect 8220 40344 9864 40372
rect 9858 40332 9864 40344
rect 9916 40332 9922 40384
rect 10321 40375 10379 40381
rect 10321 40341 10333 40375
rect 10367 40372 10379 40375
rect 10594 40372 10600 40384
rect 10367 40344 10600 40372
rect 10367 40341 10379 40344
rect 10321 40335 10379 40341
rect 10594 40332 10600 40344
rect 10652 40332 10658 40384
rect 11517 40375 11575 40381
rect 11517 40341 11529 40375
rect 11563 40372 11575 40375
rect 12434 40372 12440 40384
rect 11563 40344 12440 40372
rect 11563 40341 11575 40344
rect 11517 40335 11575 40341
rect 12434 40332 12440 40344
rect 12492 40332 12498 40384
rect 15562 40332 15568 40384
rect 15620 40372 15626 40384
rect 16298 40372 16304 40384
rect 15620 40344 16304 40372
rect 15620 40332 15626 40344
rect 16298 40332 16304 40344
rect 16356 40332 16362 40384
rect 18782 40332 18788 40384
rect 18840 40372 18846 40384
rect 20625 40375 20683 40381
rect 20625 40372 20637 40375
rect 18840 40344 20637 40372
rect 18840 40332 18846 40344
rect 20625 40341 20637 40344
rect 20671 40341 20683 40375
rect 20625 40335 20683 40341
rect 22465 40375 22523 40381
rect 22465 40341 22477 40375
rect 22511 40372 22523 40375
rect 22646 40372 22652 40384
rect 22511 40344 22652 40372
rect 22511 40341 22523 40344
rect 22465 40335 22523 40341
rect 22646 40332 22652 40344
rect 22704 40332 22710 40384
rect 24302 40332 24308 40384
rect 24360 40372 24366 40384
rect 24397 40375 24455 40381
rect 24397 40372 24409 40375
rect 24360 40344 24409 40372
rect 24360 40332 24366 40344
rect 24397 40341 24409 40344
rect 24443 40341 24455 40375
rect 28184 40372 28212 40471
rect 28276 40440 28304 40471
rect 28442 40468 28448 40480
rect 28500 40468 28506 40520
rect 58158 40508 58164 40520
rect 58119 40480 58164 40508
rect 58158 40468 58164 40480
rect 58216 40468 58222 40520
rect 29546 40440 29552 40452
rect 28276 40412 29552 40440
rect 29546 40400 29552 40412
rect 29604 40400 29610 40452
rect 30184 40443 30242 40449
rect 30184 40409 30196 40443
rect 30230 40440 30242 40443
rect 30282 40440 30288 40452
rect 30230 40412 30288 40440
rect 30230 40409 30242 40412
rect 30184 40403 30242 40409
rect 30282 40400 30288 40412
rect 30340 40400 30346 40452
rect 28902 40372 28908 40384
rect 28184 40344 28908 40372
rect 24397 40335 24455 40341
rect 28902 40332 28908 40344
rect 28960 40332 28966 40384
rect 28997 40375 29055 40381
rect 28997 40341 29009 40375
rect 29043 40372 29055 40375
rect 29086 40372 29092 40384
rect 29043 40344 29092 40372
rect 29043 40341 29055 40344
rect 28997 40335 29055 40341
rect 29086 40332 29092 40344
rect 29144 40372 29150 40384
rect 30006 40372 30012 40384
rect 29144 40344 30012 40372
rect 29144 40332 29150 40344
rect 30006 40332 30012 40344
rect 30064 40332 30070 40384
rect 31297 40375 31355 40381
rect 31297 40341 31309 40375
rect 31343 40372 31355 40375
rect 31846 40372 31852 40384
rect 31343 40344 31852 40372
rect 31343 40341 31355 40344
rect 31297 40335 31355 40341
rect 31846 40332 31852 40344
rect 31904 40332 31910 40384
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 5994 40168 6000 40180
rect 5460 40140 6000 40168
rect 5460 40109 5488 40140
rect 5994 40128 6000 40140
rect 6052 40128 6058 40180
rect 9766 40168 9772 40180
rect 9727 40140 9772 40168
rect 9766 40128 9772 40140
rect 9824 40128 9830 40180
rect 27706 40168 27712 40180
rect 27632 40140 27712 40168
rect 5445 40103 5503 40109
rect 5445 40069 5457 40103
rect 5491 40069 5503 40103
rect 5445 40063 5503 40069
rect 5534 40060 5540 40112
rect 5592 40100 5598 40112
rect 5629 40103 5687 40109
rect 5629 40100 5641 40103
rect 5592 40072 5641 40100
rect 5592 40060 5598 40072
rect 5629 40069 5641 40072
rect 5675 40100 5687 40103
rect 8570 40100 8576 40112
rect 5675 40072 8576 40100
rect 5675 40069 5687 40072
rect 5629 40063 5687 40069
rect 8570 40060 8576 40072
rect 8628 40060 8634 40112
rect 9030 40060 9036 40112
rect 9088 40100 9094 40112
rect 10318 40100 10324 40112
rect 9088 40072 10324 40100
rect 9088 40060 9094 40072
rect 10318 40060 10324 40072
rect 10376 40060 10382 40112
rect 10520 40072 11100 40100
rect 2406 40041 2412 40044
rect 2400 39995 2412 40041
rect 2464 40032 2470 40044
rect 6365 40035 6423 40041
rect 6365 40032 6377 40035
rect 2464 40004 2500 40032
rect 5552 40004 6377 40032
rect 2406 39992 2412 39995
rect 2464 39992 2470 40004
rect 2133 39967 2191 39973
rect 2133 39933 2145 39967
rect 2179 39933 2191 39967
rect 2133 39927 2191 39933
rect 3973 39967 4031 39973
rect 3973 39933 3985 39967
rect 4019 39964 4031 39967
rect 4062 39964 4068 39976
rect 4019 39936 4068 39964
rect 4019 39933 4031 39936
rect 3973 39927 4031 39933
rect 2148 39828 2176 39927
rect 4062 39924 4068 39936
rect 4120 39924 4126 39976
rect 4249 39967 4307 39973
rect 4249 39933 4261 39967
rect 4295 39964 4307 39967
rect 4430 39964 4436 39976
rect 4295 39936 4436 39964
rect 4295 39933 4307 39936
rect 4249 39927 4307 39933
rect 3234 39856 3240 39908
rect 3292 39896 3298 39908
rect 4264 39896 4292 39927
rect 4430 39924 4436 39936
rect 4488 39964 4494 39976
rect 5552 39964 5580 40004
rect 6365 40001 6377 40004
rect 6411 40001 6423 40035
rect 6365 39995 6423 40001
rect 6549 40035 6607 40041
rect 6549 40001 6561 40035
rect 6595 40001 6607 40035
rect 6549 39995 6607 40001
rect 6641 40035 6699 40041
rect 6641 40001 6653 40035
rect 6687 40001 6699 40035
rect 6641 39995 6699 40001
rect 6779 40035 6837 40041
rect 6779 40001 6791 40035
rect 6825 40032 6837 40035
rect 7098 40032 7104 40044
rect 6825 40004 7104 40032
rect 6825 40001 6837 40004
rect 6779 39995 6837 40001
rect 4488 39936 5580 39964
rect 5813 39967 5871 39973
rect 4488 39924 4494 39936
rect 5813 39933 5825 39967
rect 5859 39964 5871 39967
rect 6564 39964 6592 39995
rect 5859 39936 6592 39964
rect 5859 39933 5871 39936
rect 5813 39927 5871 39933
rect 6656 39908 6684 39995
rect 7098 39992 7104 40004
rect 7156 40032 7162 40044
rect 7469 40035 7527 40041
rect 7469 40032 7481 40035
rect 7156 40004 7481 40032
rect 7156 39992 7162 40004
rect 7469 40001 7481 40004
rect 7515 40001 7527 40035
rect 7469 39995 7527 40001
rect 8389 40035 8447 40041
rect 8389 40001 8401 40035
rect 8435 40032 8447 40035
rect 8478 40032 8484 40044
rect 8435 40004 8484 40032
rect 8435 40001 8447 40004
rect 8389 39995 8447 40001
rect 8478 39992 8484 40004
rect 8536 39992 8542 40044
rect 8656 40035 8714 40041
rect 8656 40001 8668 40035
rect 8702 40032 8714 40035
rect 9214 40032 9220 40044
rect 8702 40004 9220 40032
rect 8702 40001 8714 40004
rect 8656 39995 8714 40001
rect 9214 39992 9220 40004
rect 9272 39992 9278 40044
rect 10520 40041 10548 40072
rect 10505 40035 10563 40041
rect 10505 40001 10517 40035
rect 10551 40001 10563 40035
rect 10505 39995 10563 40001
rect 10597 40035 10655 40041
rect 10597 40001 10609 40035
rect 10643 40001 10655 40035
rect 10597 39995 10655 40001
rect 7006 39964 7012 39976
rect 6967 39936 7012 39964
rect 7006 39924 7012 39936
rect 7064 39924 7070 39976
rect 10226 39964 10232 39976
rect 10187 39936 10232 39964
rect 10226 39924 10232 39936
rect 10284 39924 10290 39976
rect 3292 39868 4292 39896
rect 3292 39856 3298 39868
rect 4706 39856 4712 39908
rect 4764 39896 4770 39908
rect 6638 39896 6644 39908
rect 4764 39868 6644 39896
rect 4764 39856 4770 39868
rect 6638 39856 6644 39868
rect 6696 39856 6702 39908
rect 9950 39856 9956 39908
rect 10008 39896 10014 39908
rect 10612 39896 10640 39995
rect 10686 39992 10692 40044
rect 10744 40032 10750 40044
rect 10873 40035 10931 40041
rect 10744 40004 10789 40032
rect 10744 39992 10750 40004
rect 10873 40001 10885 40035
rect 10919 40001 10931 40035
rect 11072 40032 11100 40072
rect 11422 40060 11428 40112
rect 11480 40100 11486 40112
rect 18782 40100 18788 40112
rect 11480 40072 12848 40100
rect 18743 40072 18788 40100
rect 11480 40060 11486 40072
rect 11606 40032 11612 40044
rect 11072 40004 11612 40032
rect 10873 39995 10931 40001
rect 10888 39964 10916 39995
rect 11606 39992 11612 40004
rect 11664 39992 11670 40044
rect 12820 40041 12848 40072
rect 18782 40060 18788 40072
rect 18840 40060 18846 40112
rect 23106 40100 23112 40112
rect 22756 40072 23112 40100
rect 12621 40035 12679 40041
rect 12621 40001 12633 40035
rect 12667 40001 12679 40035
rect 12621 39995 12679 40001
rect 12713 40035 12771 40041
rect 12713 40001 12725 40035
rect 12759 40001 12771 40035
rect 12713 39995 12771 40001
rect 12805 40035 12863 40041
rect 12805 40001 12817 40035
rect 12851 40001 12863 40035
rect 12986 40032 12992 40044
rect 12947 40004 12992 40032
rect 12805 39995 12863 40001
rect 10008 39868 10640 39896
rect 10796 39936 10916 39964
rect 12345 39967 12403 39973
rect 10008 39856 10014 39868
rect 2774 39828 2780 39840
rect 2148 39800 2780 39828
rect 2774 39788 2780 39800
rect 2832 39788 2838 39840
rect 3513 39831 3571 39837
rect 3513 39797 3525 39831
rect 3559 39828 3571 39831
rect 3970 39828 3976 39840
rect 3559 39800 3976 39828
rect 3559 39797 3571 39800
rect 3513 39791 3571 39797
rect 3970 39788 3976 39800
rect 4028 39788 4034 39840
rect 10226 39788 10232 39840
rect 10284 39828 10290 39840
rect 10796 39828 10824 39936
rect 12345 39933 12357 39967
rect 12391 39964 12403 39967
rect 12526 39964 12532 39976
rect 12391 39936 12532 39964
rect 12391 39933 12403 39936
rect 12345 39927 12403 39933
rect 12526 39924 12532 39936
rect 12584 39924 12590 39976
rect 12636 39896 12664 39995
rect 12728 39964 12756 39995
rect 12986 39992 12992 40004
rect 13044 39992 13050 40044
rect 18414 39992 18420 40044
rect 18472 40032 18478 40044
rect 18601 40035 18659 40041
rect 18601 40032 18613 40035
rect 18472 40004 18613 40032
rect 18472 39992 18478 40004
rect 18601 40001 18613 40004
rect 18647 40001 18659 40035
rect 18966 40032 18972 40044
rect 18879 40004 18972 40032
rect 18601 39995 18659 40001
rect 18966 39992 18972 40004
rect 19024 40032 19030 40044
rect 19150 40032 19156 40044
rect 19024 40004 19156 40032
rect 19024 39992 19030 40004
rect 19150 39992 19156 40004
rect 19208 39992 19214 40044
rect 19334 39992 19340 40044
rect 19392 40032 19398 40044
rect 20162 40041 20168 40044
rect 19889 40035 19947 40041
rect 19889 40032 19901 40035
rect 19392 40004 19901 40032
rect 19392 39992 19398 40004
rect 19889 40001 19901 40004
rect 19935 40001 19947 40035
rect 19889 39995 19947 40001
rect 20156 39995 20168 40041
rect 20220 40032 20226 40044
rect 20220 40004 20256 40032
rect 20162 39992 20168 39995
rect 20220 39992 20226 40004
rect 22278 39992 22284 40044
rect 22336 40032 22342 40044
rect 22373 40035 22431 40041
rect 22373 40032 22385 40035
rect 22336 40004 22385 40032
rect 22336 39992 22342 40004
rect 22373 40001 22385 40004
rect 22419 40001 22431 40035
rect 22554 40032 22560 40044
rect 22515 40004 22560 40032
rect 22373 39995 22431 40001
rect 22554 39992 22560 40004
rect 22612 39992 22618 40044
rect 22756 40041 22784 40072
rect 23106 40060 23112 40072
rect 23164 40100 23170 40112
rect 24946 40100 24952 40112
rect 23164 40072 24952 40100
rect 23164 40060 23170 40072
rect 24946 40060 24952 40072
rect 25004 40060 25010 40112
rect 22649 40035 22707 40041
rect 22649 40001 22661 40035
rect 22695 40001 22707 40035
rect 22649 39995 22707 40001
rect 22741 40035 22799 40041
rect 22741 40001 22753 40035
rect 22787 40001 22799 40035
rect 22741 39995 22799 40001
rect 12894 39964 12900 39976
rect 12728 39936 12900 39964
rect 12894 39924 12900 39936
rect 12952 39964 12958 39976
rect 13354 39964 13360 39976
rect 12952 39936 13360 39964
rect 12952 39924 12958 39936
rect 13354 39924 13360 39936
rect 13412 39924 13418 39976
rect 22664 39964 22692 39995
rect 23198 39992 23204 40044
rect 23256 40032 23262 40044
rect 24590 40035 24648 40041
rect 24590 40032 24602 40035
rect 23256 40004 24602 40032
rect 23256 39992 23262 40004
rect 24590 40001 24602 40004
rect 24636 40001 24648 40035
rect 27632 40032 27660 40140
rect 27706 40128 27712 40140
rect 27764 40128 27770 40180
rect 28813 40171 28871 40177
rect 28813 40137 28825 40171
rect 28859 40168 28871 40171
rect 28994 40168 29000 40180
rect 28859 40140 29000 40168
rect 28859 40137 28871 40140
rect 28813 40131 28871 40137
rect 28994 40128 29000 40140
rect 29052 40128 29058 40180
rect 30282 40168 30288 40180
rect 30243 40140 30288 40168
rect 30282 40128 30288 40140
rect 30340 40128 30346 40180
rect 30745 40103 30803 40109
rect 30745 40100 30757 40103
rect 29840 40072 30757 40100
rect 27706 40041 27712 40044
rect 24590 39995 24648 40001
rect 27448 40004 27660 40032
rect 22830 39964 22836 39976
rect 13464 39936 19932 39964
rect 22664 39936 22836 39964
rect 13464 39905 13492 39936
rect 13449 39899 13507 39905
rect 13449 39896 13461 39899
rect 12636 39868 13461 39896
rect 13449 39865 13461 39868
rect 13495 39865 13507 39899
rect 19426 39896 19432 39908
rect 13449 39859 13507 39865
rect 18524 39868 19432 39896
rect 18524 39840 18552 39868
rect 19426 39856 19432 39868
rect 19484 39856 19490 39908
rect 11606 39828 11612 39840
rect 10284 39800 10824 39828
rect 11567 39800 11612 39828
rect 10284 39788 10290 39800
rect 11606 39788 11612 39800
rect 11664 39788 11670 39840
rect 16666 39828 16672 39840
rect 16627 39800 16672 39828
rect 16666 39788 16672 39800
rect 16724 39828 16730 39840
rect 18506 39828 18512 39840
rect 16724 39800 18512 39828
rect 16724 39788 16730 39800
rect 18506 39788 18512 39800
rect 18564 39788 18570 39840
rect 19904 39828 19932 39936
rect 22830 39924 22836 39936
rect 22888 39924 22894 39976
rect 23017 39967 23075 39973
rect 23017 39933 23029 39967
rect 23063 39964 23075 39967
rect 23750 39964 23756 39976
rect 23063 39936 23756 39964
rect 23063 39933 23075 39936
rect 23017 39927 23075 39933
rect 23750 39924 23756 39936
rect 23808 39924 23814 39976
rect 24857 39967 24915 39973
rect 24857 39933 24869 39967
rect 24903 39964 24915 39967
rect 25958 39964 25964 39976
rect 24903 39936 25964 39964
rect 24903 39933 24915 39936
rect 24857 39927 24915 39933
rect 25958 39924 25964 39936
rect 26016 39964 26022 39976
rect 27448 39973 27476 40004
rect 27700 39995 27712 40041
rect 27764 40032 27770 40044
rect 27764 40004 27800 40032
rect 27706 39992 27712 39995
rect 27764 39992 27770 40004
rect 28442 39992 28448 40044
rect 28500 40032 28506 40044
rect 29840 40041 29868 40072
rect 30745 40069 30757 40072
rect 30791 40069 30803 40103
rect 30745 40063 30803 40069
rect 30929 40103 30987 40109
rect 30929 40069 30941 40103
rect 30975 40100 30987 40103
rect 31846 40100 31852 40112
rect 30975 40072 31852 40100
rect 30975 40069 30987 40072
rect 30929 40063 30987 40069
rect 31846 40060 31852 40072
rect 31904 40060 31910 40112
rect 29641 40035 29699 40041
rect 29641 40032 29653 40035
rect 28500 40004 29653 40032
rect 28500 39992 28506 40004
rect 29641 40001 29653 40004
rect 29687 40001 29699 40035
rect 29641 39995 29699 40001
rect 29825 40035 29883 40041
rect 29825 40001 29837 40035
rect 29871 40001 29883 40035
rect 29825 39995 29883 40001
rect 29917 40035 29975 40041
rect 29917 40001 29929 40035
rect 29963 40001 29975 40035
rect 29917 39995 29975 40001
rect 27433 39967 27491 39973
rect 27433 39964 27445 39967
rect 26016 39936 27445 39964
rect 26016 39924 26022 39936
rect 27433 39933 27445 39936
rect 27479 39933 27491 39967
rect 27433 39927 27491 39933
rect 29178 39856 29184 39908
rect 29236 39896 29242 39908
rect 29932 39896 29960 39995
rect 30006 39992 30012 40044
rect 30064 40032 30070 40044
rect 31113 40035 31171 40041
rect 30064 40004 30109 40032
rect 30064 39992 30070 40004
rect 31113 40001 31125 40035
rect 31159 40032 31171 40035
rect 31202 40032 31208 40044
rect 31159 40004 31208 40032
rect 31159 40001 31171 40004
rect 31113 39995 31171 40001
rect 31202 39992 31208 40004
rect 31260 39992 31266 40044
rect 30098 39896 30104 39908
rect 29236 39868 30104 39896
rect 29236 39856 29242 39868
rect 30098 39856 30104 39868
rect 30156 39856 30162 39908
rect 20254 39828 20260 39840
rect 19904 39800 20260 39828
rect 20254 39788 20260 39800
rect 20312 39788 20318 39840
rect 21266 39828 21272 39840
rect 21227 39800 21272 39828
rect 21266 39788 21272 39800
rect 21324 39788 21330 39840
rect 23477 39831 23535 39837
rect 23477 39797 23489 39831
rect 23523 39828 23535 39831
rect 23658 39828 23664 39840
rect 23523 39800 23664 39828
rect 23523 39797 23535 39800
rect 23477 39791 23535 39797
rect 23658 39788 23664 39800
rect 23716 39788 23722 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 2406 39584 2412 39636
rect 2464 39624 2470 39636
rect 2593 39627 2651 39633
rect 2593 39624 2605 39627
rect 2464 39596 2605 39624
rect 2464 39584 2470 39596
rect 2593 39593 2605 39596
rect 2639 39593 2651 39627
rect 6362 39624 6368 39636
rect 6323 39596 6368 39624
rect 2593 39587 2651 39593
rect 6362 39584 6368 39596
rect 6420 39584 6426 39636
rect 9214 39624 9220 39636
rect 9175 39596 9220 39624
rect 9214 39584 9220 39596
rect 9272 39584 9278 39636
rect 10686 39624 10692 39636
rect 10647 39596 10692 39624
rect 10686 39584 10692 39596
rect 10744 39584 10750 39636
rect 20073 39627 20131 39633
rect 20073 39593 20085 39627
rect 20119 39624 20131 39627
rect 20162 39624 20168 39636
rect 20119 39596 20168 39624
rect 20119 39593 20131 39596
rect 20073 39587 20131 39593
rect 20162 39584 20168 39596
rect 20220 39584 20226 39636
rect 20346 39584 20352 39636
rect 20404 39624 20410 39636
rect 20533 39627 20591 39633
rect 20533 39624 20545 39627
rect 20404 39596 20545 39624
rect 20404 39584 20410 39596
rect 20533 39593 20545 39596
rect 20579 39593 20591 39627
rect 20533 39587 20591 39593
rect 22097 39627 22155 39633
rect 22097 39593 22109 39627
rect 22143 39624 22155 39627
rect 22554 39624 22560 39636
rect 22143 39596 22560 39624
rect 22143 39593 22155 39596
rect 22097 39587 22155 39593
rect 22554 39584 22560 39596
rect 22612 39584 22618 39636
rect 23198 39624 23204 39636
rect 23159 39596 23204 39624
rect 23198 39584 23204 39596
rect 23256 39584 23262 39636
rect 29546 39624 29552 39636
rect 29507 39596 29552 39624
rect 29546 39584 29552 39596
rect 29604 39584 29610 39636
rect 19978 39556 19984 39568
rect 19444 39528 19984 39556
rect 4706 39488 4712 39500
rect 2976 39460 4712 39488
rect 2866 39420 2872 39432
rect 2827 39392 2872 39420
rect 2866 39380 2872 39392
rect 2924 39380 2930 39432
rect 2976 39429 3004 39460
rect 4706 39448 4712 39460
rect 4764 39448 4770 39500
rect 11149 39491 11207 39497
rect 11149 39488 11161 39491
rect 9508 39460 11161 39488
rect 2961 39423 3019 39429
rect 2961 39389 2973 39423
rect 3007 39389 3019 39423
rect 2961 39383 3019 39389
rect 3053 39423 3111 39429
rect 3053 39389 3065 39423
rect 3099 39389 3111 39423
rect 3234 39420 3240 39432
rect 3195 39392 3240 39420
rect 3053 39383 3111 39389
rect 2590 39312 2596 39364
rect 2648 39352 2654 39364
rect 2976 39352 3004 39383
rect 2648 39324 3004 39352
rect 3068 39352 3096 39383
rect 3234 39380 3240 39392
rect 3292 39380 3298 39432
rect 3786 39380 3792 39432
rect 3844 39420 3850 39432
rect 4985 39423 5043 39429
rect 4985 39420 4997 39423
rect 3844 39392 4997 39420
rect 3844 39380 3850 39392
rect 4985 39389 4997 39392
rect 5031 39389 5043 39423
rect 4985 39383 5043 39389
rect 5074 39380 5080 39432
rect 5132 39420 5138 39432
rect 9508 39429 9536 39460
rect 11149 39457 11161 39460
rect 11195 39488 11207 39491
rect 11195 39460 12434 39488
rect 11195 39457 11207 39460
rect 11149 39451 11207 39457
rect 5241 39423 5299 39429
rect 5241 39420 5253 39423
rect 5132 39392 5253 39420
rect 5132 39380 5138 39392
rect 5241 39389 5253 39392
rect 5287 39389 5299 39423
rect 5241 39383 5299 39389
rect 9493 39423 9551 39429
rect 9493 39389 9505 39423
rect 9539 39389 9551 39423
rect 9493 39383 9551 39389
rect 9585 39423 9643 39429
rect 9585 39389 9597 39423
rect 9631 39389 9643 39423
rect 9585 39383 9643 39389
rect 3970 39352 3976 39364
rect 3068 39324 3832 39352
rect 3931 39324 3976 39352
rect 2648 39312 2654 39324
rect 3804 39293 3832 39324
rect 3970 39312 3976 39324
rect 4028 39312 4034 39364
rect 4157 39355 4215 39361
rect 4157 39321 4169 39355
rect 4203 39352 4215 39355
rect 5994 39352 6000 39364
rect 4203 39324 6000 39352
rect 4203 39321 4215 39324
rect 4157 39315 4215 39321
rect 5994 39312 6000 39324
rect 6052 39312 6058 39364
rect 9600 39352 9628 39383
rect 9674 39380 9680 39432
rect 9732 39420 9738 39432
rect 9861 39423 9919 39429
rect 9732 39392 9777 39420
rect 9732 39380 9738 39392
rect 9861 39389 9873 39423
rect 9907 39420 9919 39423
rect 10318 39420 10324 39432
rect 9907 39392 10088 39420
rect 10279 39392 10324 39420
rect 9907 39389 9919 39392
rect 9861 39383 9919 39389
rect 9950 39352 9956 39364
rect 9600 39324 9956 39352
rect 9950 39312 9956 39324
rect 10008 39312 10014 39364
rect 10060 39352 10088 39392
rect 10318 39380 10324 39392
rect 10376 39380 10382 39432
rect 10226 39352 10232 39364
rect 10060 39324 10232 39352
rect 10226 39312 10232 39324
rect 10284 39312 10290 39364
rect 10505 39355 10563 39361
rect 10505 39321 10517 39355
rect 10551 39352 10563 39355
rect 10594 39352 10600 39364
rect 10551 39324 10600 39352
rect 10551 39321 10563 39324
rect 10505 39315 10563 39321
rect 10594 39312 10600 39324
rect 10652 39312 10658 39364
rect 3789 39287 3847 39293
rect 3789 39253 3801 39287
rect 3835 39253 3847 39287
rect 12406 39284 12434 39460
rect 19444 39429 19472 39528
rect 19978 39516 19984 39528
rect 20036 39516 20042 39568
rect 19518 39448 19524 39500
rect 19576 39488 19582 39500
rect 24302 39488 24308 39500
rect 19576 39460 19748 39488
rect 19576 39448 19582 39460
rect 19720 39429 19748 39460
rect 22664 39460 24308 39488
rect 19429 39423 19487 39429
rect 19429 39420 19441 39423
rect 19260 39392 19441 39420
rect 19260 39296 19288 39392
rect 19429 39389 19441 39392
rect 19475 39389 19487 39423
rect 19429 39383 19487 39389
rect 19613 39423 19671 39429
rect 19613 39389 19625 39423
rect 19659 39389 19671 39423
rect 19613 39383 19671 39389
rect 19705 39423 19763 39429
rect 19705 39389 19717 39423
rect 19751 39389 19763 39423
rect 19705 39383 19763 39389
rect 19797 39423 19855 39429
rect 19797 39389 19809 39423
rect 19843 39420 19855 39423
rect 20346 39420 20352 39432
rect 19843 39392 20352 39420
rect 19843 39389 19855 39392
rect 19797 39383 19855 39389
rect 19334 39312 19340 39364
rect 19392 39352 19398 39364
rect 19628 39352 19656 39383
rect 19392 39324 19656 39352
rect 19720 39352 19748 39383
rect 20346 39380 20352 39392
rect 20404 39380 20410 39432
rect 21729 39423 21787 39429
rect 21729 39389 21741 39423
rect 21775 39420 21787 39423
rect 22094 39420 22100 39432
rect 21775 39392 22100 39420
rect 21775 39389 21787 39392
rect 21729 39383 21787 39389
rect 22094 39380 22100 39392
rect 22152 39380 22158 39432
rect 22278 39380 22284 39432
rect 22336 39420 22342 39432
rect 22557 39423 22615 39429
rect 22557 39420 22569 39423
rect 22336 39392 22569 39420
rect 22336 39380 22342 39392
rect 22557 39389 22569 39392
rect 22603 39389 22615 39423
rect 22557 39383 22615 39389
rect 19978 39352 19984 39364
rect 19720 39324 19984 39352
rect 19392 39312 19398 39324
rect 19978 39312 19984 39324
rect 20036 39312 20042 39364
rect 21913 39355 21971 39361
rect 21913 39321 21925 39355
rect 21959 39352 21971 39355
rect 22664 39352 22692 39460
rect 24302 39448 24308 39460
rect 24360 39448 24366 39500
rect 22741 39423 22799 39429
rect 22741 39389 22753 39423
rect 22787 39389 22799 39423
rect 22741 39383 22799 39389
rect 21959 39324 22692 39352
rect 22756 39352 22784 39383
rect 22830 39380 22836 39432
rect 22888 39420 22894 39432
rect 22971 39423 23029 39429
rect 22888 39392 22933 39420
rect 22888 39380 22894 39392
rect 22971 39389 22983 39423
rect 23017 39420 23029 39423
rect 23106 39420 23112 39432
rect 23017 39392 23112 39420
rect 23017 39389 23029 39392
rect 22971 39383 23029 39389
rect 23106 39380 23112 39392
rect 23164 39420 23170 39432
rect 23661 39423 23719 39429
rect 23661 39420 23673 39423
rect 23164 39392 23673 39420
rect 23164 39380 23170 39392
rect 23661 39389 23673 39392
rect 23707 39389 23719 39423
rect 23661 39383 23719 39389
rect 26789 39423 26847 39429
rect 26789 39389 26801 39423
rect 26835 39420 26847 39423
rect 30377 39423 30435 39429
rect 30377 39420 30389 39423
rect 26835 39392 30389 39420
rect 26835 39389 26847 39392
rect 26789 39383 26847 39389
rect 30377 39389 30389 39392
rect 30423 39420 30435 39423
rect 31754 39420 31760 39432
rect 30423 39392 31760 39420
rect 30423 39389 30435 39392
rect 30377 39383 30435 39389
rect 31754 39380 31760 39392
rect 31812 39380 31818 39432
rect 31849 39423 31907 39429
rect 31849 39389 31861 39423
rect 31895 39420 31907 39423
rect 33318 39420 33324 39432
rect 31895 39392 33324 39420
rect 31895 39389 31907 39392
rect 31849 39383 31907 39389
rect 33318 39380 33324 39392
rect 33376 39380 33382 39432
rect 23842 39352 23848 39364
rect 22756 39324 23848 39352
rect 21959 39321 21971 39324
rect 21913 39315 21971 39321
rect 23842 39312 23848 39324
rect 23900 39312 23906 39364
rect 29270 39312 29276 39364
rect 29328 39352 29334 39364
rect 32122 39361 32128 39364
rect 29733 39355 29791 39361
rect 29733 39352 29745 39355
rect 29328 39324 29745 39352
rect 29328 39312 29334 39324
rect 29733 39321 29745 39324
rect 29779 39321 29791 39355
rect 29733 39315 29791 39321
rect 29917 39355 29975 39361
rect 29917 39321 29929 39355
rect 29963 39321 29975 39355
rect 29917 39315 29975 39321
rect 32116 39315 32128 39361
rect 32180 39352 32186 39364
rect 32180 39324 32216 39352
rect 14366 39284 14372 39296
rect 12406 39256 14372 39284
rect 3789 39247 3847 39253
rect 14366 39244 14372 39256
rect 14424 39244 14430 39296
rect 17954 39244 17960 39296
rect 18012 39284 18018 39296
rect 18693 39287 18751 39293
rect 18693 39284 18705 39287
rect 18012 39256 18705 39284
rect 18012 39244 18018 39256
rect 18693 39253 18705 39256
rect 18739 39284 18751 39287
rect 19242 39284 19248 39296
rect 18739 39256 19248 39284
rect 18739 39253 18751 39256
rect 18693 39247 18751 39253
rect 19242 39244 19248 39256
rect 19300 39244 19306 39296
rect 25958 39244 25964 39296
rect 26016 39284 26022 39296
rect 28077 39287 28135 39293
rect 28077 39284 28089 39287
rect 26016 39256 28089 39284
rect 26016 39244 26022 39256
rect 28077 39253 28089 39256
rect 28123 39253 28135 39287
rect 29932 39284 29960 39315
rect 32122 39312 32128 39315
rect 32180 39312 32186 39324
rect 30374 39284 30380 39296
rect 29932 39256 30380 39284
rect 28077 39247 28135 39253
rect 30374 39244 30380 39256
rect 30432 39244 30438 39296
rect 31389 39287 31447 39293
rect 31389 39253 31401 39287
rect 31435 39284 31447 39287
rect 31662 39284 31668 39296
rect 31435 39256 31668 39284
rect 31435 39253 31447 39256
rect 31389 39247 31447 39253
rect 31662 39244 31668 39256
rect 31720 39244 31726 39296
rect 33226 39284 33232 39296
rect 33187 39256 33232 39284
rect 33226 39244 33232 39256
rect 33284 39244 33290 39296
rect 33781 39287 33839 39293
rect 33781 39253 33793 39287
rect 33827 39284 33839 39287
rect 34514 39284 34520 39296
rect 33827 39256 34520 39284
rect 33827 39253 33839 39256
rect 33781 39247 33839 39253
rect 34514 39244 34520 39256
rect 34572 39244 34578 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 4062 39040 4068 39092
rect 4120 39080 4126 39092
rect 4893 39083 4951 39089
rect 4893 39080 4905 39083
rect 4120 39052 4905 39080
rect 4120 39040 4126 39052
rect 4893 39049 4905 39052
rect 4939 39080 4951 39083
rect 12066 39080 12072 39092
rect 4939 39052 12072 39080
rect 4939 39049 4951 39052
rect 4893 39043 4951 39049
rect 12066 39040 12072 39052
rect 12124 39040 12130 39092
rect 19334 39040 19340 39092
rect 19392 39080 19398 39092
rect 19521 39083 19579 39089
rect 19521 39080 19533 39083
rect 19392 39052 19533 39080
rect 19392 39040 19398 39052
rect 19521 39049 19533 39052
rect 19567 39049 19579 39083
rect 19521 39043 19579 39049
rect 23017 39083 23075 39089
rect 23017 39049 23029 39083
rect 23063 39080 23075 39083
rect 23474 39080 23480 39092
rect 23063 39052 23480 39080
rect 23063 39049 23075 39052
rect 23017 39043 23075 39049
rect 23474 39040 23480 39052
rect 23532 39040 23538 39092
rect 23842 39080 23848 39092
rect 23803 39052 23848 39080
rect 23842 39040 23848 39052
rect 23900 39040 23906 39092
rect 27706 39080 27712 39092
rect 27667 39052 27712 39080
rect 27706 39040 27712 39052
rect 27764 39040 27770 39092
rect 32122 39080 32128 39092
rect 32083 39052 32128 39080
rect 32122 39040 32128 39052
rect 32180 39040 32186 39092
rect 21910 38972 21916 39024
rect 21968 39012 21974 39024
rect 29181 39015 29239 39021
rect 21968 38984 22784 39012
rect 21968 38972 21974 38984
rect 5718 38904 5724 38956
rect 5776 38944 5782 38956
rect 8941 38947 8999 38953
rect 8941 38944 8953 38947
rect 5776 38916 8953 38944
rect 5776 38904 5782 38916
rect 8941 38913 8953 38916
rect 8987 38944 8999 38947
rect 11517 38947 11575 38953
rect 11517 38944 11529 38947
rect 8987 38916 11529 38944
rect 8987 38913 8999 38916
rect 8941 38907 8999 38913
rect 11517 38913 11529 38916
rect 11563 38944 11575 38947
rect 16666 38944 16672 38956
rect 11563 38916 16672 38944
rect 11563 38913 11575 38916
rect 11517 38907 11575 38913
rect 16666 38904 16672 38916
rect 16724 38904 16730 38956
rect 19150 38944 19156 38956
rect 19111 38916 19156 38944
rect 19150 38904 19156 38916
rect 19208 38904 19214 38956
rect 19334 38944 19340 38956
rect 19295 38916 19340 38944
rect 19334 38904 19340 38916
rect 19392 38944 19398 38956
rect 21266 38944 21272 38956
rect 19392 38916 21272 38944
rect 19392 38904 19398 38916
rect 21266 38904 21272 38916
rect 21324 38904 21330 38956
rect 22278 38904 22284 38956
rect 22336 38944 22342 38956
rect 22373 38947 22431 38953
rect 22373 38944 22385 38947
rect 22336 38916 22385 38944
rect 22336 38904 22342 38916
rect 22373 38913 22385 38916
rect 22419 38913 22431 38947
rect 22554 38944 22560 38956
rect 22515 38916 22560 38944
rect 22373 38907 22431 38913
rect 22554 38904 22560 38916
rect 22612 38904 22618 38956
rect 22756 38953 22784 38984
rect 29181 38981 29193 39015
rect 29227 39012 29239 39015
rect 30374 39012 30380 39024
rect 29227 38984 30380 39012
rect 29227 38981 29239 38984
rect 29181 38975 29239 38981
rect 30374 38972 30380 38984
rect 30432 39012 30438 39024
rect 31202 39012 31208 39024
rect 30432 38984 31208 39012
rect 30432 38972 30438 38984
rect 31202 38972 31208 38984
rect 31260 38972 31266 39024
rect 33134 39012 33140 39024
rect 32508 38984 33140 39012
rect 22649 38947 22707 38953
rect 22649 38913 22661 38947
rect 22695 38913 22707 38947
rect 22649 38907 22707 38913
rect 22741 38947 22799 38953
rect 22741 38913 22753 38947
rect 22787 38913 22799 38947
rect 22741 38907 22799 38913
rect 13081 38879 13139 38885
rect 13081 38845 13093 38879
rect 13127 38845 13139 38879
rect 13354 38876 13360 38888
rect 13315 38848 13360 38876
rect 13081 38839 13139 38845
rect 13096 38808 13124 38839
rect 13354 38836 13360 38848
rect 13412 38836 13418 38888
rect 20346 38836 20352 38888
rect 20404 38876 20410 38888
rect 20404 38848 22094 38876
rect 20404 38836 20410 38848
rect 13262 38808 13268 38820
rect 13096 38780 13268 38808
rect 13262 38768 13268 38780
rect 13320 38768 13326 38820
rect 22066 38808 22094 38848
rect 22186 38836 22192 38888
rect 22244 38876 22250 38888
rect 22664 38876 22692 38907
rect 22922 38904 22928 38956
rect 22980 38944 22986 38956
rect 23477 38947 23535 38953
rect 23477 38944 23489 38947
rect 22980 38916 23489 38944
rect 22980 38904 22986 38916
rect 23477 38913 23489 38916
rect 23523 38913 23535 38947
rect 23658 38944 23664 38956
rect 23619 38916 23664 38944
rect 23477 38907 23535 38913
rect 23658 38904 23664 38916
rect 23716 38904 23722 38956
rect 27985 38947 28043 38953
rect 27985 38944 27997 38947
rect 27172 38916 27997 38944
rect 22830 38876 22836 38888
rect 22244 38848 22836 38876
rect 22244 38836 22250 38848
rect 22830 38836 22836 38848
rect 22888 38836 22894 38888
rect 23566 38808 23572 38820
rect 22066 38780 23572 38808
rect 23566 38768 23572 38780
rect 23624 38768 23630 38820
rect 2866 38700 2872 38752
rect 2924 38740 2930 38752
rect 3421 38743 3479 38749
rect 3421 38740 3433 38743
rect 2924 38712 3433 38740
rect 2924 38700 2930 38712
rect 3421 38709 3433 38712
rect 3467 38740 3479 38743
rect 4706 38740 4712 38752
rect 3467 38712 4712 38740
rect 3467 38709 3479 38712
rect 3421 38703 3479 38709
rect 4706 38700 4712 38712
rect 4764 38700 4770 38752
rect 10413 38743 10471 38749
rect 10413 38709 10425 38743
rect 10459 38740 10471 38743
rect 10502 38740 10508 38752
rect 10459 38712 10508 38740
rect 10459 38709 10471 38712
rect 10413 38703 10471 38709
rect 10502 38700 10508 38712
rect 10560 38700 10566 38752
rect 11606 38700 11612 38752
rect 11664 38740 11670 38752
rect 16390 38740 16396 38752
rect 11664 38712 16396 38740
rect 11664 38700 11670 38712
rect 16390 38700 16396 38712
rect 16448 38700 16454 38752
rect 21910 38740 21916 38752
rect 21871 38712 21916 38740
rect 21910 38700 21916 38712
rect 21968 38700 21974 38752
rect 26970 38700 26976 38752
rect 27028 38740 27034 38752
rect 27172 38749 27200 38916
rect 27985 38913 27997 38916
rect 28031 38913 28043 38947
rect 27985 38907 28043 38913
rect 28077 38947 28135 38953
rect 28077 38913 28089 38947
rect 28123 38913 28135 38947
rect 28077 38907 28135 38913
rect 28169 38947 28227 38953
rect 28169 38913 28181 38947
rect 28215 38913 28227 38947
rect 28169 38907 28227 38913
rect 28353 38947 28411 38953
rect 28353 38913 28365 38947
rect 28399 38944 28411 38947
rect 28442 38944 28448 38956
rect 28399 38916 28448 38944
rect 28399 38913 28411 38916
rect 28353 38907 28411 38913
rect 28092 38808 28120 38907
rect 28184 38876 28212 38907
rect 28442 38904 28448 38916
rect 28500 38904 28506 38956
rect 28994 38944 29000 38956
rect 28955 38916 29000 38944
rect 28994 38904 29000 38916
rect 29052 38904 29058 38956
rect 29914 38904 29920 38956
rect 29972 38944 29978 38956
rect 30466 38953 30472 38956
rect 30193 38947 30251 38953
rect 30193 38944 30205 38947
rect 29972 38916 30205 38944
rect 29972 38904 29978 38916
rect 30193 38913 30205 38916
rect 30239 38913 30251 38947
rect 30193 38907 30251 38913
rect 30460 38907 30472 38953
rect 30524 38944 30530 38956
rect 30524 38916 30560 38944
rect 30466 38904 30472 38907
rect 30524 38904 30530 38916
rect 31662 38904 31668 38956
rect 31720 38944 31726 38956
rect 32508 38953 32536 38984
rect 33134 38972 33140 38984
rect 33192 39012 33198 39024
rect 34057 39015 34115 39021
rect 33192 38984 33732 39012
rect 33192 38972 33198 38984
rect 32401 38947 32459 38953
rect 32401 38944 32413 38947
rect 31720 38916 32413 38944
rect 31720 38904 31726 38916
rect 32401 38913 32413 38916
rect 32447 38913 32459 38947
rect 32401 38907 32459 38913
rect 32493 38947 32551 38953
rect 32493 38913 32505 38947
rect 32539 38913 32551 38947
rect 32493 38907 32551 38913
rect 32582 38904 32588 38956
rect 32640 38944 32646 38956
rect 32769 38947 32827 38953
rect 32640 38916 32685 38944
rect 32640 38904 32646 38916
rect 32769 38913 32781 38947
rect 32815 38913 32827 38947
rect 32769 38907 32827 38913
rect 33413 38947 33471 38953
rect 33413 38913 33425 38947
rect 33459 38944 33471 38947
rect 33502 38944 33508 38956
rect 33459 38916 33508 38944
rect 33459 38913 33471 38916
rect 33413 38907 33471 38913
rect 28813 38879 28871 38885
rect 28813 38876 28825 38879
rect 28184 38848 28825 38876
rect 28813 38845 28825 38848
rect 28859 38845 28871 38879
rect 28813 38839 28871 38845
rect 30098 38808 30104 38820
rect 28092 38780 30104 38808
rect 30098 38768 30104 38780
rect 30156 38768 30162 38820
rect 32784 38808 32812 38907
rect 33502 38904 33508 38916
rect 33560 38904 33566 38956
rect 33704 38953 33732 38984
rect 34057 38981 34069 39015
rect 34103 39012 34115 39015
rect 35630 39015 35688 39021
rect 35630 39012 35642 39015
rect 34103 38984 35642 39012
rect 34103 38981 34115 38984
rect 34057 38975 34115 38981
rect 35630 38981 35642 38984
rect 35676 38981 35688 39015
rect 35630 38975 35688 38981
rect 33597 38947 33655 38953
rect 33597 38913 33609 38947
rect 33643 38913 33655 38947
rect 33597 38907 33655 38913
rect 33689 38947 33747 38953
rect 33689 38913 33701 38947
rect 33735 38913 33747 38947
rect 33689 38907 33747 38913
rect 33781 38947 33839 38953
rect 33781 38913 33793 38947
rect 33827 38944 33839 38947
rect 34514 38944 34520 38956
rect 33827 38916 34520 38944
rect 33827 38913 33839 38916
rect 33781 38907 33839 38913
rect 33612 38876 33640 38907
rect 34514 38904 34520 38916
rect 34572 38944 34578 38956
rect 35342 38944 35348 38956
rect 34572 38916 35348 38944
rect 34572 38904 34578 38916
rect 35342 38904 35348 38916
rect 35400 38904 35406 38956
rect 34790 38876 34796 38888
rect 33612 38848 34796 38876
rect 34790 38836 34796 38848
rect 34848 38836 34854 38888
rect 35897 38879 35955 38885
rect 35897 38845 35909 38879
rect 35943 38876 35955 38879
rect 36078 38876 36084 38888
rect 35943 38848 36084 38876
rect 35943 38845 35955 38848
rect 35897 38839 35955 38845
rect 36078 38836 36084 38848
rect 36136 38836 36142 38888
rect 58158 38808 58164 38820
rect 31128 38780 32812 38808
rect 58119 38780 58164 38808
rect 31128 38752 31156 38780
rect 58158 38768 58164 38780
rect 58216 38768 58222 38820
rect 27157 38743 27215 38749
rect 27157 38740 27169 38743
rect 27028 38712 27169 38740
rect 27028 38700 27034 38712
rect 27157 38709 27169 38712
rect 27203 38709 27215 38743
rect 27157 38703 27215 38709
rect 28442 38700 28448 38752
rect 28500 38740 28506 38752
rect 31110 38740 31116 38752
rect 28500 38712 31116 38740
rect 28500 38700 28506 38712
rect 31110 38700 31116 38712
rect 31168 38700 31174 38752
rect 31573 38743 31631 38749
rect 31573 38709 31585 38743
rect 31619 38740 31631 38743
rect 31938 38740 31944 38752
rect 31619 38712 31944 38740
rect 31619 38709 31631 38712
rect 31573 38703 31631 38709
rect 31938 38700 31944 38712
rect 31996 38700 32002 38752
rect 34517 38743 34575 38749
rect 34517 38709 34529 38743
rect 34563 38740 34575 38743
rect 34698 38740 34704 38752
rect 34563 38712 34704 38740
rect 34563 38709 34575 38712
rect 34517 38703 34575 38709
rect 34698 38700 34704 38712
rect 34756 38700 34762 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 9674 38496 9680 38548
rect 9732 38536 9738 38548
rect 9861 38539 9919 38545
rect 9861 38536 9873 38539
rect 9732 38508 9873 38536
rect 9732 38496 9738 38508
rect 9861 38505 9873 38508
rect 9907 38505 9919 38539
rect 13262 38536 13268 38548
rect 9861 38499 9919 38505
rect 11992 38508 13268 38536
rect 11992 38468 12020 38508
rect 13262 38496 13268 38508
rect 13320 38496 13326 38548
rect 13538 38496 13544 38548
rect 13596 38536 13602 38548
rect 19334 38536 19340 38548
rect 13596 38508 19340 38536
rect 13596 38496 13602 38508
rect 19334 38496 19340 38508
rect 19392 38496 19398 38548
rect 22554 38496 22560 38548
rect 22612 38536 22618 38548
rect 22833 38539 22891 38545
rect 22833 38536 22845 38539
rect 22612 38508 22845 38536
rect 22612 38496 22618 38508
rect 22833 38505 22845 38508
rect 22879 38505 22891 38539
rect 22833 38499 22891 38505
rect 23566 38496 23572 38548
rect 23624 38536 23630 38548
rect 24489 38539 24547 38545
rect 24489 38536 24501 38539
rect 23624 38508 24501 38536
rect 23624 38496 23630 38508
rect 24489 38505 24501 38508
rect 24535 38536 24547 38539
rect 30466 38536 30472 38548
rect 24535 38508 28304 38536
rect 30427 38508 30472 38536
rect 24535 38505 24547 38508
rect 24489 38499 24547 38505
rect 12158 38468 12164 38480
rect 7300 38440 12020 38468
rect 12119 38440 12164 38468
rect 6638 38360 6644 38412
rect 6696 38400 6702 38412
rect 7300 38409 7328 38440
rect 12158 38428 12164 38440
rect 12216 38428 12222 38480
rect 12268 38440 12756 38468
rect 7009 38403 7067 38409
rect 7009 38400 7021 38403
rect 6696 38372 7021 38400
rect 6696 38360 6702 38372
rect 7009 38369 7021 38372
rect 7055 38369 7067 38403
rect 7009 38363 7067 38369
rect 7285 38403 7343 38409
rect 7285 38369 7297 38403
rect 7331 38369 7343 38403
rect 9766 38400 9772 38412
rect 9679 38372 9772 38400
rect 7285 38363 7343 38369
rect 3786 38332 3792 38344
rect 3747 38304 3792 38332
rect 3786 38292 3792 38304
rect 3844 38292 3850 38344
rect 9692 38341 9720 38372
rect 9766 38360 9772 38372
rect 9824 38400 9830 38412
rect 12268 38400 12296 38440
rect 9824 38372 12296 38400
rect 12728 38400 12756 38440
rect 13630 38428 13636 38480
rect 13688 38468 13694 38480
rect 13688 38440 17356 38468
rect 13688 38428 13694 38440
rect 12728 38372 15240 38400
rect 9824 38360 9830 38372
rect 9677 38335 9735 38341
rect 9677 38301 9689 38335
rect 9723 38301 9735 38335
rect 10318 38332 10324 38344
rect 9677 38295 9735 38301
rect 9784 38304 10324 38332
rect 3878 38224 3884 38276
rect 3936 38264 3942 38276
rect 4034 38267 4092 38273
rect 4034 38264 4046 38267
rect 3936 38236 4046 38264
rect 3936 38224 3942 38236
rect 4034 38233 4046 38236
rect 4080 38233 4092 38267
rect 5813 38267 5871 38273
rect 5813 38264 5825 38267
rect 4034 38227 4092 38233
rect 5276 38236 5825 38264
rect 5276 38208 5304 38236
rect 5813 38233 5825 38236
rect 5859 38233 5871 38267
rect 5994 38264 6000 38276
rect 5955 38236 6000 38264
rect 5813 38227 5871 38233
rect 5994 38224 6000 38236
rect 6052 38224 6058 38276
rect 9493 38267 9551 38273
rect 9493 38233 9505 38267
rect 9539 38264 9551 38267
rect 9784 38264 9812 38304
rect 10318 38292 10324 38304
rect 10376 38292 10382 38344
rect 11977 38335 12035 38341
rect 11977 38301 11989 38335
rect 12023 38332 12035 38335
rect 12434 38332 12440 38344
rect 12023 38304 12440 38332
rect 12023 38301 12035 38304
rect 11977 38295 12035 38301
rect 12434 38292 12440 38304
rect 12492 38292 12498 38344
rect 12618 38332 12624 38344
rect 12579 38304 12624 38332
rect 12618 38292 12624 38304
rect 12676 38292 12682 38344
rect 12986 38332 12992 38344
rect 12947 38304 12992 38332
rect 12986 38292 12992 38304
rect 13044 38332 13050 38344
rect 15212 38341 15240 38372
rect 15378 38360 15384 38412
rect 15436 38360 15442 38412
rect 17328 38400 17356 38440
rect 17402 38428 17408 38480
rect 17460 38468 17466 38480
rect 18690 38468 18696 38480
rect 17460 38440 18696 38468
rect 17460 38428 17466 38440
rect 18690 38428 18696 38440
rect 18748 38428 18754 38480
rect 28276 38468 28304 38508
rect 30466 38496 30472 38508
rect 30524 38496 30530 38548
rect 32401 38539 32459 38545
rect 32401 38505 32413 38539
rect 32447 38536 32459 38539
rect 32582 38536 32588 38548
rect 32447 38508 32588 38536
rect 32447 38505 32459 38508
rect 32401 38499 32459 38505
rect 32582 38496 32588 38508
rect 32640 38496 32646 38548
rect 31662 38468 31668 38480
rect 28276 38440 31668 38468
rect 31662 38428 31668 38440
rect 31720 38428 31726 38480
rect 33502 38428 33508 38480
rect 33560 38428 33566 38480
rect 18322 38400 18328 38412
rect 17328 38372 18328 38400
rect 15197 38335 15255 38341
rect 13044 38304 15056 38332
rect 13044 38292 13050 38304
rect 12802 38264 12808 38276
rect 9539 38236 9812 38264
rect 12763 38236 12808 38264
rect 9539 38233 9551 38236
rect 9493 38227 9551 38233
rect 12802 38224 12808 38236
rect 12860 38224 12866 38276
rect 12897 38267 12955 38273
rect 12897 38233 12909 38267
rect 12943 38264 12955 38267
rect 13814 38264 13820 38276
rect 12943 38236 13820 38264
rect 12943 38233 12955 38236
rect 12897 38227 12955 38233
rect 13814 38224 13820 38236
rect 13872 38224 13878 38276
rect 3142 38196 3148 38208
rect 3103 38168 3148 38196
rect 3142 38156 3148 38168
rect 3200 38156 3206 38208
rect 5169 38199 5227 38205
rect 5169 38165 5181 38199
rect 5215 38196 5227 38199
rect 5258 38196 5264 38208
rect 5215 38168 5264 38196
rect 5215 38165 5227 38168
rect 5169 38159 5227 38165
rect 5258 38156 5264 38168
rect 5316 38156 5322 38208
rect 5534 38156 5540 38208
rect 5592 38196 5598 38208
rect 5629 38199 5687 38205
rect 5629 38196 5641 38199
rect 5592 38168 5641 38196
rect 5592 38156 5598 38168
rect 5629 38165 5641 38168
rect 5675 38165 5687 38199
rect 5629 38159 5687 38165
rect 9858 38156 9864 38208
rect 9916 38196 9922 38208
rect 12618 38196 12624 38208
rect 9916 38168 12624 38196
rect 9916 38156 9922 38168
rect 12618 38156 12624 38168
rect 12676 38156 12682 38208
rect 13173 38199 13231 38205
rect 13173 38165 13185 38199
rect 13219 38196 13231 38199
rect 13354 38196 13360 38208
rect 13219 38168 13360 38196
rect 13219 38165 13231 38168
rect 13173 38159 13231 38165
rect 13354 38156 13360 38168
rect 13412 38156 13418 38208
rect 15028 38196 15056 38304
rect 15197 38301 15209 38335
rect 15243 38301 15255 38335
rect 15396 38332 15424 38360
rect 17328 38341 17356 38372
rect 18322 38360 18328 38372
rect 18380 38360 18386 38412
rect 31941 38403 31999 38409
rect 31941 38400 31953 38403
rect 30944 38372 31953 38400
rect 15473 38335 15531 38341
rect 15473 38332 15485 38335
rect 15396 38304 15485 38332
rect 15197 38295 15255 38301
rect 15473 38301 15485 38304
rect 15519 38301 15531 38335
rect 15473 38295 15531 38301
rect 15565 38335 15623 38341
rect 15565 38301 15577 38335
rect 15611 38301 15623 38335
rect 17037 38335 17095 38341
rect 17037 38332 17049 38335
rect 15565 38295 15623 38301
rect 15764 38304 17049 38332
rect 15102 38224 15108 38276
rect 15160 38264 15166 38276
rect 15381 38267 15439 38273
rect 15381 38264 15393 38267
rect 15160 38236 15393 38264
rect 15160 38224 15166 38236
rect 15381 38233 15393 38236
rect 15427 38233 15439 38267
rect 15381 38227 15439 38233
rect 15470 38196 15476 38208
rect 15028 38168 15476 38196
rect 15470 38156 15476 38168
rect 15528 38196 15534 38208
rect 15580 38196 15608 38295
rect 15764 38205 15792 38304
rect 17037 38301 17049 38304
rect 17083 38301 17095 38335
rect 17037 38295 17095 38301
rect 17130 38335 17188 38341
rect 17130 38301 17142 38335
rect 17176 38301 17188 38335
rect 17130 38295 17188 38301
rect 17313 38335 17371 38341
rect 17313 38301 17325 38335
rect 17359 38301 17371 38335
rect 17313 38295 17371 38301
rect 17502 38335 17560 38341
rect 17502 38301 17514 38335
rect 17548 38332 17560 38335
rect 22646 38332 22652 38344
rect 17548 38304 17632 38332
rect 22607 38304 22652 38332
rect 17548 38301 17560 38304
rect 17502 38295 17560 38301
rect 15838 38224 15844 38276
rect 15896 38264 15902 38276
rect 17144 38264 17172 38295
rect 17402 38264 17408 38276
rect 15896 38236 17172 38264
rect 17363 38236 17408 38264
rect 15896 38224 15902 38236
rect 17402 38224 17408 38236
rect 17460 38224 17466 38276
rect 17604 38264 17632 38304
rect 22646 38292 22652 38304
rect 22704 38292 22710 38344
rect 25958 38292 25964 38344
rect 26016 38332 26022 38344
rect 30944 38341 30972 38372
rect 31941 38369 31953 38372
rect 31987 38369 31999 38403
rect 31941 38363 31999 38369
rect 33134 38360 33140 38412
rect 33192 38400 33198 38412
rect 33520 38400 33548 38428
rect 36078 38400 36084 38412
rect 33192 38372 33824 38400
rect 36039 38372 36084 38400
rect 33192 38360 33198 38372
rect 27341 38335 27399 38341
rect 27341 38332 27353 38335
rect 26016 38304 27353 38332
rect 26016 38292 26022 38304
rect 27341 38301 27353 38304
rect 27387 38301 27399 38335
rect 30745 38335 30803 38341
rect 30745 38332 30757 38335
rect 27341 38295 27399 38301
rect 29932 38304 30757 38332
rect 18598 38264 18604 38276
rect 17604 38236 18604 38264
rect 15528 38168 15608 38196
rect 15749 38199 15807 38205
rect 15528 38156 15534 38168
rect 15749 38165 15761 38199
rect 15795 38165 15807 38199
rect 15749 38159 15807 38165
rect 16482 38156 16488 38208
rect 16540 38196 16546 38208
rect 17604 38196 17632 38236
rect 18598 38224 18604 38236
rect 18656 38264 18662 38276
rect 18966 38264 18972 38276
rect 18656 38236 18972 38264
rect 18656 38224 18662 38236
rect 18966 38224 18972 38236
rect 19024 38224 19030 38276
rect 22094 38224 22100 38276
rect 22152 38264 22158 38276
rect 22465 38267 22523 38273
rect 22465 38264 22477 38267
rect 22152 38236 22477 38264
rect 22152 38224 22158 38236
rect 22465 38233 22477 38236
rect 22511 38264 22523 38267
rect 22830 38264 22836 38276
rect 22511 38236 22836 38264
rect 22511 38233 22523 38236
rect 22465 38227 22523 38233
rect 22830 38224 22836 38236
rect 22888 38224 22894 38276
rect 27608 38267 27666 38273
rect 27608 38233 27620 38267
rect 27654 38264 27666 38267
rect 27706 38264 27712 38276
rect 27654 38236 27712 38264
rect 27654 38233 27666 38236
rect 27608 38227 27666 38233
rect 27706 38224 27712 38236
rect 27764 38224 27770 38276
rect 29932 38208 29960 38304
rect 30745 38301 30757 38304
rect 30791 38301 30803 38335
rect 30745 38295 30803 38301
rect 30837 38335 30895 38341
rect 30837 38301 30849 38335
rect 30883 38301 30895 38335
rect 30837 38295 30895 38301
rect 30929 38335 30987 38341
rect 30929 38301 30941 38335
rect 30975 38301 30987 38335
rect 31110 38332 31116 38344
rect 31071 38304 31116 38332
rect 30929 38295 30987 38301
rect 30098 38224 30104 38276
rect 30156 38264 30162 38276
rect 30852 38264 30880 38295
rect 31110 38292 31116 38304
rect 31168 38292 31174 38344
rect 32585 38335 32643 38341
rect 32585 38301 32597 38335
rect 32631 38332 32643 38335
rect 33226 38332 33232 38344
rect 32631 38304 33232 38332
rect 32631 38301 32643 38304
rect 32585 38295 32643 38301
rect 33226 38292 33232 38304
rect 33284 38292 33290 38344
rect 33505 38335 33563 38341
rect 33505 38301 33517 38335
rect 33551 38301 33563 38335
rect 33686 38332 33692 38344
rect 33647 38304 33692 38332
rect 33505 38295 33563 38301
rect 30156 38236 30880 38264
rect 30156 38224 30162 38236
rect 31202 38224 31208 38276
rect 31260 38264 31266 38276
rect 31573 38267 31631 38273
rect 31573 38264 31585 38267
rect 31260 38236 31585 38264
rect 31260 38224 31266 38236
rect 31573 38233 31585 38236
rect 31619 38233 31631 38267
rect 31573 38227 31631 38233
rect 31757 38267 31815 38273
rect 31757 38233 31769 38267
rect 31803 38264 31815 38267
rect 31938 38264 31944 38276
rect 31803 38236 31944 38264
rect 31803 38233 31815 38236
rect 31757 38227 31815 38233
rect 31938 38224 31944 38236
rect 31996 38264 32002 38276
rect 32674 38264 32680 38276
rect 31996 38236 32680 38264
rect 31996 38224 32002 38236
rect 32674 38224 32680 38236
rect 32732 38224 32738 38276
rect 32769 38267 32827 38273
rect 32769 38233 32781 38267
rect 32815 38264 32827 38267
rect 33410 38264 33416 38276
rect 32815 38236 33416 38264
rect 32815 38233 32827 38236
rect 32769 38227 32827 38233
rect 33410 38224 33416 38236
rect 33468 38224 33474 38276
rect 33520 38264 33548 38295
rect 33686 38292 33692 38304
rect 33744 38292 33750 38344
rect 33796 38341 33824 38372
rect 36078 38360 36084 38372
rect 36136 38360 36142 38412
rect 33781 38335 33839 38341
rect 33781 38301 33793 38335
rect 33827 38301 33839 38335
rect 33781 38295 33839 38301
rect 33919 38335 33977 38341
rect 33919 38301 33931 38335
rect 33965 38332 33977 38335
rect 34514 38332 34520 38344
rect 33965 38304 34520 38332
rect 33965 38301 33977 38304
rect 33919 38295 33977 38301
rect 34514 38292 34520 38304
rect 34572 38292 34578 38344
rect 33594 38264 33600 38276
rect 33520 38236 33600 38264
rect 33594 38224 33600 38236
rect 33652 38224 33658 38276
rect 34149 38267 34207 38273
rect 34149 38233 34161 38267
rect 34195 38264 34207 38267
rect 35814 38267 35872 38273
rect 35814 38264 35826 38267
rect 34195 38236 35826 38264
rect 34195 38233 34207 38236
rect 34149 38227 34207 38233
rect 35814 38233 35826 38236
rect 35860 38233 35872 38267
rect 35814 38227 35872 38233
rect 16540 38168 17632 38196
rect 17681 38199 17739 38205
rect 16540 38156 16546 38168
rect 17681 38165 17693 38199
rect 17727 38196 17739 38199
rect 18506 38196 18512 38208
rect 17727 38168 18512 38196
rect 17727 38165 17739 38168
rect 17681 38159 17739 38165
rect 18506 38156 18512 38168
rect 18564 38156 18570 38208
rect 19334 38156 19340 38208
rect 19392 38196 19398 38208
rect 19429 38199 19487 38205
rect 19429 38196 19441 38199
rect 19392 38168 19441 38196
rect 19392 38156 19398 38168
rect 19429 38165 19441 38168
rect 19475 38165 19487 38199
rect 19429 38159 19487 38165
rect 28721 38199 28779 38205
rect 28721 38165 28733 38199
rect 28767 38196 28779 38199
rect 28994 38196 29000 38208
rect 28767 38168 29000 38196
rect 28767 38165 28779 38168
rect 28721 38159 28779 38165
rect 28994 38156 29000 38168
rect 29052 38156 29058 38208
rect 29914 38196 29920 38208
rect 29875 38168 29920 38196
rect 29914 38156 29920 38168
rect 29972 38156 29978 38208
rect 34054 38156 34060 38208
rect 34112 38196 34118 38208
rect 34701 38199 34759 38205
rect 34701 38196 34713 38199
rect 34112 38168 34713 38196
rect 34112 38156 34118 38168
rect 34701 38165 34713 38168
rect 34747 38165 34759 38199
rect 34701 38159 34759 38165
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 2590 37952 2596 38004
rect 2648 37952 2654 38004
rect 15102 37992 15108 38004
rect 12820 37964 15108 37992
rect 2608 37924 2636 37952
rect 12820 37936 12848 37964
rect 15102 37952 15108 37964
rect 15160 37992 15166 38004
rect 15657 37995 15715 38001
rect 15160 37964 15249 37992
rect 15160 37952 15166 37964
rect 2608 37896 2728 37924
rect 2700 37865 2728 37896
rect 6362 37884 6368 37936
rect 6420 37924 6426 37936
rect 7469 37927 7527 37933
rect 6420 37896 7420 37924
rect 6420 37884 6426 37896
rect 2593 37859 2651 37865
rect 2593 37825 2605 37859
rect 2639 37825 2651 37859
rect 2593 37819 2651 37825
rect 2685 37859 2743 37865
rect 2685 37825 2697 37859
rect 2731 37825 2743 37859
rect 2685 37819 2743 37825
rect 2777 37859 2835 37865
rect 2777 37825 2789 37859
rect 2823 37856 2835 37859
rect 2866 37856 2872 37868
rect 2823 37828 2872 37856
rect 2823 37825 2835 37828
rect 2777 37819 2835 37825
rect 2608 37788 2636 37819
rect 2866 37816 2872 37828
rect 2924 37816 2930 37868
rect 2961 37859 3019 37865
rect 2961 37825 2973 37859
rect 3007 37856 3019 37859
rect 3234 37856 3240 37868
rect 3007 37828 3240 37856
rect 3007 37825 3019 37828
rect 2961 37819 3019 37825
rect 3234 37816 3240 37828
rect 3292 37856 3298 37868
rect 4614 37856 4620 37868
rect 3292 37828 4620 37856
rect 3292 37816 3298 37828
rect 4614 37816 4620 37828
rect 4672 37816 4678 37868
rect 5169 37859 5227 37865
rect 5169 37825 5181 37859
rect 5215 37856 5227 37859
rect 5718 37856 5724 37868
rect 5215 37828 5724 37856
rect 5215 37825 5227 37828
rect 5169 37819 5227 37825
rect 5718 37816 5724 37828
rect 5776 37816 5782 37868
rect 6822 37816 6828 37868
rect 6880 37856 6886 37868
rect 7285 37859 7343 37865
rect 7285 37856 7297 37859
rect 6880 37828 7297 37856
rect 6880 37816 6886 37828
rect 7285 37825 7297 37828
rect 7331 37825 7343 37859
rect 7392 37856 7420 37896
rect 7469 37893 7481 37927
rect 7515 37924 7527 37927
rect 8481 37927 8539 37933
rect 8481 37924 8493 37927
rect 7515 37896 8493 37924
rect 7515 37893 7527 37896
rect 7469 37887 7527 37893
rect 8481 37893 8493 37896
rect 8527 37924 8539 37927
rect 11974 37924 11980 37936
rect 8527 37896 11980 37924
rect 8527 37893 8539 37896
rect 8481 37887 8539 37893
rect 11974 37884 11980 37896
rect 12032 37924 12038 37936
rect 12802 37924 12808 37936
rect 12032 37896 12808 37924
rect 12032 37884 12038 37896
rect 12802 37884 12808 37896
rect 12860 37884 12866 37936
rect 7561 37859 7619 37865
rect 7561 37856 7573 37859
rect 7392 37828 7573 37856
rect 7285 37819 7343 37825
rect 7561 37825 7573 37828
rect 7607 37825 7619 37859
rect 7561 37819 7619 37825
rect 7653 37859 7711 37865
rect 7653 37825 7665 37859
rect 7699 37825 7711 37859
rect 8294 37856 8300 37868
rect 8255 37828 8300 37856
rect 7653 37819 7711 37825
rect 3142 37788 3148 37800
rect 2608 37760 3148 37788
rect 3142 37748 3148 37760
rect 3200 37748 3206 37800
rect 3421 37791 3479 37797
rect 3421 37757 3433 37791
rect 3467 37788 3479 37791
rect 3786 37788 3792 37800
rect 3467 37760 3792 37788
rect 3467 37757 3479 37760
rect 3421 37751 3479 37757
rect 2774 37680 2780 37732
rect 2832 37720 2838 37732
rect 3436 37720 3464 37751
rect 3786 37748 3792 37760
rect 3844 37748 3850 37800
rect 7668 37788 7696 37819
rect 8294 37816 8300 37828
rect 8352 37816 8358 37868
rect 8570 37856 8576 37868
rect 8531 37828 8576 37856
rect 8570 37816 8576 37828
rect 8628 37816 8634 37868
rect 8665 37859 8723 37865
rect 8665 37825 8677 37859
rect 8711 37856 8723 37859
rect 12253 37859 12311 37865
rect 12253 37856 12265 37859
rect 8711 37828 12265 37856
rect 8711 37825 8723 37828
rect 8665 37819 8723 37825
rect 12253 37825 12265 37828
rect 12299 37856 12311 37859
rect 12986 37856 12992 37868
rect 12299 37828 12992 37856
rect 12299 37825 12311 37828
rect 12253 37819 12311 37825
rect 8680 37788 8708 37819
rect 12986 37816 12992 37828
rect 13044 37816 13050 37868
rect 13354 37856 13360 37868
rect 13315 37828 13360 37856
rect 13354 37816 13360 37828
rect 13412 37816 13418 37868
rect 13446 37816 13452 37868
rect 13504 37856 13510 37868
rect 13630 37856 13636 37868
rect 13504 37828 13549 37856
rect 13591 37828 13636 37856
rect 13504 37816 13510 37828
rect 13630 37816 13636 37828
rect 13688 37816 13694 37868
rect 13725 37859 13783 37865
rect 13725 37825 13737 37859
rect 13771 37825 13783 37859
rect 13725 37819 13783 37825
rect 13822 37859 13880 37865
rect 13822 37825 13834 37859
rect 13868 37856 13880 37859
rect 13868 37828 13952 37856
rect 13868 37825 13880 37828
rect 13822 37819 13880 37825
rect 7668 37760 8708 37788
rect 12529 37791 12587 37797
rect 12529 37757 12541 37791
rect 12575 37788 12587 37791
rect 12802 37788 12808 37800
rect 12575 37760 12808 37788
rect 12575 37757 12587 37760
rect 12529 37751 12587 37757
rect 12802 37748 12808 37760
rect 12860 37748 12866 37800
rect 13538 37748 13544 37800
rect 13596 37788 13602 37800
rect 13740 37788 13768 37819
rect 13596 37760 13768 37788
rect 13924 37788 13952 37828
rect 13998 37816 14004 37868
rect 14056 37856 14062 37868
rect 15221 37865 15249 37964
rect 15657 37961 15669 37995
rect 15703 37961 15715 37995
rect 15657 37955 15715 37961
rect 15381 37927 15439 37933
rect 15381 37893 15393 37927
rect 15427 37924 15439 37927
rect 15562 37924 15568 37936
rect 15427 37896 15568 37924
rect 15427 37893 15439 37896
rect 15381 37887 15439 37893
rect 15562 37884 15568 37896
rect 15620 37884 15626 37936
rect 15672 37924 15700 37955
rect 18782 37952 18788 38004
rect 18840 37992 18846 38004
rect 18840 37964 18920 37992
rect 18840 37952 18846 37964
rect 18892 37933 18920 37964
rect 20438 37952 20444 38004
rect 20496 37992 20502 38004
rect 20717 37995 20775 38001
rect 20717 37992 20729 37995
rect 20496 37964 20729 37992
rect 20496 37952 20502 37964
rect 20717 37961 20729 37964
rect 20763 37961 20775 37995
rect 20717 37955 20775 37961
rect 33686 37952 33692 38004
rect 33744 37992 33750 38004
rect 33781 37995 33839 38001
rect 33781 37992 33793 37995
rect 33744 37964 33793 37992
rect 33744 37952 33750 37964
rect 33781 37961 33793 37964
rect 33827 37961 33839 37995
rect 33781 37955 33839 37961
rect 34790 37952 34796 38004
rect 34848 37992 34854 38004
rect 34977 37995 35035 38001
rect 34977 37992 34989 37995
rect 34848 37964 34989 37992
rect 34848 37952 34854 37964
rect 34977 37961 34989 37964
rect 35023 37961 35035 37995
rect 34977 37955 35035 37961
rect 18877 37927 18935 37933
rect 15672 37896 18552 37924
rect 15105 37859 15163 37865
rect 15105 37856 15117 37859
rect 14056 37828 15117 37856
rect 14056 37816 14062 37828
rect 15105 37825 15117 37828
rect 15151 37825 15163 37859
rect 15221 37859 15301 37865
rect 15221 37828 15255 37859
rect 15105 37819 15163 37825
rect 15243 37825 15255 37828
rect 15289 37825 15301 37859
rect 15470 37856 15476 37868
rect 15431 37828 15476 37856
rect 15243 37819 15301 37825
rect 15470 37816 15476 37828
rect 15528 37816 15534 37868
rect 16758 37816 16764 37868
rect 16816 37856 16822 37868
rect 18524 37865 18552 37896
rect 18877 37893 18889 37927
rect 18923 37893 18935 37927
rect 18877 37887 18935 37893
rect 16925 37859 16983 37865
rect 16925 37856 16937 37859
rect 16816 37828 16937 37856
rect 16816 37816 16822 37828
rect 16925 37825 16937 37828
rect 16971 37825 16983 37859
rect 16925 37819 16983 37825
rect 18509 37859 18567 37865
rect 18509 37825 18521 37859
rect 18555 37825 18567 37859
rect 18509 37819 18567 37825
rect 18602 37859 18660 37865
rect 18602 37825 18614 37859
rect 18648 37825 18660 37859
rect 18602 37819 18660 37825
rect 18785 37859 18843 37865
rect 18785 37825 18797 37859
rect 18831 37825 18843 37859
rect 18785 37819 18843 37825
rect 13924 37760 14044 37788
rect 13596 37748 13602 37760
rect 2832 37692 3464 37720
rect 2832 37680 2838 37692
rect 10594 37680 10600 37732
rect 10652 37720 10658 37732
rect 13906 37720 13912 37732
rect 10652 37692 13912 37720
rect 10652 37680 10658 37692
rect 13906 37680 13912 37692
rect 13964 37680 13970 37732
rect 14016 37720 14044 37760
rect 14090 37748 14096 37800
rect 14148 37788 14154 37800
rect 14918 37788 14924 37800
rect 14148 37760 14924 37788
rect 14148 37748 14154 37760
rect 14918 37748 14924 37760
rect 14976 37788 14982 37800
rect 16669 37791 16727 37797
rect 16669 37788 16681 37791
rect 14976 37760 16681 37788
rect 14976 37748 14982 37760
rect 16669 37757 16681 37760
rect 16715 37757 16727 37791
rect 18616 37788 18644 37819
rect 16669 37751 16727 37757
rect 18064 37760 18644 37788
rect 15194 37720 15200 37732
rect 14016 37692 15200 37720
rect 15194 37680 15200 37692
rect 15252 37720 15258 37732
rect 16482 37720 16488 37732
rect 15252 37692 16488 37720
rect 15252 37680 15258 37692
rect 16482 37680 16488 37692
rect 16540 37680 16546 37732
rect 2314 37652 2320 37664
rect 2275 37624 2320 37652
rect 2314 37612 2320 37624
rect 2372 37612 2378 37664
rect 5718 37652 5724 37664
rect 5679 37624 5724 37652
rect 5718 37612 5724 37624
rect 5776 37612 5782 37664
rect 7837 37655 7895 37661
rect 7837 37621 7849 37655
rect 7883 37652 7895 37655
rect 8662 37652 8668 37664
rect 7883 37624 8668 37652
rect 7883 37621 7895 37624
rect 7837 37615 7895 37621
rect 8662 37612 8668 37624
rect 8720 37612 8726 37664
rect 8849 37655 8907 37661
rect 8849 37621 8861 37655
rect 8895 37652 8907 37655
rect 8938 37652 8944 37664
rect 8895 37624 8944 37652
rect 8895 37621 8907 37624
rect 8849 37615 8907 37621
rect 8938 37612 8944 37624
rect 8996 37612 9002 37664
rect 14001 37655 14059 37661
rect 14001 37621 14013 37655
rect 14047 37652 14059 37655
rect 14458 37652 14464 37664
rect 14047 37624 14464 37652
rect 14047 37621 14059 37624
rect 14001 37615 14059 37621
rect 14458 37612 14464 37624
rect 14516 37612 14522 37664
rect 17954 37612 17960 37664
rect 18012 37652 18018 37664
rect 18064 37661 18092 37760
rect 18322 37680 18328 37732
rect 18380 37720 18386 37732
rect 18800 37720 18828 37819
rect 18966 37816 18972 37868
rect 19024 37865 19030 37868
rect 19024 37856 19032 37865
rect 19024 37828 19069 37856
rect 19024 37819 19032 37828
rect 19024 37816 19030 37819
rect 19334 37816 19340 37868
rect 19392 37856 19398 37868
rect 19613 37859 19671 37865
rect 19613 37856 19625 37859
rect 19392 37828 19625 37856
rect 19392 37816 19398 37828
rect 19613 37825 19625 37828
rect 19659 37825 19671 37859
rect 19794 37856 19800 37868
rect 19755 37828 19800 37856
rect 19613 37819 19671 37825
rect 19794 37816 19800 37828
rect 19852 37816 19858 37868
rect 19889 37859 19947 37865
rect 19889 37825 19901 37859
rect 19935 37825 19947 37859
rect 19889 37819 19947 37825
rect 19981 37859 20039 37865
rect 19981 37825 19993 37859
rect 20027 37856 20039 37859
rect 20456 37856 20484 37952
rect 33410 37884 33416 37936
rect 33468 37924 33474 37936
rect 34149 37927 34207 37933
rect 34149 37924 34161 37927
rect 33468 37896 34161 37924
rect 33468 37884 33474 37896
rect 34149 37893 34161 37896
rect 34195 37924 34207 37927
rect 34609 37927 34667 37933
rect 34609 37924 34621 37927
rect 34195 37896 34621 37924
rect 34195 37893 34207 37896
rect 34149 37887 34207 37893
rect 34609 37893 34621 37896
rect 34655 37893 34667 37927
rect 34609 37887 34667 37893
rect 24210 37856 24216 37868
rect 20027 37828 24216 37856
rect 20027 37825 20039 37828
rect 19981 37819 20039 37825
rect 19904 37788 19932 37819
rect 24210 37816 24216 37828
rect 24268 37816 24274 37868
rect 25130 37816 25136 37868
rect 25188 37856 25194 37868
rect 25694 37859 25752 37865
rect 25694 37856 25706 37859
rect 25188 37828 25706 37856
rect 25188 37816 25194 37828
rect 25694 37825 25706 37828
rect 25740 37825 25752 37859
rect 25694 37819 25752 37825
rect 31021 37859 31079 37865
rect 31021 37825 31033 37859
rect 31067 37856 31079 37859
rect 31110 37856 31116 37868
rect 31067 37828 31116 37856
rect 31067 37825 31079 37828
rect 31021 37819 31079 37825
rect 31110 37816 31116 37828
rect 31168 37816 31174 37868
rect 32585 37859 32643 37865
rect 32585 37825 32597 37859
rect 32631 37825 32643 37859
rect 32585 37819 32643 37825
rect 33965 37859 34023 37865
rect 33965 37825 33977 37859
rect 34011 37856 34023 37859
rect 34054 37856 34060 37868
rect 34011 37828 34060 37856
rect 34011 37825 34023 37828
rect 33965 37819 34023 37825
rect 25958 37788 25964 37800
rect 19904 37760 20024 37788
rect 25919 37760 25964 37788
rect 19996 37732 20024 37760
rect 25958 37748 25964 37760
rect 26016 37748 26022 37800
rect 31297 37791 31355 37797
rect 31297 37788 31309 37791
rect 29932 37760 31309 37788
rect 18380 37692 18828 37720
rect 18380 37680 18386 37692
rect 19978 37680 19984 37732
rect 20036 37680 20042 37732
rect 20257 37723 20315 37729
rect 20257 37689 20269 37723
rect 20303 37720 20315 37723
rect 21174 37720 21180 37732
rect 20303 37692 21180 37720
rect 20303 37689 20315 37692
rect 20257 37683 20315 37689
rect 21174 37680 21180 37692
rect 21232 37680 21238 37732
rect 18049 37655 18107 37661
rect 18049 37652 18061 37655
rect 18012 37624 18061 37652
rect 18012 37612 18018 37624
rect 18049 37621 18061 37624
rect 18095 37621 18107 37655
rect 18049 37615 18107 37621
rect 18782 37612 18788 37664
rect 18840 37652 18846 37664
rect 19153 37655 19211 37661
rect 19153 37652 19165 37655
rect 18840 37624 19165 37652
rect 18840 37612 18846 37624
rect 19153 37621 19165 37624
rect 19199 37621 19211 37655
rect 19153 37615 19211 37621
rect 23569 37655 23627 37661
rect 23569 37621 23581 37655
rect 23615 37652 23627 37655
rect 24026 37652 24032 37664
rect 23615 37624 24032 37652
rect 23615 37621 23627 37624
rect 23569 37615 23627 37621
rect 24026 37612 24032 37624
rect 24084 37612 24090 37664
rect 24486 37612 24492 37664
rect 24544 37652 24550 37664
rect 24581 37655 24639 37661
rect 24581 37652 24593 37655
rect 24544 37624 24593 37652
rect 24544 37612 24550 37624
rect 24581 37621 24593 37624
rect 24627 37621 24639 37655
rect 24581 37615 24639 37621
rect 29822 37612 29828 37664
rect 29880 37652 29886 37664
rect 29932 37661 29960 37760
rect 31297 37757 31309 37760
rect 31343 37788 31355 37791
rect 32306 37788 32312 37800
rect 31343 37760 32312 37788
rect 31343 37757 31355 37760
rect 31297 37751 31355 37757
rect 32306 37748 32312 37760
rect 32364 37788 32370 37800
rect 32600 37788 32628 37819
rect 34054 37816 34060 37828
rect 34112 37816 34118 37868
rect 34698 37816 34704 37868
rect 34756 37856 34762 37868
rect 34793 37859 34851 37865
rect 34793 37856 34805 37859
rect 34756 37828 34805 37856
rect 34756 37816 34762 37828
rect 34793 37825 34805 37828
rect 34839 37825 34851 37859
rect 34793 37819 34851 37825
rect 32364 37760 32628 37788
rect 32364 37748 32370 37760
rect 32769 37723 32827 37729
rect 32769 37689 32781 37723
rect 32815 37720 32827 37723
rect 33594 37720 33600 37732
rect 32815 37692 33600 37720
rect 32815 37689 32827 37692
rect 32769 37683 32827 37689
rect 33594 37680 33600 37692
rect 33652 37680 33658 37732
rect 29917 37655 29975 37661
rect 29917 37652 29929 37655
rect 29880 37624 29929 37652
rect 29880 37612 29886 37624
rect 29917 37621 29929 37624
rect 29963 37621 29975 37655
rect 29917 37615 29975 37621
rect 33321 37655 33379 37661
rect 33321 37621 33333 37655
rect 33367 37652 33379 37655
rect 34514 37652 34520 37664
rect 33367 37624 34520 37652
rect 33367 37621 33379 37624
rect 33321 37615 33379 37621
rect 34514 37612 34520 37624
rect 34572 37652 34578 37664
rect 35526 37652 35532 37664
rect 34572 37624 35532 37652
rect 34572 37612 34578 37624
rect 35526 37612 35532 37624
rect 35584 37612 35590 37664
rect 58158 37652 58164 37664
rect 58119 37624 58164 37652
rect 58158 37612 58164 37624
rect 58216 37612 58222 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 2590 37408 2596 37460
rect 2648 37448 2654 37460
rect 3789 37451 3847 37457
rect 2648 37420 3464 37448
rect 2648 37408 2654 37420
rect 3436 37380 3464 37420
rect 3789 37417 3801 37451
rect 3835 37448 3847 37451
rect 3878 37448 3884 37460
rect 3835 37420 3884 37448
rect 3835 37417 3847 37420
rect 3789 37411 3847 37417
rect 3878 37408 3884 37420
rect 3936 37408 3942 37460
rect 15473 37451 15531 37457
rect 15473 37417 15485 37451
rect 15519 37448 15531 37451
rect 15838 37448 15844 37460
rect 15519 37420 15844 37448
rect 15519 37417 15531 37420
rect 15473 37411 15531 37417
rect 15838 37408 15844 37420
rect 15896 37408 15902 37460
rect 19613 37451 19671 37457
rect 19613 37417 19625 37451
rect 19659 37448 19671 37451
rect 19794 37448 19800 37460
rect 19659 37420 19800 37448
rect 19659 37417 19671 37420
rect 19613 37411 19671 37417
rect 19794 37408 19800 37420
rect 19852 37408 19858 37460
rect 24670 37448 24676 37460
rect 23492 37420 24676 37448
rect 3436 37352 4200 37380
rect 4172 37253 4200 37352
rect 11974 37312 11980 37324
rect 4264 37284 4568 37312
rect 11935 37284 11980 37312
rect 4264 37253 4292 37284
rect 1857 37247 1915 37253
rect 1857 37213 1869 37247
rect 1903 37244 1915 37247
rect 4065 37247 4123 37253
rect 4065 37244 4077 37247
rect 1903 37216 2774 37244
rect 1903 37213 1915 37216
rect 1857 37207 1915 37213
rect 2746 37188 2774 37216
rect 3988 37216 4077 37244
rect 2124 37179 2182 37185
rect 2124 37145 2136 37179
rect 2170 37176 2182 37179
rect 2314 37176 2320 37188
rect 2170 37148 2320 37176
rect 2170 37145 2182 37148
rect 2124 37139 2182 37145
rect 2314 37136 2320 37148
rect 2372 37136 2378 37188
rect 2746 37148 2780 37188
rect 2774 37136 2780 37148
rect 2832 37136 2838 37188
rect 3988 37176 4016 37216
rect 4065 37213 4077 37216
rect 4111 37213 4123 37247
rect 4065 37207 4123 37213
rect 4157 37247 4215 37253
rect 4157 37213 4169 37247
rect 4203 37213 4215 37247
rect 4157 37207 4215 37213
rect 4249 37247 4307 37253
rect 4249 37213 4261 37247
rect 4295 37213 4307 37247
rect 4430 37244 4436 37256
rect 4391 37216 4436 37244
rect 4249 37207 4307 37213
rect 4430 37204 4436 37216
rect 4488 37204 4494 37256
rect 4540 37244 4568 37284
rect 11974 37272 11980 37284
rect 12032 37272 12038 37324
rect 14090 37312 14096 37324
rect 14051 37284 14096 37312
rect 14090 37272 14096 37284
rect 14148 37272 14154 37324
rect 17954 37312 17960 37324
rect 17880 37284 17960 37312
rect 5350 37244 5356 37256
rect 4540 37216 5356 37244
rect 5350 37204 5356 37216
rect 5408 37204 5414 37256
rect 5445 37247 5503 37253
rect 5445 37213 5457 37247
rect 5491 37213 5503 37247
rect 5445 37207 5503 37213
rect 10229 37247 10287 37253
rect 10229 37213 10241 37247
rect 10275 37244 10287 37247
rect 10318 37244 10324 37256
rect 10275 37216 10324 37244
rect 10275 37213 10287 37216
rect 10229 37207 10287 37213
rect 4982 37176 4988 37188
rect 3988 37148 4988 37176
rect 4982 37136 4988 37148
rect 5040 37136 5046 37188
rect 3050 37068 3056 37120
rect 3108 37108 3114 37120
rect 3237 37111 3295 37117
rect 3237 37108 3249 37111
rect 3108 37080 3249 37108
rect 3108 37068 3114 37080
rect 3237 37077 3249 37080
rect 3283 37077 3295 37111
rect 3237 37071 3295 37077
rect 3786 37068 3792 37120
rect 3844 37108 3850 37120
rect 5460 37108 5488 37207
rect 10318 37204 10324 37216
rect 10376 37204 10382 37256
rect 12253 37247 12311 37253
rect 12253 37213 12265 37247
rect 12299 37244 12311 37247
rect 12618 37244 12624 37256
rect 12299 37216 12624 37244
rect 12299 37213 12311 37216
rect 12253 37207 12311 37213
rect 12618 37204 12624 37216
rect 12676 37204 12682 37256
rect 16761 37247 16819 37253
rect 16761 37213 16773 37247
rect 16807 37244 16819 37247
rect 17880 37244 17908 37284
rect 17954 37272 17960 37284
rect 18012 37272 18018 37324
rect 18432 37284 18736 37312
rect 18046 37244 18052 37256
rect 16807 37216 17908 37244
rect 18007 37216 18052 37244
rect 16807 37213 16819 37216
rect 16761 37207 16819 37213
rect 18046 37204 18052 37216
rect 18104 37204 18110 37256
rect 18197 37247 18255 37253
rect 18197 37213 18209 37247
rect 18243 37244 18255 37247
rect 18432 37244 18460 37284
rect 18708 37256 18736 37284
rect 18598 37253 18604 37256
rect 18243 37216 18460 37244
rect 18555 37247 18604 37253
rect 18243 37213 18255 37216
rect 18197 37207 18255 37213
rect 18555 37213 18567 37247
rect 18601 37213 18604 37247
rect 18555 37207 18604 37213
rect 18598 37204 18604 37207
rect 18656 37204 18662 37256
rect 18690 37204 18696 37256
rect 18748 37204 18754 37256
rect 19150 37204 19156 37256
rect 19208 37244 19214 37256
rect 19245 37247 19303 37253
rect 19245 37244 19257 37247
rect 19208 37216 19257 37244
rect 19208 37204 19214 37216
rect 19245 37213 19257 37216
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 21453 37247 21511 37253
rect 21453 37244 21465 37247
rect 20772 37216 21465 37244
rect 20772 37204 20778 37216
rect 21453 37213 21465 37216
rect 21499 37213 21511 37247
rect 21453 37207 21511 37213
rect 23201 37247 23259 37253
rect 23201 37213 23213 37247
rect 23247 37213 23259 37247
rect 23382 37244 23388 37256
rect 23343 37216 23388 37244
rect 23201 37207 23259 37213
rect 5712 37179 5770 37185
rect 5712 37145 5724 37179
rect 5758 37145 5770 37179
rect 10410 37176 10416 37188
rect 10371 37148 10416 37176
rect 5712 37139 5770 37145
rect 3844 37080 5488 37108
rect 3844 37068 3850 37080
rect 5626 37068 5632 37120
rect 5684 37108 5690 37120
rect 5736 37108 5764 37139
rect 10410 37136 10416 37148
rect 10468 37136 10474 37188
rect 14090 37136 14096 37188
rect 14148 37176 14154 37188
rect 14338 37179 14396 37185
rect 14338 37176 14350 37179
rect 14148 37148 14350 37176
rect 14148 37136 14154 37148
rect 14338 37145 14350 37148
rect 14384 37145 14396 37179
rect 16942 37176 16948 37188
rect 16903 37148 16948 37176
rect 14338 37139 14396 37145
rect 16942 37136 16948 37148
rect 17000 37136 17006 37188
rect 18322 37176 18328 37188
rect 18283 37148 18328 37176
rect 18322 37136 18328 37148
rect 18380 37136 18386 37188
rect 18417 37179 18475 37185
rect 18417 37145 18429 37179
rect 18463 37176 18475 37179
rect 19429 37179 19487 37185
rect 18463 37148 19196 37176
rect 18463 37145 18475 37148
rect 18417 37139 18475 37145
rect 5684 37080 5764 37108
rect 5684 37068 5690 37080
rect 6178 37068 6184 37120
rect 6236 37108 6242 37120
rect 6822 37108 6828 37120
rect 6236 37080 6828 37108
rect 6236 37068 6242 37080
rect 6822 37068 6828 37080
rect 6880 37068 6886 37120
rect 10594 37108 10600 37120
rect 10555 37080 10600 37108
rect 10594 37068 10600 37080
rect 10652 37068 10658 37120
rect 16206 37068 16212 37120
rect 16264 37108 16270 37120
rect 16577 37111 16635 37117
rect 16577 37108 16589 37111
rect 16264 37080 16589 37108
rect 16264 37068 16270 37080
rect 16577 37077 16589 37080
rect 16623 37077 16635 37111
rect 16577 37071 16635 37077
rect 18598 37068 18604 37120
rect 18656 37108 18662 37120
rect 18693 37111 18751 37117
rect 18693 37108 18705 37111
rect 18656 37080 18705 37108
rect 18656 37068 18662 37080
rect 18693 37077 18705 37080
rect 18739 37077 18751 37111
rect 19168 37108 19196 37148
rect 19429 37145 19441 37179
rect 19475 37145 19487 37179
rect 19429 37139 19487 37145
rect 19444 37108 19472 37139
rect 21174 37136 21180 37188
rect 21232 37185 21238 37188
rect 21232 37176 21244 37185
rect 21232 37148 21277 37176
rect 21232 37139 21244 37148
rect 21232 37136 21238 37139
rect 20073 37111 20131 37117
rect 20073 37108 20085 37111
rect 19168 37080 20085 37108
rect 18693 37071 18751 37077
rect 20073 37077 20085 37080
rect 20119 37077 20131 37111
rect 22738 37108 22744 37120
rect 22699 37080 22744 37108
rect 20073 37071 20131 37077
rect 22738 37068 22744 37080
rect 22796 37068 22802 37120
rect 23216 37108 23244 37207
rect 23382 37204 23388 37216
rect 23440 37204 23446 37256
rect 23492 37253 23520 37420
rect 24670 37408 24676 37420
rect 24728 37408 24734 37460
rect 32306 37448 32312 37460
rect 32267 37420 32312 37448
rect 32306 37408 32312 37420
rect 32364 37408 32370 37460
rect 23477 37247 23535 37253
rect 23477 37213 23489 37247
rect 23523 37213 23535 37247
rect 23477 37207 23535 37213
rect 23566 37204 23572 37256
rect 23624 37244 23630 37256
rect 24397 37247 24455 37253
rect 23624 37216 23669 37244
rect 23624 37204 23630 37216
rect 24397 37213 24409 37247
rect 24443 37244 24455 37247
rect 25958 37244 25964 37256
rect 24443 37216 25964 37244
rect 24443 37213 24455 37216
rect 24397 37207 24455 37213
rect 25958 37204 25964 37216
rect 26016 37244 26022 37256
rect 27617 37247 27675 37253
rect 27617 37244 27629 37247
rect 26016 37216 27629 37244
rect 26016 37204 26022 37216
rect 27617 37213 27629 37216
rect 27663 37213 27675 37247
rect 27617 37207 27675 37213
rect 27890 37185 27896 37188
rect 23845 37179 23903 37185
rect 23845 37145 23857 37179
rect 23891 37176 23903 37179
rect 24642 37179 24700 37185
rect 24642 37176 24654 37179
rect 23891 37148 24654 37176
rect 23891 37145 23903 37148
rect 23845 37139 23903 37145
rect 24642 37145 24654 37148
rect 24688 37145 24700 37179
rect 24642 37139 24700 37145
rect 27884 37139 27896 37185
rect 27948 37176 27954 37188
rect 27948 37148 27984 37176
rect 27890 37136 27896 37139
rect 27948 37136 27954 37148
rect 24026 37108 24032 37120
rect 23216 37080 24032 37108
rect 24026 37068 24032 37080
rect 24084 37068 24090 37120
rect 25682 37068 25688 37120
rect 25740 37108 25746 37120
rect 25777 37111 25835 37117
rect 25777 37108 25789 37111
rect 25740 37080 25789 37108
rect 25740 37068 25746 37080
rect 25777 37077 25789 37080
rect 25823 37077 25835 37111
rect 25777 37071 25835 37077
rect 28626 37068 28632 37120
rect 28684 37108 28690 37120
rect 28997 37111 29055 37117
rect 28997 37108 29009 37111
rect 28684 37080 29009 37108
rect 28684 37068 28690 37080
rect 28997 37077 29009 37080
rect 29043 37077 29055 37111
rect 28997 37071 29055 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 2866 36904 2872 36916
rect 2827 36876 2872 36904
rect 2866 36864 2872 36876
rect 2924 36864 2930 36916
rect 6365 36907 6423 36913
rect 6365 36873 6377 36907
rect 6411 36873 6423 36907
rect 6365 36867 6423 36873
rect 10321 36907 10379 36913
rect 10321 36873 10333 36907
rect 10367 36904 10379 36907
rect 10410 36904 10416 36916
rect 10367 36876 10416 36904
rect 10367 36873 10379 36876
rect 10321 36867 10379 36873
rect 3237 36839 3295 36845
rect 3237 36805 3249 36839
rect 3283 36836 3295 36839
rect 5994 36836 6000 36848
rect 3283 36808 6000 36836
rect 3283 36805 3295 36808
rect 3237 36799 3295 36805
rect 5994 36796 6000 36808
rect 6052 36836 6058 36848
rect 6380 36836 6408 36867
rect 10410 36864 10416 36876
rect 10468 36904 10474 36916
rect 10468 36876 11652 36904
rect 10468 36864 10474 36876
rect 10502 36836 10508 36848
rect 6052 36808 6408 36836
rect 8956 36808 10508 36836
rect 6052 36796 6058 36808
rect 3050 36768 3056 36780
rect 3011 36740 3056 36768
rect 3050 36728 3056 36740
rect 3108 36728 3114 36780
rect 8956 36777 8984 36808
rect 10502 36796 10508 36808
rect 10560 36796 10566 36848
rect 6549 36771 6607 36777
rect 6549 36737 6561 36771
rect 6595 36737 6607 36771
rect 6549 36731 6607 36737
rect 8941 36771 8999 36777
rect 8941 36737 8953 36771
rect 8987 36737 8999 36771
rect 8941 36731 8999 36737
rect 9208 36771 9266 36777
rect 9208 36737 9220 36771
rect 9254 36768 9266 36771
rect 10134 36768 10140 36780
rect 9254 36740 10140 36768
rect 9254 36737 9266 36740
rect 9208 36731 9266 36737
rect 6564 36564 6592 36731
rect 10134 36728 10140 36740
rect 10192 36728 10198 36780
rect 11624 36777 11652 36876
rect 11698 36864 11704 36916
rect 11756 36904 11762 36916
rect 12161 36907 12219 36913
rect 11756 36876 11928 36904
rect 11756 36864 11762 36876
rect 11900 36845 11928 36876
rect 12161 36873 12173 36907
rect 12207 36904 12219 36907
rect 18046 36904 18052 36916
rect 12207 36876 18052 36904
rect 12207 36873 12219 36876
rect 12161 36867 12219 36873
rect 18046 36864 18052 36876
rect 18104 36864 18110 36916
rect 24486 36904 24492 36916
rect 23216 36876 24492 36904
rect 11885 36839 11943 36845
rect 11885 36805 11897 36839
rect 11931 36805 11943 36839
rect 11885 36799 11943 36805
rect 12250 36796 12256 36848
rect 12308 36836 12314 36848
rect 12434 36836 12440 36848
rect 12308 36808 12440 36836
rect 12308 36796 12314 36808
rect 12434 36796 12440 36808
rect 12492 36836 12498 36848
rect 12710 36836 12716 36848
rect 12492 36808 12716 36836
rect 12492 36796 12498 36808
rect 12710 36796 12716 36808
rect 12768 36796 12774 36848
rect 13357 36839 13415 36845
rect 13357 36805 13369 36839
rect 13403 36836 13415 36839
rect 13446 36836 13452 36848
rect 13403 36808 13452 36836
rect 13403 36805 13415 36808
rect 13357 36799 13415 36805
rect 13446 36796 13452 36808
rect 13504 36796 13510 36848
rect 14645 36839 14703 36845
rect 14645 36805 14657 36839
rect 14691 36836 14703 36839
rect 15838 36836 15844 36848
rect 14691 36808 15844 36836
rect 14691 36805 14703 36808
rect 14645 36799 14703 36805
rect 15838 36796 15844 36808
rect 15896 36796 15902 36848
rect 23216 36845 23244 36876
rect 24486 36864 24492 36876
rect 24544 36864 24550 36916
rect 24670 36904 24676 36916
rect 24657 36864 24676 36904
rect 24728 36864 24734 36916
rect 25041 36907 25099 36913
rect 25041 36873 25053 36907
rect 25087 36904 25099 36907
rect 25130 36904 25136 36916
rect 25087 36876 25136 36904
rect 25087 36873 25099 36876
rect 25041 36867 25099 36873
rect 25130 36864 25136 36876
rect 25188 36864 25194 36916
rect 27246 36904 27252 36916
rect 27207 36876 27252 36904
rect 27246 36864 27252 36876
rect 27304 36864 27310 36916
rect 27706 36904 27712 36916
rect 27667 36876 27712 36904
rect 27706 36864 27712 36876
rect 27764 36864 27770 36916
rect 17773 36839 17831 36845
rect 17773 36805 17785 36839
rect 17819 36836 17831 36839
rect 19898 36839 19956 36845
rect 19898 36836 19910 36839
rect 17819 36808 19910 36836
rect 17819 36805 17831 36808
rect 17773 36799 17831 36805
rect 19898 36805 19910 36808
rect 19944 36805 19956 36839
rect 19898 36799 19956 36805
rect 23201 36839 23259 36845
rect 23201 36805 23213 36839
rect 23247 36805 23259 36839
rect 24657 36836 24685 36864
rect 24657 36808 24716 36836
rect 23201 36799 23259 36805
rect 11609 36771 11667 36777
rect 11609 36737 11621 36771
rect 11655 36737 11667 36771
rect 11609 36731 11667 36737
rect 11793 36771 11851 36777
rect 11793 36737 11805 36771
rect 11839 36737 11851 36771
rect 11793 36731 11851 36737
rect 11977 36771 12035 36777
rect 11977 36737 11989 36771
rect 12023 36768 12035 36771
rect 12802 36768 12808 36780
rect 12023 36740 12808 36768
rect 12023 36737 12035 36740
rect 11977 36731 12035 36737
rect 11808 36700 11836 36731
rect 12802 36728 12808 36740
rect 12860 36728 12866 36780
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36768 13599 36771
rect 14826 36768 14832 36780
rect 13587 36740 14832 36768
rect 13587 36737 13599 36740
rect 13541 36731 13599 36737
rect 14826 36728 14832 36740
rect 14884 36768 14890 36780
rect 16942 36768 16948 36780
rect 14884 36740 16948 36768
rect 14884 36728 14890 36740
rect 16942 36728 16948 36740
rect 17000 36728 17006 36780
rect 17126 36768 17132 36780
rect 17087 36740 17132 36768
rect 17126 36728 17132 36740
rect 17184 36728 17190 36780
rect 17310 36768 17316 36780
rect 17271 36740 17316 36768
rect 17310 36728 17316 36740
rect 17368 36728 17374 36780
rect 17405 36771 17463 36777
rect 17405 36737 17417 36771
rect 17451 36737 17463 36771
rect 17405 36731 17463 36737
rect 17497 36771 17555 36777
rect 17497 36737 17509 36771
rect 17543 36737 17555 36771
rect 17497 36731 17555 36737
rect 12618 36700 12624 36712
rect 11808 36672 12624 36700
rect 12618 36660 12624 36672
rect 12676 36660 12682 36712
rect 16666 36660 16672 36712
rect 16724 36700 16730 36712
rect 17420 36700 17448 36731
rect 16724 36672 17448 36700
rect 16724 36660 16730 36672
rect 13078 36592 13084 36644
rect 13136 36632 13142 36644
rect 17512 36632 17540 36731
rect 22738 36728 22744 36780
rect 22796 36768 22802 36780
rect 23109 36771 23167 36777
rect 23109 36768 23121 36771
rect 22796 36740 23121 36768
rect 22796 36728 22802 36740
rect 23109 36737 23121 36740
rect 23155 36737 23167 36771
rect 23290 36768 23296 36780
rect 23251 36740 23296 36768
rect 23109 36731 23167 36737
rect 20165 36703 20223 36709
rect 20165 36669 20177 36703
rect 20211 36700 20223 36703
rect 20714 36700 20720 36712
rect 20211 36672 20720 36700
rect 20211 36669 20223 36672
rect 20165 36663 20223 36669
rect 20714 36660 20720 36672
rect 20772 36660 20778 36712
rect 23124 36700 23152 36731
rect 23290 36728 23296 36740
rect 23348 36728 23354 36780
rect 23477 36771 23535 36777
rect 23477 36737 23489 36771
rect 23523 36768 23535 36771
rect 23658 36768 23664 36780
rect 23523 36740 23664 36768
rect 23523 36737 23535 36740
rect 23477 36731 23535 36737
rect 23658 36728 23664 36740
rect 23716 36728 23722 36780
rect 24026 36728 24032 36780
rect 24084 36768 24090 36780
rect 24688 36777 24716 36808
rect 24397 36771 24455 36777
rect 24397 36768 24409 36771
rect 24084 36740 24409 36768
rect 24084 36728 24090 36740
rect 24397 36737 24409 36740
rect 24443 36737 24455 36771
rect 24397 36731 24455 36737
rect 24581 36771 24639 36777
rect 24581 36737 24593 36771
rect 24627 36737 24639 36771
rect 24581 36731 24639 36737
rect 24676 36771 24734 36777
rect 24676 36737 24688 36771
rect 24722 36737 24734 36771
rect 24676 36731 24734 36737
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36768 24823 36771
rect 24854 36768 24860 36780
rect 24811 36740 24860 36768
rect 24811 36737 24823 36740
rect 24765 36731 24823 36737
rect 23382 36700 23388 36712
rect 23124 36672 23388 36700
rect 23382 36660 23388 36672
rect 23440 36660 23446 36712
rect 24118 36660 24124 36712
rect 24176 36700 24182 36712
rect 24596 36700 24624 36731
rect 24854 36728 24860 36740
rect 24912 36728 24918 36780
rect 25498 36768 25504 36780
rect 25459 36740 25504 36768
rect 25498 36728 25504 36740
rect 25556 36728 25562 36780
rect 25682 36768 25688 36780
rect 25643 36740 25688 36768
rect 25682 36728 25688 36740
rect 25740 36728 25746 36780
rect 27264 36768 27292 36864
rect 28071 36777 28077 36780
rect 27939 36771 27997 36777
rect 27939 36768 27951 36771
rect 27264 36740 27951 36768
rect 27939 36737 27951 36740
rect 27985 36737 27997 36771
rect 27939 36731 27997 36737
rect 28058 36771 28077 36777
rect 28058 36737 28070 36771
rect 28058 36731 28077 36737
rect 28071 36728 28077 36731
rect 28129 36728 28135 36780
rect 28174 36771 28232 36777
rect 28174 36737 28186 36771
rect 28220 36737 28232 36771
rect 28174 36731 28232 36737
rect 28353 36771 28411 36777
rect 28353 36737 28365 36771
rect 28399 36768 28411 36771
rect 28813 36771 28871 36777
rect 28813 36768 28825 36771
rect 28399 36740 28825 36768
rect 28399 36737 28411 36740
rect 28353 36731 28411 36737
rect 28813 36737 28825 36740
rect 28859 36737 28871 36771
rect 33410 36768 33416 36780
rect 33371 36740 33416 36768
rect 28813 36731 28871 36737
rect 24176 36672 24624 36700
rect 24176 36660 24182 36672
rect 28189 36644 28217 36731
rect 28258 36660 28264 36712
rect 28316 36700 28322 36712
rect 28368 36700 28396 36731
rect 33410 36728 33416 36740
rect 33468 36728 33474 36780
rect 33597 36771 33655 36777
rect 33597 36737 33609 36771
rect 33643 36768 33655 36771
rect 34514 36768 34520 36780
rect 33643 36740 34520 36768
rect 33643 36737 33655 36740
rect 33597 36731 33655 36737
rect 34514 36728 34520 36740
rect 34572 36728 34578 36780
rect 28316 36672 28396 36700
rect 28316 36660 28322 36672
rect 18233 36635 18291 36641
rect 18233 36632 18245 36635
rect 13136 36604 18245 36632
rect 13136 36592 13142 36604
rect 18233 36601 18245 36604
rect 18279 36632 18291 36635
rect 18279 36604 19288 36632
rect 18279 36601 18291 36604
rect 18233 36595 18291 36601
rect 12250 36564 12256 36576
rect 6564 36536 12256 36564
rect 12250 36524 12256 36536
rect 12308 36524 12314 36576
rect 12894 36524 12900 36576
rect 12952 36564 12958 36576
rect 13173 36567 13231 36573
rect 13173 36564 13185 36567
rect 12952 36536 13185 36564
rect 12952 36524 12958 36536
rect 13173 36533 13185 36536
rect 13219 36533 13231 36567
rect 13173 36527 13231 36533
rect 14461 36567 14519 36573
rect 14461 36533 14473 36567
rect 14507 36564 14519 36567
rect 14550 36564 14556 36576
rect 14507 36536 14556 36564
rect 14507 36533 14519 36536
rect 14461 36527 14519 36533
rect 14550 36524 14556 36536
rect 14608 36524 14614 36576
rect 18690 36524 18696 36576
rect 18748 36564 18754 36576
rect 18785 36567 18843 36573
rect 18785 36564 18797 36567
rect 18748 36536 18797 36564
rect 18748 36524 18754 36536
rect 18785 36533 18797 36536
rect 18831 36533 18843 36567
rect 19260 36564 19288 36604
rect 28166 36592 28172 36644
rect 28224 36592 28230 36644
rect 31754 36592 31760 36644
rect 31812 36632 31818 36644
rect 32030 36632 32036 36644
rect 31812 36604 32036 36632
rect 31812 36592 31818 36604
rect 32030 36592 32036 36604
rect 32088 36632 32094 36644
rect 34241 36635 34299 36641
rect 34241 36632 34253 36635
rect 32088 36604 34253 36632
rect 32088 36592 32094 36604
rect 34241 36601 34253 36604
rect 34287 36632 34299 36635
rect 36630 36632 36636 36644
rect 34287 36604 36636 36632
rect 34287 36601 34299 36604
rect 34241 36595 34299 36601
rect 36630 36592 36636 36604
rect 36688 36592 36694 36644
rect 20806 36564 20812 36576
rect 19260 36536 20812 36564
rect 18785 36527 18843 36533
rect 20806 36524 20812 36536
rect 20864 36524 20870 36576
rect 22462 36564 22468 36576
rect 22423 36536 22468 36564
rect 22462 36524 22468 36536
rect 22520 36524 22526 36576
rect 22554 36524 22560 36576
rect 22612 36564 22618 36576
rect 22925 36567 22983 36573
rect 22925 36564 22937 36567
rect 22612 36536 22937 36564
rect 22612 36524 22618 36536
rect 22925 36533 22937 36536
rect 22971 36533 22983 36567
rect 22925 36527 22983 36533
rect 23474 36524 23480 36576
rect 23532 36564 23538 36576
rect 25869 36567 25927 36573
rect 25869 36564 25881 36567
rect 23532 36536 25881 36564
rect 23532 36524 23538 36536
rect 25869 36533 25881 36536
rect 25915 36533 25927 36567
rect 33778 36564 33784 36576
rect 33739 36536 33784 36564
rect 25869 36527 25927 36533
rect 33778 36524 33784 36536
rect 33836 36524 33842 36576
rect 34885 36567 34943 36573
rect 34885 36533 34897 36567
rect 34931 36564 34943 36567
rect 35342 36564 35348 36576
rect 34931 36536 35348 36564
rect 34931 36533 34943 36536
rect 34885 36527 34943 36533
rect 35342 36524 35348 36536
rect 35400 36524 35406 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 10134 36360 10140 36372
rect 10095 36332 10140 36360
rect 10134 36320 10140 36332
rect 10192 36320 10198 36372
rect 11333 36363 11391 36369
rect 11333 36329 11345 36363
rect 11379 36360 11391 36363
rect 13078 36360 13084 36372
rect 11379 36332 13084 36360
rect 11379 36329 11391 36332
rect 11333 36323 11391 36329
rect 7469 36295 7527 36301
rect 7469 36261 7481 36295
rect 7515 36261 7527 36295
rect 11348 36292 11376 36323
rect 13078 36320 13084 36332
rect 13136 36320 13142 36372
rect 13173 36363 13231 36369
rect 13173 36329 13185 36363
rect 13219 36360 13231 36363
rect 13446 36360 13452 36372
rect 13219 36332 13452 36360
rect 13219 36329 13231 36332
rect 13173 36323 13231 36329
rect 13446 36320 13452 36332
rect 13504 36320 13510 36372
rect 14090 36360 14096 36372
rect 14051 36332 14096 36360
rect 14090 36320 14096 36332
rect 14148 36320 14154 36372
rect 16669 36363 16727 36369
rect 16669 36329 16681 36363
rect 16715 36360 16727 36363
rect 16758 36360 16764 36372
rect 16715 36332 16764 36360
rect 16715 36329 16727 36332
rect 16669 36323 16727 36329
rect 16758 36320 16764 36332
rect 16816 36320 16822 36372
rect 17310 36360 17316 36372
rect 17271 36332 17316 36360
rect 17310 36320 17316 36332
rect 17368 36320 17374 36372
rect 20806 36360 20812 36372
rect 20767 36332 20812 36360
rect 20806 36320 20812 36332
rect 20864 36320 20870 36372
rect 24118 36320 24124 36372
rect 24176 36360 24182 36372
rect 24397 36363 24455 36369
rect 24397 36360 24409 36363
rect 24176 36332 24409 36360
rect 24176 36320 24182 36332
rect 24397 36329 24409 36332
rect 24443 36329 24455 36363
rect 24397 36323 24455 36329
rect 27617 36363 27675 36369
rect 27617 36329 27629 36363
rect 27663 36360 27675 36363
rect 27890 36360 27896 36372
rect 27663 36332 27896 36360
rect 27663 36329 27675 36332
rect 27617 36323 27675 36329
rect 27890 36320 27896 36332
rect 27948 36320 27954 36372
rect 33318 36360 33324 36372
rect 33279 36332 33324 36360
rect 33318 36320 33324 36332
rect 33376 36320 33382 36372
rect 36630 36360 36636 36372
rect 36591 36332 36636 36360
rect 36630 36320 36636 36332
rect 36688 36320 36694 36372
rect 7469 36255 7527 36261
rect 10428 36264 11376 36292
rect 7484 36224 7512 36255
rect 8294 36224 8300 36236
rect 7484 36196 8300 36224
rect 8294 36184 8300 36196
rect 8352 36184 8358 36236
rect 6086 36156 6092 36168
rect 6047 36128 6092 36156
rect 6086 36116 6092 36128
rect 6144 36116 6150 36168
rect 8113 36159 8171 36165
rect 8113 36125 8125 36159
rect 8159 36156 8171 36159
rect 8312 36156 8340 36184
rect 10428 36165 10456 36264
rect 28074 36252 28080 36304
rect 28132 36252 28138 36304
rect 14642 36224 14648 36236
rect 14476 36196 14648 36224
rect 8159 36128 8340 36156
rect 10413 36159 10471 36165
rect 8159 36125 8171 36128
rect 8113 36119 8171 36125
rect 10413 36125 10425 36159
rect 10459 36125 10471 36159
rect 10413 36119 10471 36125
rect 10505 36159 10563 36165
rect 10505 36125 10517 36159
rect 10551 36125 10563 36159
rect 10505 36119 10563 36125
rect 6356 36091 6414 36097
rect 6356 36057 6368 36091
rect 6402 36088 6414 36091
rect 6914 36088 6920 36100
rect 6402 36060 6920 36088
rect 6402 36057 6414 36060
rect 6356 36051 6414 36057
rect 6914 36048 6920 36060
rect 6972 36048 6978 36100
rect 7374 36048 7380 36100
rect 7432 36088 7438 36100
rect 7929 36091 7987 36097
rect 7929 36088 7941 36091
rect 7432 36060 7941 36088
rect 7432 36048 7438 36060
rect 7929 36057 7941 36060
rect 7975 36057 7987 36091
rect 8294 36088 8300 36100
rect 8255 36060 8300 36088
rect 7929 36051 7987 36057
rect 8294 36048 8300 36060
rect 8352 36048 8358 36100
rect 9950 36048 9956 36100
rect 10008 36088 10014 36100
rect 10520 36088 10548 36119
rect 10594 36116 10600 36168
rect 10652 36156 10658 36168
rect 10781 36159 10839 36165
rect 10652 36128 10697 36156
rect 10652 36116 10658 36128
rect 10781 36125 10793 36159
rect 10827 36156 10839 36159
rect 10870 36156 10876 36168
rect 10827 36128 10876 36156
rect 10827 36125 10839 36128
rect 10781 36119 10839 36125
rect 10870 36116 10876 36128
rect 10928 36116 10934 36168
rect 11793 36159 11851 36165
rect 11793 36125 11805 36159
rect 11839 36125 11851 36159
rect 14366 36156 14372 36168
rect 14327 36128 14372 36156
rect 11793 36119 11851 36125
rect 10008 36060 10548 36088
rect 10008 36048 10014 36060
rect 10428 36032 10456 36060
rect 4982 35980 4988 36032
rect 5040 36020 5046 36032
rect 5534 36020 5540 36032
rect 5040 35992 5540 36020
rect 5040 35980 5046 35992
rect 5534 35980 5540 35992
rect 5592 35980 5598 36032
rect 10410 35980 10416 36032
rect 10468 35980 10474 36032
rect 10502 35980 10508 36032
rect 10560 36020 10566 36032
rect 11808 36020 11836 36119
rect 14366 36116 14372 36128
rect 14424 36116 14430 36168
rect 14476 36165 14504 36196
rect 14642 36184 14648 36196
rect 14700 36224 14706 36236
rect 16666 36224 16672 36236
rect 14700 36196 16672 36224
rect 14700 36184 14706 36196
rect 14461 36159 14519 36165
rect 14461 36125 14473 36159
rect 14507 36125 14519 36159
rect 14461 36119 14519 36125
rect 14550 36116 14556 36168
rect 14608 36156 14614 36168
rect 14737 36159 14795 36165
rect 14608 36128 14653 36156
rect 14608 36116 14614 36128
rect 14737 36125 14749 36159
rect 14783 36156 14795 36159
rect 16025 36159 16083 36165
rect 16025 36156 16037 36159
rect 14783 36128 16037 36156
rect 14783 36125 14795 36128
rect 14737 36119 14795 36125
rect 16025 36125 16037 36128
rect 16071 36125 16083 36159
rect 16206 36156 16212 36168
rect 16167 36128 16212 36156
rect 16025 36119 16083 36125
rect 12060 36091 12118 36097
rect 12060 36057 12072 36091
rect 12106 36088 12118 36091
rect 12434 36088 12440 36100
rect 12106 36060 12440 36088
rect 12106 36057 12118 36060
rect 12060 36051 12118 36057
rect 12434 36048 12440 36060
rect 12492 36048 12498 36100
rect 13906 36048 13912 36100
rect 13964 36088 13970 36100
rect 14752 36088 14780 36119
rect 13964 36060 14780 36088
rect 16040 36088 16068 36119
rect 16206 36116 16212 36128
rect 16264 36116 16270 36168
rect 16316 36165 16344 36196
rect 16666 36184 16672 36196
rect 16724 36184 16730 36236
rect 25682 36224 25688 36236
rect 23400 36196 25688 36224
rect 16301 36159 16359 36165
rect 16301 36125 16313 36159
rect 16347 36125 16359 36159
rect 16301 36119 16359 36125
rect 16390 36116 16396 36168
rect 16448 36156 16454 36168
rect 16448 36128 16493 36156
rect 16448 36116 16454 36128
rect 17034 36116 17040 36168
rect 17092 36156 17098 36168
rect 17497 36159 17555 36165
rect 17092 36128 17264 36156
rect 17092 36116 17098 36128
rect 17126 36088 17132 36100
rect 16040 36060 17132 36088
rect 13964 36048 13970 36060
rect 17126 36048 17132 36060
rect 17184 36048 17190 36100
rect 17236 36088 17264 36128
rect 17497 36125 17509 36159
rect 17543 36156 17555 36159
rect 18690 36156 18696 36168
rect 17543 36128 18696 36156
rect 17543 36125 17555 36128
rect 17497 36119 17555 36125
rect 18690 36116 18696 36128
rect 18748 36116 18754 36168
rect 20806 36116 20812 36168
rect 20864 36156 20870 36168
rect 21637 36159 21695 36165
rect 21637 36156 21649 36159
rect 20864 36128 21649 36156
rect 20864 36116 20870 36128
rect 21637 36125 21649 36128
rect 21683 36125 21695 36159
rect 21637 36119 21695 36125
rect 21729 36159 21787 36165
rect 21729 36125 21741 36159
rect 21775 36125 21787 36159
rect 21729 36119 21787 36125
rect 17678 36088 17684 36100
rect 17236 36060 17684 36088
rect 17678 36048 17684 36060
rect 17736 36048 17742 36100
rect 21744 36088 21772 36119
rect 21818 36116 21824 36168
rect 21876 36156 21882 36168
rect 22005 36159 22063 36165
rect 21876 36128 21921 36156
rect 21876 36116 21882 36128
rect 22005 36125 22017 36159
rect 22051 36156 22063 36159
rect 22278 36156 22284 36168
rect 22051 36128 22284 36156
rect 22051 36125 22063 36128
rect 22005 36119 22063 36125
rect 22278 36116 22284 36128
rect 22336 36116 22342 36168
rect 22646 36116 22652 36168
rect 22704 36156 22710 36168
rect 23400 36165 23428 36196
rect 25682 36184 25688 36196
rect 25740 36184 25746 36236
rect 28092 36224 28120 36252
rect 28442 36224 28448 36236
rect 28000 36196 28448 36224
rect 23109 36159 23167 36165
rect 23109 36156 23121 36159
rect 22704 36128 23121 36156
rect 22704 36116 22710 36128
rect 23109 36125 23121 36128
rect 23155 36125 23167 36159
rect 23109 36119 23167 36125
rect 23385 36159 23443 36165
rect 23385 36125 23397 36159
rect 23431 36125 23443 36159
rect 23385 36119 23443 36125
rect 23474 36116 23480 36168
rect 23532 36156 23538 36168
rect 23532 36128 23577 36156
rect 23532 36116 23538 36128
rect 24486 36116 24492 36168
rect 24544 36156 24550 36168
rect 24581 36159 24639 36165
rect 24581 36156 24593 36159
rect 24544 36128 24593 36156
rect 24544 36116 24550 36128
rect 24581 36125 24593 36128
rect 24627 36125 24639 36159
rect 24581 36119 24639 36125
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36156 24823 36159
rect 24854 36156 24860 36168
rect 24811 36128 24860 36156
rect 24811 36125 24823 36128
rect 24765 36119 24823 36125
rect 24854 36116 24860 36128
rect 24912 36156 24918 36168
rect 25498 36156 25504 36168
rect 24912 36128 25504 36156
rect 24912 36116 24918 36128
rect 25498 36116 25504 36128
rect 25556 36116 25562 36168
rect 27798 36116 27804 36168
rect 27856 36165 27862 36168
rect 28000 36165 28028 36196
rect 28442 36184 28448 36196
rect 28500 36184 28506 36236
rect 33502 36184 33508 36236
rect 33560 36224 33566 36236
rect 33560 36196 35020 36224
rect 33560 36184 33566 36196
rect 27856 36159 27905 36165
rect 27856 36125 27859 36159
rect 27893 36125 27905 36159
rect 27856 36119 27905 36125
rect 27985 36159 28043 36165
rect 27985 36125 27997 36159
rect 28031 36125 28043 36159
rect 27985 36119 28043 36125
rect 28077 36159 28135 36165
rect 28077 36125 28089 36159
rect 28123 36125 28135 36159
rect 28258 36156 28264 36168
rect 28219 36128 28264 36156
rect 28077 36119 28135 36125
rect 27856 36116 27862 36119
rect 22186 36088 22192 36100
rect 21744 36060 22192 36088
rect 22186 36048 22192 36060
rect 22244 36048 22250 36100
rect 22462 36048 22468 36100
rect 22520 36088 22526 36100
rect 23290 36088 23296 36100
rect 22520 36060 23296 36088
rect 22520 36048 22526 36060
rect 22664 36032 22692 36060
rect 23290 36048 23296 36060
rect 23348 36048 23354 36100
rect 26605 36091 26663 36097
rect 26605 36057 26617 36091
rect 26651 36088 26663 36091
rect 27614 36088 27620 36100
rect 26651 36060 27620 36088
rect 26651 36057 26663 36060
rect 26605 36051 26663 36057
rect 27614 36048 27620 36060
rect 27672 36048 27678 36100
rect 10560 35992 11836 36020
rect 10560 35980 10566 35992
rect 14366 35980 14372 36032
rect 14424 36020 14430 36032
rect 15289 36023 15347 36029
rect 15289 36020 15301 36023
rect 14424 35992 15301 36020
rect 14424 35980 14430 35992
rect 15289 35989 15301 35992
rect 15335 36020 15347 36023
rect 15562 36020 15568 36032
rect 15335 35992 15568 36020
rect 15335 35989 15347 35992
rect 15289 35983 15347 35989
rect 15562 35980 15568 35992
rect 15620 35980 15626 36032
rect 21361 36023 21419 36029
rect 21361 35989 21373 36023
rect 21407 36020 21419 36023
rect 22370 36020 22376 36032
rect 21407 35992 22376 36020
rect 21407 35989 21419 35992
rect 21361 35983 21419 35989
rect 22370 35980 22376 35992
rect 22428 35980 22434 36032
rect 22646 36020 22652 36032
rect 22607 35992 22652 36020
rect 22646 35980 22652 35992
rect 22704 35980 22710 36032
rect 23658 36020 23664 36032
rect 23619 35992 23664 36020
rect 23658 35980 23664 35992
rect 23716 35980 23722 36032
rect 24486 35980 24492 36032
rect 24544 36020 24550 36032
rect 24762 36020 24768 36032
rect 24544 35992 24768 36020
rect 24544 35980 24550 35992
rect 24762 35980 24768 35992
rect 24820 35980 24826 36032
rect 27157 36023 27215 36029
rect 27157 35989 27169 36023
rect 27203 36020 27215 36023
rect 27798 36020 27804 36032
rect 27203 35992 27804 36020
rect 27203 35989 27215 35992
rect 27157 35983 27215 35989
rect 27798 35980 27804 35992
rect 27856 35980 27862 36032
rect 28092 36020 28120 36119
rect 28258 36116 28264 36128
rect 28316 36116 28322 36168
rect 33594 36116 33600 36168
rect 33652 36156 33658 36168
rect 34992 36165 35020 36196
rect 34701 36159 34759 36165
rect 34701 36156 34713 36159
rect 33652 36128 34713 36156
rect 33652 36116 33658 36128
rect 34701 36125 34713 36128
rect 34747 36125 34759 36159
rect 34701 36119 34759 36125
rect 34885 36159 34943 36165
rect 34885 36125 34897 36159
rect 34931 36125 34943 36159
rect 34885 36119 34943 36125
rect 34977 36159 35035 36165
rect 34977 36125 34989 36159
rect 35023 36125 35035 36159
rect 34977 36119 35035 36125
rect 35069 36159 35127 36165
rect 35069 36125 35081 36159
rect 35115 36156 35127 36159
rect 35342 36156 35348 36168
rect 35115 36128 35348 36156
rect 35115 36125 35127 36128
rect 35069 36119 35127 36125
rect 30098 36088 30104 36100
rect 30059 36060 30104 36088
rect 30098 36048 30104 36060
rect 30156 36048 30162 36100
rect 30285 36091 30343 36097
rect 30285 36057 30297 36091
rect 30331 36088 30343 36091
rect 30926 36088 30932 36100
rect 30331 36060 30932 36088
rect 30331 36057 30343 36060
rect 30285 36051 30343 36057
rect 30926 36048 30932 36060
rect 30984 36048 30990 36100
rect 31021 36091 31079 36097
rect 31021 36057 31033 36091
rect 31067 36057 31079 36091
rect 31021 36051 31079 36057
rect 28534 36020 28540 36032
rect 28092 35992 28540 36020
rect 28534 35980 28540 35992
rect 28592 35980 28598 36032
rect 30834 36020 30840 36032
rect 30795 35992 30840 36020
rect 30834 35980 30840 35992
rect 30892 35980 30898 36032
rect 31036 36020 31064 36051
rect 31110 36048 31116 36100
rect 31168 36088 31174 36100
rect 31205 36091 31263 36097
rect 31205 36088 31217 36091
rect 31168 36060 31217 36088
rect 31168 36048 31174 36060
rect 31205 36057 31217 36060
rect 31251 36057 31263 36091
rect 32030 36088 32036 36100
rect 31991 36060 32036 36088
rect 31205 36051 31263 36057
rect 32030 36048 32036 36060
rect 32088 36048 32094 36100
rect 33134 36048 33140 36100
rect 33192 36088 33198 36100
rect 34900 36088 34928 36119
rect 35342 36116 35348 36128
rect 35400 36116 35406 36168
rect 36648 36156 36676 36320
rect 38933 36159 38991 36165
rect 38933 36156 38945 36159
rect 36648 36128 38945 36156
rect 38933 36125 38945 36128
rect 38979 36125 38991 36159
rect 58158 36156 58164 36168
rect 58119 36128 58164 36156
rect 38933 36119 38991 36125
rect 58158 36116 58164 36128
rect 58216 36116 58222 36168
rect 33192 36060 34928 36088
rect 33192 36048 33198 36060
rect 36078 36048 36084 36100
rect 36136 36088 36142 36100
rect 37277 36091 37335 36097
rect 37277 36088 37289 36091
rect 36136 36060 37289 36088
rect 36136 36048 36142 36060
rect 37277 36057 37289 36060
rect 37323 36088 37335 36091
rect 38562 36088 38568 36100
rect 37323 36060 38568 36088
rect 37323 36057 37335 36060
rect 37277 36051 37335 36057
rect 38562 36048 38568 36060
rect 38620 36048 38626 36100
rect 32398 36020 32404 36032
rect 31036 35992 32404 36020
rect 32398 35980 32404 35992
rect 32456 35980 32462 36032
rect 34606 35980 34612 36032
rect 34664 36020 34670 36032
rect 35345 36023 35403 36029
rect 35345 36020 35357 36023
rect 34664 35992 35357 36020
rect 34664 35980 34670 35992
rect 35345 35989 35357 35992
rect 35391 35989 35403 36023
rect 35345 35983 35403 35989
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 6914 35816 6920 35828
rect 6875 35788 6920 35816
rect 6914 35776 6920 35788
rect 6972 35776 6978 35828
rect 12434 35776 12440 35828
rect 12492 35816 12498 35828
rect 12492 35788 12537 35816
rect 12728 35788 13676 35816
rect 12492 35776 12498 35788
rect 10318 35708 10324 35760
rect 10376 35748 10382 35760
rect 10413 35751 10471 35757
rect 10413 35748 10425 35751
rect 10376 35720 10425 35748
rect 10376 35708 10382 35720
rect 10413 35717 10425 35720
rect 10459 35717 10471 35751
rect 10870 35748 10876 35760
rect 10413 35711 10471 35717
rect 10520 35720 10876 35748
rect 3044 35683 3102 35689
rect 3044 35649 3056 35683
rect 3090 35680 3102 35683
rect 4062 35680 4068 35692
rect 3090 35652 4068 35680
rect 3090 35649 3102 35652
rect 3044 35643 3102 35649
rect 4062 35640 4068 35652
rect 4120 35640 4126 35692
rect 7193 35683 7251 35689
rect 7193 35680 7205 35683
rect 6380 35652 7205 35680
rect 2774 35572 2780 35624
rect 2832 35612 2838 35624
rect 2832 35584 2877 35612
rect 2832 35572 2838 35584
rect 4157 35479 4215 35485
rect 4157 35445 4169 35479
rect 4203 35476 4215 35479
rect 4706 35476 4712 35488
rect 4203 35448 4712 35476
rect 4203 35445 4215 35448
rect 4157 35439 4215 35445
rect 4706 35436 4712 35448
rect 4764 35436 4770 35488
rect 6270 35436 6276 35488
rect 6328 35476 6334 35488
rect 6380 35485 6408 35652
rect 7193 35649 7205 35652
rect 7239 35649 7251 35683
rect 7193 35643 7251 35649
rect 7285 35683 7343 35689
rect 7285 35649 7297 35683
rect 7331 35649 7343 35683
rect 7285 35643 7343 35649
rect 7300 35612 7328 35643
rect 7374 35640 7380 35692
rect 7432 35680 7438 35692
rect 7561 35683 7619 35689
rect 7432 35652 7477 35680
rect 7432 35640 7438 35652
rect 7561 35649 7573 35683
rect 7607 35680 7619 35683
rect 10226 35680 10232 35692
rect 7607 35652 10232 35680
rect 7607 35649 7619 35652
rect 7561 35643 7619 35649
rect 10226 35640 10232 35652
rect 10284 35680 10290 35692
rect 10520 35680 10548 35720
rect 10870 35708 10876 35720
rect 10928 35708 10934 35760
rect 10962 35708 10968 35760
rect 11020 35748 11026 35760
rect 12728 35748 12756 35788
rect 11020 35720 12756 35748
rect 11020 35708 11026 35720
rect 10284 35652 10548 35680
rect 10597 35683 10655 35689
rect 10284 35640 10290 35652
rect 10597 35649 10609 35683
rect 10643 35680 10655 35683
rect 11882 35680 11888 35692
rect 10643 35652 11888 35680
rect 10643 35649 10655 35652
rect 10597 35643 10655 35649
rect 11882 35640 11888 35652
rect 11940 35640 11946 35692
rect 12728 35689 12756 35720
rect 12820 35720 13584 35748
rect 12820 35689 12848 35720
rect 12713 35683 12771 35689
rect 12713 35649 12725 35683
rect 12759 35649 12771 35683
rect 12713 35643 12771 35649
rect 12805 35683 12863 35689
rect 12805 35649 12817 35683
rect 12851 35649 12863 35683
rect 12805 35643 12863 35649
rect 12894 35640 12900 35692
rect 12952 35680 12958 35692
rect 13081 35683 13139 35689
rect 12952 35652 12997 35680
rect 12952 35640 12958 35652
rect 13081 35649 13093 35683
rect 13127 35649 13139 35683
rect 13081 35643 13139 35649
rect 7650 35612 7656 35624
rect 7300 35584 7656 35612
rect 7650 35572 7656 35584
rect 7708 35572 7714 35624
rect 7558 35504 7564 35556
rect 7616 35544 7622 35556
rect 11885 35547 11943 35553
rect 11885 35544 11897 35547
rect 7616 35516 11897 35544
rect 7616 35504 7622 35516
rect 11885 35513 11897 35516
rect 11931 35544 11943 35547
rect 13096 35544 13124 35643
rect 13556 35612 13584 35720
rect 13648 35689 13676 35788
rect 16574 35776 16580 35828
rect 16632 35816 16638 35828
rect 16761 35819 16819 35825
rect 16761 35816 16773 35819
rect 16632 35788 16773 35816
rect 16632 35776 16638 35788
rect 16761 35785 16773 35788
rect 16807 35785 16819 35819
rect 16761 35779 16819 35785
rect 16776 35748 16804 35779
rect 19334 35776 19340 35828
rect 19392 35816 19398 35828
rect 19518 35816 19524 35828
rect 19392 35788 19524 35816
rect 19392 35776 19398 35788
rect 19518 35776 19524 35788
rect 19576 35776 19582 35828
rect 21818 35816 21824 35828
rect 21779 35788 21824 35816
rect 21818 35776 21824 35788
rect 21876 35776 21882 35828
rect 24946 35816 24952 35828
rect 21928 35788 24952 35816
rect 21928 35748 21956 35788
rect 24946 35776 24952 35788
rect 25004 35816 25010 35828
rect 25682 35816 25688 35828
rect 25004 35788 25688 35816
rect 25004 35776 25010 35788
rect 25682 35776 25688 35788
rect 25740 35776 25746 35828
rect 28166 35776 28172 35828
rect 28224 35816 28230 35828
rect 29181 35819 29239 35825
rect 29181 35816 29193 35819
rect 28224 35788 29193 35816
rect 28224 35776 28230 35788
rect 29181 35785 29193 35788
rect 29227 35785 29239 35819
rect 29181 35779 29239 35785
rect 32861 35819 32919 35825
rect 32861 35785 32873 35819
rect 32907 35816 32919 35819
rect 33134 35816 33140 35828
rect 32907 35788 33140 35816
rect 32907 35785 32919 35788
rect 32861 35779 32919 35785
rect 33134 35776 33140 35788
rect 33192 35776 33198 35828
rect 16776 35720 21956 35748
rect 22005 35751 22063 35757
rect 22005 35717 22017 35751
rect 22051 35748 22063 35751
rect 22094 35748 22100 35760
rect 22051 35720 22100 35748
rect 22051 35717 22063 35720
rect 22005 35711 22063 35717
rect 22094 35708 22100 35720
rect 22152 35708 22158 35760
rect 33318 35708 33324 35760
rect 33376 35748 33382 35760
rect 33376 35720 34744 35748
rect 33376 35708 33382 35720
rect 13633 35683 13691 35689
rect 13633 35649 13645 35683
rect 13679 35680 13691 35683
rect 21910 35680 21916 35692
rect 13679 35652 21916 35680
rect 13679 35649 13691 35652
rect 13633 35643 13691 35649
rect 21910 35640 21916 35652
rect 21968 35640 21974 35692
rect 22189 35683 22247 35689
rect 22189 35649 22201 35683
rect 22235 35680 22247 35683
rect 22830 35680 22836 35692
rect 22235 35652 22836 35680
rect 22235 35649 22247 35652
rect 22189 35643 22247 35649
rect 22830 35640 22836 35652
rect 22888 35640 22894 35692
rect 27430 35640 27436 35692
rect 27488 35680 27494 35692
rect 27597 35683 27655 35689
rect 27597 35680 27609 35683
rect 27488 35652 27609 35680
rect 27488 35640 27494 35652
rect 27597 35649 27609 35652
rect 27643 35649 27655 35683
rect 27597 35643 27655 35649
rect 28994 35640 29000 35692
rect 29052 35680 29058 35692
rect 29365 35683 29423 35689
rect 29365 35680 29377 35683
rect 29052 35652 29377 35680
rect 29052 35640 29058 35652
rect 29365 35649 29377 35652
rect 29411 35649 29423 35683
rect 29365 35643 29423 35649
rect 29546 35640 29552 35692
rect 29604 35680 29610 35692
rect 31110 35680 31116 35692
rect 29604 35652 31116 35680
rect 29604 35640 29610 35652
rect 31110 35640 31116 35652
rect 31168 35640 31174 35692
rect 32493 35683 32551 35689
rect 32493 35649 32505 35683
rect 32539 35649 32551 35683
rect 32493 35643 32551 35649
rect 32677 35683 32735 35689
rect 32677 35649 32689 35683
rect 32723 35680 32735 35683
rect 33042 35680 33048 35692
rect 32723 35652 33048 35680
rect 32723 35649 32735 35652
rect 32677 35643 32735 35649
rect 14642 35612 14648 35624
rect 13556 35584 14648 35612
rect 14642 35572 14648 35584
rect 14700 35572 14706 35624
rect 27338 35612 27344 35624
rect 27299 35584 27344 35612
rect 27338 35572 27344 35584
rect 27396 35572 27402 35624
rect 30466 35572 30472 35624
rect 30524 35612 30530 35624
rect 31021 35615 31079 35621
rect 31021 35612 31033 35615
rect 30524 35584 31033 35612
rect 30524 35572 30530 35584
rect 31021 35581 31033 35584
rect 31067 35612 31079 35615
rect 31202 35612 31208 35624
rect 31067 35584 31208 35612
rect 31067 35581 31079 35584
rect 31021 35575 31079 35581
rect 31202 35572 31208 35584
rect 31260 35572 31266 35624
rect 31297 35615 31355 35621
rect 31297 35581 31309 35615
rect 31343 35612 31355 35615
rect 31570 35612 31576 35624
rect 31343 35584 31576 35612
rect 31343 35581 31355 35584
rect 31297 35575 31355 35581
rect 31570 35572 31576 35584
rect 31628 35572 31634 35624
rect 32508 35612 32536 35643
rect 33042 35640 33048 35652
rect 33100 35640 33106 35692
rect 34445 35683 34503 35689
rect 34445 35649 34457 35683
rect 34491 35680 34503 35683
rect 34606 35680 34612 35692
rect 34491 35652 34612 35680
rect 34491 35649 34503 35652
rect 34445 35643 34503 35649
rect 34606 35640 34612 35652
rect 34664 35640 34670 35692
rect 34716 35689 34744 35720
rect 36078 35708 36084 35760
rect 36136 35748 36142 35760
rect 36136 35720 36584 35748
rect 36136 35708 36142 35720
rect 34701 35683 34759 35689
rect 34701 35649 34713 35683
rect 34747 35649 34759 35683
rect 34701 35643 34759 35649
rect 34790 35640 34796 35692
rect 34848 35680 34854 35692
rect 36556 35689 36584 35720
rect 36274 35683 36332 35689
rect 36274 35680 36286 35683
rect 34848 35652 36286 35680
rect 34848 35640 34854 35652
rect 36274 35649 36286 35652
rect 36320 35649 36332 35683
rect 36274 35643 36332 35649
rect 36541 35683 36599 35689
rect 36541 35649 36553 35683
rect 36587 35649 36599 35683
rect 36541 35643 36599 35649
rect 33134 35612 33140 35624
rect 32508 35584 33140 35612
rect 33134 35572 33140 35584
rect 33192 35612 33198 35624
rect 33410 35612 33416 35624
rect 33192 35584 33416 35612
rect 33192 35572 33198 35584
rect 33410 35572 33416 35584
rect 33468 35572 33474 35624
rect 11931 35516 13124 35544
rect 11931 35513 11943 35516
rect 11885 35507 11943 35513
rect 19334 35504 19340 35556
rect 19392 35544 19398 35556
rect 19705 35547 19763 35553
rect 19705 35544 19717 35547
rect 19392 35516 19717 35544
rect 19392 35504 19398 35516
rect 19705 35513 19717 35516
rect 19751 35544 19763 35547
rect 23658 35544 23664 35556
rect 19751 35516 23664 35544
rect 19751 35513 19763 35516
rect 19705 35507 19763 35513
rect 23658 35504 23664 35516
rect 23716 35504 23722 35556
rect 6365 35479 6423 35485
rect 6365 35476 6377 35479
rect 6328 35448 6377 35476
rect 6328 35436 6334 35448
rect 6365 35445 6377 35448
rect 6411 35445 6423 35479
rect 6365 35439 6423 35445
rect 10686 35436 10692 35488
rect 10744 35476 10750 35488
rect 10781 35479 10839 35485
rect 10781 35476 10793 35479
rect 10744 35448 10793 35476
rect 10744 35436 10750 35448
rect 10781 35445 10793 35448
rect 10827 35445 10839 35479
rect 10781 35439 10839 35445
rect 16850 35436 16856 35488
rect 16908 35476 16914 35488
rect 17313 35479 17371 35485
rect 17313 35476 17325 35479
rect 16908 35448 17325 35476
rect 16908 35436 16914 35448
rect 17313 35445 17325 35448
rect 17359 35445 17371 35479
rect 17313 35439 17371 35445
rect 23382 35436 23388 35488
rect 23440 35476 23446 35488
rect 23753 35479 23811 35485
rect 23753 35476 23765 35479
rect 23440 35448 23765 35476
rect 23440 35436 23446 35448
rect 23753 35445 23765 35448
rect 23799 35445 23811 35479
rect 23753 35439 23811 35445
rect 24397 35479 24455 35485
rect 24397 35445 24409 35479
rect 24443 35476 24455 35479
rect 24486 35476 24492 35488
rect 24443 35448 24492 35476
rect 24443 35445 24455 35448
rect 24397 35439 24455 35445
rect 24486 35436 24492 35448
rect 24544 35436 24550 35488
rect 28258 35436 28264 35488
rect 28316 35476 28322 35488
rect 28721 35479 28779 35485
rect 28721 35476 28733 35479
rect 28316 35448 28733 35476
rect 28316 35436 28322 35448
rect 28721 35445 28733 35448
rect 28767 35445 28779 35479
rect 28721 35439 28779 35445
rect 33042 35436 33048 35488
rect 33100 35476 33106 35488
rect 33321 35479 33379 35485
rect 33321 35476 33333 35479
rect 33100 35448 33333 35476
rect 33100 35436 33106 35448
rect 33321 35445 33333 35448
rect 33367 35445 33379 35479
rect 33321 35439 33379 35445
rect 34514 35436 34520 35488
rect 34572 35476 34578 35488
rect 35161 35479 35219 35485
rect 35161 35476 35173 35479
rect 34572 35448 35173 35476
rect 34572 35436 34578 35448
rect 35161 35445 35173 35448
rect 35207 35445 35219 35479
rect 35161 35439 35219 35445
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 11882 35272 11888 35284
rect 11843 35244 11888 35272
rect 11882 35232 11888 35244
rect 11940 35232 11946 35284
rect 17218 35232 17224 35284
rect 17276 35272 17282 35284
rect 27154 35272 27160 35284
rect 17276 35244 27160 35272
rect 17276 35232 17282 35244
rect 27154 35232 27160 35244
rect 27212 35232 27218 35284
rect 27430 35272 27436 35284
rect 27391 35244 27436 35272
rect 27430 35232 27436 35244
rect 27488 35232 27494 35284
rect 28534 35272 28540 35284
rect 28495 35244 28540 35272
rect 28534 35232 28540 35244
rect 28592 35232 28598 35284
rect 30926 35232 30932 35284
rect 30984 35272 30990 35284
rect 30984 35244 33456 35272
rect 30984 35232 30990 35244
rect 10502 35136 10508 35148
rect 4264 35108 6776 35136
rect 10463 35108 10508 35136
rect 4264 35077 4292 35108
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35037 4307 35071
rect 6178 35068 6184 35080
rect 6139 35040 6184 35068
rect 4249 35031 4307 35037
rect 6178 35028 6184 35040
rect 6236 35028 6242 35080
rect 6748 35012 6776 35108
rect 10502 35096 10508 35108
rect 10560 35096 10566 35148
rect 8294 35068 8300 35080
rect 7392 35040 8300 35068
rect 4433 35003 4491 35009
rect 4433 34969 4445 35003
rect 4479 35000 4491 35003
rect 4706 35000 4712 35012
rect 4479 34972 4712 35000
rect 4479 34969 4491 34972
rect 4433 34963 4491 34969
rect 4706 34960 4712 34972
rect 4764 35000 4770 35012
rect 5258 35000 5264 35012
rect 4764 34972 5264 35000
rect 4764 34960 4770 34972
rect 5258 34960 5264 34972
rect 5316 34960 5322 35012
rect 5442 34960 5448 35012
rect 5500 35000 5506 35012
rect 6365 35003 6423 35009
rect 6365 35000 6377 35003
rect 5500 34972 6377 35000
rect 5500 34960 5506 34972
rect 6365 34969 6377 34972
rect 6411 34969 6423 35003
rect 6365 34963 6423 34969
rect 4617 34935 4675 34941
rect 4617 34901 4629 34935
rect 4663 34932 4675 34935
rect 4798 34932 4804 34944
rect 4663 34904 4804 34932
rect 4663 34901 4675 34904
rect 4617 34895 4675 34901
rect 4798 34892 4804 34904
rect 4856 34892 4862 34944
rect 5074 34932 5080 34944
rect 5035 34904 5080 34932
rect 5074 34892 5080 34904
rect 5132 34892 5138 34944
rect 5994 34932 6000 34944
rect 5955 34904 6000 34932
rect 5994 34892 6000 34904
rect 6052 34892 6058 34944
rect 6380 34932 6408 34963
rect 6730 34960 6736 35012
rect 6788 35000 6794 35012
rect 7285 35003 7343 35009
rect 7285 35000 7297 35003
rect 6788 34972 7297 35000
rect 6788 34960 6794 34972
rect 7285 34969 7297 34972
rect 7331 34969 7343 35003
rect 7285 34963 7343 34969
rect 7392 34932 7420 35040
rect 8294 35028 8300 35040
rect 8352 35028 8358 35080
rect 11900 35068 11928 35232
rect 12897 35207 12955 35213
rect 12897 35173 12909 35207
rect 12943 35204 12955 35207
rect 17310 35204 17316 35216
rect 12943 35176 17316 35204
rect 12943 35173 12955 35176
rect 12897 35167 12955 35173
rect 17310 35164 17316 35176
rect 17368 35164 17374 35216
rect 30282 35164 30288 35216
rect 30340 35164 30346 35216
rect 12526 35096 12532 35148
rect 12584 35136 12590 35148
rect 18049 35139 18107 35145
rect 18049 35136 18061 35139
rect 12584 35108 12664 35136
rect 12584 35096 12590 35108
rect 12636 35077 12664 35108
rect 17052 35108 18061 35136
rect 12345 35071 12403 35077
rect 12345 35068 12357 35071
rect 11900 35040 12357 35068
rect 12345 35037 12357 35040
rect 12391 35037 12403 35071
rect 12345 35031 12403 35037
rect 12621 35071 12679 35077
rect 12621 35037 12633 35071
rect 12667 35037 12679 35071
rect 12621 35031 12679 35037
rect 12713 35071 12771 35077
rect 12713 35037 12725 35071
rect 12759 35068 12771 35071
rect 12802 35068 12808 35080
rect 12759 35040 12808 35068
rect 12759 35037 12771 35040
rect 12713 35031 12771 35037
rect 12802 35028 12808 35040
rect 12860 35028 12866 35080
rect 16850 35068 16856 35080
rect 16811 35040 16856 35068
rect 16850 35028 16856 35040
rect 16908 35028 16914 35080
rect 17052 35077 17080 35108
rect 18049 35105 18061 35108
rect 18095 35105 18107 35139
rect 28442 35136 28448 35148
rect 18049 35099 18107 35105
rect 27816 35108 28448 35136
rect 16945 35071 17003 35077
rect 16945 35037 16957 35071
rect 16991 35037 17003 35071
rect 16945 35031 17003 35037
rect 17037 35071 17095 35077
rect 17037 35037 17049 35071
rect 17083 35037 17095 35071
rect 17037 35031 17095 35037
rect 7469 35003 7527 35009
rect 7469 34969 7481 35003
rect 7515 35000 7527 35003
rect 8570 35000 8576 35012
rect 7515 34972 8576 35000
rect 7515 34969 7527 34972
rect 7469 34963 7527 34969
rect 8570 34960 8576 34972
rect 8628 34960 8634 35012
rect 10772 35003 10830 35009
rect 10772 34969 10784 35003
rect 10818 35000 10830 35003
rect 11146 35000 11152 35012
rect 10818 34972 11152 35000
rect 10818 34969 10830 34972
rect 10772 34963 10830 34969
rect 11146 34960 11152 34972
rect 11204 34960 11210 35012
rect 12434 34960 12440 35012
rect 12492 35000 12498 35012
rect 12529 35003 12587 35009
rect 12529 35000 12541 35003
rect 12492 34972 12541 35000
rect 12492 34960 12498 34972
rect 12529 34969 12541 34972
rect 12575 34969 12587 35003
rect 12529 34963 12587 34969
rect 16666 34960 16672 35012
rect 16724 35000 16730 35012
rect 16960 35000 16988 35031
rect 17126 35028 17132 35080
rect 17184 35068 17190 35080
rect 17221 35071 17279 35077
rect 17221 35068 17233 35071
rect 17184 35040 17233 35068
rect 17184 35028 17190 35040
rect 17221 35037 17233 35040
rect 17267 35037 17279 35071
rect 17678 35068 17684 35080
rect 17639 35040 17684 35068
rect 17221 35031 17279 35037
rect 17678 35028 17684 35040
rect 17736 35028 17742 35080
rect 19334 35068 19340 35080
rect 19295 35040 19340 35068
rect 19334 35028 19340 35040
rect 19392 35028 19398 35080
rect 19426 35028 19432 35080
rect 19484 35068 19490 35080
rect 20070 35068 20076 35080
rect 19484 35040 20076 35068
rect 19484 35028 19490 35040
rect 20070 35028 20076 35040
rect 20128 35068 20134 35080
rect 27816 35077 27844 35108
rect 28442 35096 28448 35108
rect 28500 35136 28506 35148
rect 29730 35136 29736 35148
rect 28500 35108 29736 35136
rect 28500 35096 28506 35108
rect 29730 35096 29736 35108
rect 29788 35136 29794 35148
rect 30300 35136 30328 35164
rect 33318 35136 33324 35148
rect 29788 35108 30236 35136
rect 30300 35108 30972 35136
rect 29788 35096 29794 35108
rect 20257 35071 20315 35077
rect 20257 35068 20269 35071
rect 20128 35040 20269 35068
rect 20128 35028 20134 35040
rect 20257 35037 20269 35040
rect 20303 35037 20315 35071
rect 22465 35071 22523 35077
rect 22465 35068 22477 35071
rect 20257 35031 20315 35037
rect 21560 35040 22477 35068
rect 17862 35000 17868 35012
rect 16724 34972 16988 35000
rect 17823 34972 17868 35000
rect 16724 34960 16730 34972
rect 17862 34960 17868 34972
rect 17920 34960 17926 35012
rect 6380 34904 7420 34932
rect 7653 34935 7711 34941
rect 7653 34901 7665 34935
rect 7699 34932 7711 34935
rect 7926 34932 7932 34944
rect 7699 34904 7932 34932
rect 7699 34901 7711 34904
rect 7653 34895 7711 34901
rect 7926 34892 7932 34904
rect 7984 34892 7990 34944
rect 16577 34935 16635 34941
rect 16577 34901 16589 34935
rect 16623 34932 16635 34935
rect 16758 34932 16764 34944
rect 16623 34904 16764 34932
rect 16623 34901 16635 34904
rect 16577 34895 16635 34901
rect 16758 34892 16764 34904
rect 16816 34892 16822 34944
rect 19334 34892 19340 34944
rect 19392 34932 19398 34944
rect 19429 34935 19487 34941
rect 19429 34932 19441 34935
rect 19392 34904 19441 34932
rect 19392 34892 19398 34904
rect 19429 34901 19441 34904
rect 19475 34932 19487 34935
rect 19518 34932 19524 34944
rect 19475 34904 19524 34932
rect 19475 34901 19487 34904
rect 19429 34895 19487 34901
rect 19518 34892 19524 34904
rect 19576 34892 19582 34944
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 21560 34941 21588 35040
rect 22465 35037 22477 35040
rect 22511 35037 22523 35071
rect 27663 35071 27721 35077
rect 27663 35068 27675 35071
rect 22465 35031 22523 35037
rect 26988 35040 27675 35068
rect 22370 34960 22376 35012
rect 22428 35000 22434 35012
rect 22710 35003 22768 35009
rect 22710 35000 22722 35003
rect 22428 34972 22722 35000
rect 22428 34960 22434 34972
rect 22710 34969 22722 34972
rect 22756 34969 22768 35003
rect 22710 34963 22768 34969
rect 26988 34944 27016 35040
rect 27663 35037 27675 35040
rect 27709 35037 27721 35071
rect 27663 35031 27721 35037
rect 27801 35071 27859 35077
rect 27801 35037 27813 35071
rect 27847 35037 27859 35071
rect 27801 35031 27859 35037
rect 27893 35071 27951 35077
rect 27893 35037 27905 35071
rect 27939 35068 27951 35071
rect 27982 35068 27988 35080
rect 27939 35040 27988 35068
rect 27939 35037 27951 35040
rect 27893 35031 27951 35037
rect 27982 35028 27988 35040
rect 28040 35028 28046 35080
rect 28074 35028 28080 35080
rect 28132 35068 28138 35080
rect 28905 35071 28963 35077
rect 28132 35040 28177 35068
rect 28132 35028 28138 35040
rect 28905 35037 28917 35071
rect 28951 35068 28963 35071
rect 29546 35068 29552 35080
rect 28951 35040 29552 35068
rect 28951 35037 28963 35040
rect 28905 35031 28963 35037
rect 29546 35028 29552 35040
rect 29604 35028 29610 35080
rect 29914 35028 29920 35080
rect 29972 35068 29978 35080
rect 30208 35077 30236 35108
rect 30055 35071 30113 35077
rect 30055 35068 30067 35071
rect 29972 35040 30067 35068
rect 29972 35028 29978 35040
rect 30055 35037 30067 35040
rect 30101 35037 30113 35071
rect 30055 35031 30113 35037
rect 30193 35071 30251 35077
rect 30193 35037 30205 35071
rect 30239 35037 30251 35071
rect 30193 35031 30251 35037
rect 30306 35071 30364 35077
rect 30306 35037 30318 35071
rect 30352 35068 30364 35071
rect 30469 35071 30527 35077
rect 30352 35040 30420 35068
rect 30352 35037 30364 35040
rect 30306 35031 30364 35037
rect 28626 34960 28632 35012
rect 28684 35000 28690 35012
rect 28721 35003 28779 35009
rect 28721 35000 28733 35003
rect 28684 34972 28733 35000
rect 28684 34960 28690 34972
rect 28721 34969 28733 34972
rect 28767 34969 28779 35003
rect 30392 35000 30420 35040
rect 30469 35037 30481 35071
rect 30515 35068 30527 35071
rect 30558 35068 30564 35080
rect 30515 35040 30564 35068
rect 30515 35037 30527 35040
rect 30469 35031 30527 35037
rect 30558 35028 30564 35040
rect 30616 35028 30622 35080
rect 30944 35077 30972 35108
rect 32876 35108 33324 35136
rect 30929 35071 30987 35077
rect 30929 35037 30941 35071
rect 30975 35068 30987 35071
rect 32876 35068 32904 35108
rect 33318 35096 33324 35108
rect 33376 35096 33382 35148
rect 30975 35040 32904 35068
rect 33229 35071 33287 35077
rect 30975 35037 30987 35040
rect 30929 35031 30987 35037
rect 33229 35037 33241 35071
rect 33275 35068 33287 35071
rect 33428 35068 33456 35244
rect 33502 35096 33508 35148
rect 33560 35136 33566 35148
rect 33560 35108 33605 35136
rect 33560 35096 33566 35108
rect 58158 35068 58164 35080
rect 33275 35040 33456 35068
rect 58119 35040 58164 35068
rect 33275 35037 33287 35040
rect 33229 35031 33287 35037
rect 58158 35028 58164 35040
rect 58216 35028 58222 35080
rect 30834 35000 30840 35012
rect 30392 34972 30840 35000
rect 28721 34963 28779 34969
rect 30834 34960 30840 34972
rect 30892 34960 30898 35012
rect 31174 35003 31232 35009
rect 31174 35000 31186 35003
rect 31036 34972 31186 35000
rect 21545 34935 21603 34941
rect 21545 34932 21557 34935
rect 20772 34904 21557 34932
rect 20772 34892 20778 34904
rect 21545 34901 21557 34904
rect 21591 34901 21603 34935
rect 21545 34895 21603 34901
rect 22094 34892 22100 34944
rect 22152 34932 22158 34944
rect 23845 34935 23903 34941
rect 23845 34932 23857 34935
rect 22152 34904 23857 34932
rect 22152 34892 22158 34904
rect 23845 34901 23857 34904
rect 23891 34901 23903 34935
rect 26970 34932 26976 34944
rect 26931 34904 26976 34932
rect 23845 34895 23903 34901
rect 26970 34892 26976 34904
rect 27028 34892 27034 34944
rect 29825 34935 29883 34941
rect 29825 34901 29837 34935
rect 29871 34932 29883 34935
rect 31036 34932 31064 34972
rect 31174 34969 31186 34972
rect 31220 34969 31232 35003
rect 31174 34963 31232 34969
rect 29871 34904 31064 34932
rect 32309 34935 32367 34941
rect 29871 34901 29883 34904
rect 29825 34895 29883 34901
rect 32309 34901 32321 34935
rect 32355 34932 32367 34935
rect 32398 34932 32404 34944
rect 32355 34904 32404 34932
rect 32355 34901 32367 34904
rect 32309 34895 32367 34901
rect 32398 34892 32404 34904
rect 32456 34892 32462 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 2774 34728 2780 34740
rect 2516 34700 2780 34728
rect 2516 34601 2544 34700
rect 2774 34688 2780 34700
rect 2832 34688 2838 34740
rect 4062 34688 4068 34740
rect 4120 34728 4126 34740
rect 4341 34731 4399 34737
rect 4341 34728 4353 34731
rect 4120 34700 4353 34728
rect 4120 34688 4126 34700
rect 4341 34697 4353 34700
rect 4387 34697 4399 34731
rect 8570 34728 8576 34740
rect 8531 34700 8576 34728
rect 4341 34691 4399 34697
rect 8570 34688 8576 34700
rect 8628 34688 8634 34740
rect 11977 34731 12035 34737
rect 11977 34697 11989 34731
rect 12023 34728 12035 34731
rect 12066 34728 12072 34740
rect 12023 34700 12072 34728
rect 12023 34697 12035 34700
rect 11977 34691 12035 34697
rect 12066 34688 12072 34700
rect 12124 34688 12130 34740
rect 17218 34728 17224 34740
rect 12406 34700 17224 34728
rect 6457 34663 6515 34669
rect 6457 34660 6469 34663
rect 4632 34632 6469 34660
rect 4632 34604 4660 34632
rect 6457 34629 6469 34632
rect 6503 34660 6515 34663
rect 12406 34660 12434 34700
rect 17218 34688 17224 34700
rect 17276 34688 17282 34740
rect 17494 34688 17500 34740
rect 17552 34728 17558 34740
rect 17862 34728 17868 34740
rect 17552 34700 17868 34728
rect 17552 34688 17558 34700
rect 17862 34688 17868 34700
rect 17920 34728 17926 34740
rect 18049 34731 18107 34737
rect 18049 34728 18061 34731
rect 17920 34700 18061 34728
rect 17920 34688 17926 34700
rect 18049 34697 18061 34700
rect 18095 34697 18107 34731
rect 20070 34728 20076 34740
rect 20031 34700 20076 34728
rect 18049 34691 18107 34697
rect 20070 34688 20076 34700
rect 20128 34688 20134 34740
rect 27982 34728 27988 34740
rect 27943 34700 27988 34728
rect 27982 34688 27988 34700
rect 28040 34688 28046 34740
rect 29178 34688 29184 34740
rect 29236 34728 29242 34740
rect 29273 34731 29331 34737
rect 29273 34728 29285 34731
rect 29236 34700 29285 34728
rect 29236 34688 29242 34700
rect 29273 34697 29285 34700
rect 29319 34728 29331 34731
rect 29914 34728 29920 34740
rect 29319 34700 29920 34728
rect 29319 34697 29331 34700
rect 29273 34691 29331 34697
rect 29914 34688 29920 34700
rect 29972 34688 29978 34740
rect 33134 34728 33140 34740
rect 33095 34700 33140 34728
rect 33134 34688 33140 34700
rect 33192 34688 33198 34740
rect 34241 34731 34299 34737
rect 34241 34697 34253 34731
rect 34287 34728 34299 34731
rect 34790 34728 34796 34740
rect 34287 34700 34796 34728
rect 34287 34697 34299 34700
rect 34241 34691 34299 34697
rect 34790 34688 34796 34700
rect 34848 34688 34854 34740
rect 20714 34660 20720 34672
rect 6503 34632 12434 34660
rect 16684 34632 20720 34660
rect 6503 34629 6515 34632
rect 6457 34623 6515 34629
rect 2501 34595 2559 34601
rect 2501 34561 2513 34595
rect 2547 34561 2559 34595
rect 2501 34555 2559 34561
rect 2768 34595 2826 34601
rect 2768 34561 2780 34595
rect 2814 34592 2826 34595
rect 3786 34592 3792 34604
rect 2814 34564 3792 34592
rect 2814 34561 2826 34564
rect 2768 34555 2826 34561
rect 3786 34552 3792 34564
rect 3844 34552 3850 34604
rect 4614 34592 4620 34604
rect 4527 34564 4620 34592
rect 4614 34552 4620 34564
rect 4672 34552 4678 34604
rect 4706 34595 4764 34601
rect 4706 34561 4718 34595
rect 4752 34561 4764 34595
rect 4706 34555 4764 34561
rect 4724 34524 4752 34555
rect 4798 34552 4804 34604
rect 4856 34592 4862 34604
rect 4985 34595 5043 34601
rect 4856 34564 4901 34592
rect 4856 34552 4862 34564
rect 4985 34561 4997 34595
rect 5031 34592 5043 34595
rect 5074 34592 5080 34604
rect 5031 34564 5080 34592
rect 5031 34561 5043 34564
rect 4985 34555 5043 34561
rect 5074 34552 5080 34564
rect 5132 34552 5138 34604
rect 6086 34552 6092 34604
rect 6144 34592 6150 34604
rect 6822 34592 6828 34604
rect 6144 34564 6828 34592
rect 6144 34552 6150 34564
rect 6822 34552 6828 34564
rect 6880 34592 6886 34604
rect 7466 34601 7472 34604
rect 7193 34595 7251 34601
rect 7193 34592 7205 34595
rect 6880 34564 7205 34592
rect 6880 34552 6886 34564
rect 7193 34561 7205 34564
rect 7239 34561 7251 34595
rect 7193 34555 7251 34561
rect 7460 34555 7472 34601
rect 7524 34592 7530 34604
rect 7524 34564 7560 34592
rect 7466 34552 7472 34555
rect 7524 34552 7530 34564
rect 10226 34552 10232 34604
rect 10284 34592 10290 34604
rect 10321 34595 10379 34601
rect 10321 34592 10333 34595
rect 10284 34564 10333 34592
rect 10284 34552 10290 34564
rect 10321 34561 10333 34564
rect 10367 34561 10379 34595
rect 10321 34555 10379 34561
rect 12066 34552 12072 34604
rect 12124 34592 12130 34604
rect 16684 34601 16712 34632
rect 20714 34620 20720 34632
rect 20772 34620 20778 34672
rect 27065 34663 27123 34669
rect 27065 34660 27077 34663
rect 22066 34632 27077 34660
rect 12529 34595 12587 34601
rect 12529 34592 12541 34595
rect 12124 34564 12541 34592
rect 12124 34552 12130 34564
rect 12529 34561 12541 34564
rect 12575 34561 12587 34595
rect 12529 34555 12587 34561
rect 16669 34595 16727 34601
rect 16669 34561 16681 34595
rect 16715 34561 16727 34595
rect 16669 34555 16727 34561
rect 16758 34552 16764 34604
rect 16816 34592 16822 34604
rect 16925 34595 16983 34601
rect 16925 34592 16937 34595
rect 16816 34564 16937 34592
rect 16816 34552 16822 34564
rect 16925 34561 16937 34564
rect 16971 34561 16983 34595
rect 19150 34592 19156 34604
rect 19111 34564 19156 34592
rect 16925 34555 16983 34561
rect 19150 34552 19156 34564
rect 19208 34552 19214 34604
rect 19337 34595 19395 34601
rect 19337 34561 19349 34595
rect 19383 34592 19395 34595
rect 19426 34592 19432 34604
rect 19383 34564 19432 34592
rect 19383 34561 19395 34564
rect 19337 34555 19395 34561
rect 19426 34552 19432 34564
rect 19484 34552 19490 34604
rect 4890 34524 4896 34536
rect 4724 34496 4896 34524
rect 4890 34484 4896 34496
rect 4948 34484 4954 34536
rect 10594 34524 10600 34536
rect 10555 34496 10600 34524
rect 10594 34484 10600 34496
rect 10652 34484 10658 34536
rect 12713 34527 12771 34533
rect 12713 34493 12725 34527
rect 12759 34524 12771 34527
rect 13170 34524 13176 34536
rect 12759 34496 13176 34524
rect 12759 34493 12771 34496
rect 12713 34487 12771 34493
rect 13170 34484 13176 34496
rect 13228 34524 13234 34536
rect 22066 34524 22094 34632
rect 27065 34629 27077 34632
rect 27111 34660 27123 34663
rect 27614 34660 27620 34672
rect 27111 34632 27620 34660
rect 27111 34629 27123 34632
rect 27065 34623 27123 34629
rect 27614 34620 27620 34632
rect 27672 34660 27678 34672
rect 28074 34660 28080 34672
rect 27672 34632 28080 34660
rect 27672 34620 27678 34632
rect 28074 34620 28080 34632
rect 28132 34620 28138 34672
rect 28353 34663 28411 34669
rect 28353 34629 28365 34663
rect 28399 34660 28411 34663
rect 29546 34660 29552 34672
rect 28399 34632 29552 34660
rect 28399 34629 28411 34632
rect 28353 34623 28411 34629
rect 29546 34620 29552 34632
rect 29604 34620 29610 34672
rect 33502 34620 33508 34672
rect 33560 34660 33566 34672
rect 33560 34632 33916 34660
rect 33560 34620 33566 34632
rect 24118 34592 24124 34604
rect 24176 34601 24182 34604
rect 24088 34564 24124 34592
rect 24118 34552 24124 34564
rect 24176 34555 24188 34601
rect 24854 34592 24860 34604
rect 24815 34564 24860 34592
rect 24176 34552 24182 34555
rect 24854 34552 24860 34564
rect 24912 34552 24918 34604
rect 25038 34592 25044 34604
rect 24999 34564 25044 34592
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 28166 34592 28172 34604
rect 28127 34564 28172 34592
rect 28166 34552 28172 34564
rect 28224 34552 28230 34604
rect 31570 34552 31576 34604
rect 31628 34592 31634 34604
rect 32953 34595 33011 34601
rect 32953 34592 32965 34595
rect 31628 34564 32965 34592
rect 31628 34552 31634 34564
rect 32953 34561 32965 34564
rect 32999 34561 33011 34595
rect 33594 34592 33600 34604
rect 33555 34564 33600 34592
rect 32953 34555 33011 34561
rect 33594 34552 33600 34564
rect 33652 34552 33658 34604
rect 33778 34592 33784 34604
rect 33739 34564 33784 34592
rect 33778 34552 33784 34564
rect 33836 34552 33842 34604
rect 33888 34601 33916 34632
rect 33873 34595 33931 34601
rect 33873 34561 33885 34595
rect 33919 34561 33931 34595
rect 33873 34555 33931 34561
rect 33965 34595 34023 34601
rect 33965 34561 33977 34595
rect 34011 34561 34023 34595
rect 33965 34555 34023 34561
rect 13228 34496 16712 34524
rect 13228 34484 13234 34496
rect 11808 34428 12434 34456
rect 3881 34391 3939 34397
rect 3881 34357 3893 34391
rect 3927 34388 3939 34391
rect 4982 34388 4988 34400
rect 3927 34360 4988 34388
rect 3927 34357 3939 34360
rect 3881 34351 3939 34357
rect 4982 34348 4988 34360
rect 5040 34348 5046 34400
rect 5074 34348 5080 34400
rect 5132 34388 5138 34400
rect 5445 34391 5503 34397
rect 5445 34388 5457 34391
rect 5132 34360 5457 34388
rect 5132 34348 5138 34360
rect 5445 34357 5457 34360
rect 5491 34357 5503 34391
rect 5445 34351 5503 34357
rect 7098 34348 7104 34400
rect 7156 34388 7162 34400
rect 11808 34388 11836 34428
rect 7156 34360 11836 34388
rect 12406 34388 12434 34428
rect 12526 34388 12532 34400
rect 12406 34360 12532 34388
rect 7156 34348 7162 34360
rect 12526 34348 12532 34360
rect 12584 34348 12590 34400
rect 16684 34388 16712 34496
rect 17696 34496 22094 34524
rect 24397 34527 24455 34533
rect 17696 34388 17724 34496
rect 24397 34493 24409 34527
rect 24443 34524 24455 34527
rect 26234 34524 26240 34536
rect 24443 34496 26240 34524
rect 24443 34493 24455 34496
rect 24397 34487 24455 34493
rect 26234 34484 26240 34496
rect 26292 34524 26298 34536
rect 27338 34524 27344 34536
rect 26292 34496 27344 34524
rect 26292 34484 26298 34496
rect 27338 34484 27344 34496
rect 27396 34524 27402 34536
rect 27522 34524 27528 34536
rect 27396 34496 27528 34524
rect 27396 34484 27402 34496
rect 27522 34484 27528 34496
rect 27580 34484 27586 34536
rect 29822 34524 29828 34536
rect 29783 34496 29828 34524
rect 29822 34484 29828 34496
rect 29880 34524 29886 34536
rect 30285 34527 30343 34533
rect 30285 34524 30297 34527
rect 29880 34496 30297 34524
rect 29880 34484 29886 34496
rect 30285 34493 30297 34496
rect 30331 34493 30343 34527
rect 30558 34524 30564 34536
rect 30519 34496 30564 34524
rect 30285 34487 30343 34493
rect 30558 34484 30564 34496
rect 30616 34484 30622 34536
rect 33410 34484 33416 34536
rect 33468 34524 33474 34536
rect 33980 34524 34008 34555
rect 33468 34496 34008 34524
rect 33468 34484 33474 34496
rect 24486 34416 24492 34468
rect 24544 34456 24550 34468
rect 35342 34456 35348 34468
rect 24544 34428 35348 34456
rect 24544 34416 24550 34428
rect 35342 34416 35348 34428
rect 35400 34416 35406 34468
rect 16684 34360 17724 34388
rect 19334 34348 19340 34400
rect 19392 34388 19398 34400
rect 19521 34391 19579 34397
rect 19521 34388 19533 34391
rect 19392 34360 19533 34388
rect 19392 34348 19398 34360
rect 19521 34357 19533 34360
rect 19567 34357 19579 34391
rect 23014 34388 23020 34400
rect 22975 34360 23020 34388
rect 19521 34351 19579 34357
rect 23014 34348 23020 34360
rect 23072 34348 23078 34400
rect 25222 34388 25228 34400
rect 25183 34360 25228 34388
rect 25222 34348 25228 34360
rect 25280 34348 25286 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 3786 34184 3792 34196
rect 3747 34156 3792 34184
rect 3786 34144 3792 34156
rect 3844 34144 3850 34196
rect 5626 34184 5632 34196
rect 5587 34156 5632 34184
rect 5626 34144 5632 34156
rect 5684 34144 5690 34196
rect 7009 34187 7067 34193
rect 7009 34153 7021 34187
rect 7055 34184 7067 34187
rect 7098 34184 7104 34196
rect 7055 34156 7104 34184
rect 7055 34153 7067 34156
rect 7009 34147 7067 34153
rect 7098 34144 7104 34156
rect 7156 34144 7162 34196
rect 7466 34184 7472 34196
rect 7427 34156 7472 34184
rect 7466 34144 7472 34156
rect 7524 34144 7530 34196
rect 11146 34184 11152 34196
rect 11107 34156 11152 34184
rect 11146 34144 11152 34156
rect 11204 34144 11210 34196
rect 12526 34144 12532 34196
rect 12584 34184 12590 34196
rect 29178 34184 29184 34196
rect 12584 34156 29184 34184
rect 12584 34144 12590 34156
rect 29178 34144 29184 34156
rect 29236 34144 29242 34196
rect 35342 34184 35348 34196
rect 35303 34156 35348 34184
rect 35342 34144 35348 34156
rect 35400 34144 35406 34196
rect 13722 34116 13728 34128
rect 9232 34088 13728 34116
rect 3418 34008 3424 34060
rect 3476 34048 3482 34060
rect 7650 34048 7656 34060
rect 3476 34020 7656 34048
rect 3476 34008 3482 34020
rect 3142 33940 3148 33992
rect 3200 33980 3206 33992
rect 3237 33983 3295 33989
rect 3237 33980 3249 33983
rect 3200 33952 3249 33980
rect 3200 33940 3206 33952
rect 3237 33949 3249 33952
rect 3283 33980 3295 33983
rect 4062 33980 4068 33992
rect 3283 33952 4068 33980
rect 3283 33949 3295 33952
rect 3237 33943 3295 33949
rect 4062 33940 4068 33952
rect 4120 33940 4126 33992
rect 4157 33983 4215 33989
rect 4157 33949 4169 33983
rect 4203 33949 4215 33983
rect 4157 33943 4215 33949
rect 4172 33912 4200 33943
rect 4246 33940 4252 33992
rect 4304 33980 4310 33992
rect 4433 33983 4491 33989
rect 4304 33952 4349 33980
rect 4304 33940 4310 33952
rect 4433 33949 4445 33983
rect 4479 33980 4491 33983
rect 5074 33980 5080 33992
rect 4479 33952 5080 33980
rect 4479 33949 4491 33952
rect 4433 33943 4491 33949
rect 5074 33940 5080 33952
rect 5132 33940 5138 33992
rect 5169 33983 5227 33989
rect 5169 33949 5181 33983
rect 5215 33980 5227 33983
rect 5902 33980 5908 33992
rect 5215 33952 5908 33980
rect 5215 33949 5227 33952
rect 5169 33943 5227 33949
rect 5902 33940 5908 33952
rect 5960 33940 5966 33992
rect 6012 33989 6040 34020
rect 7650 34008 7656 34020
rect 7708 34008 7714 34060
rect 8202 34008 8208 34060
rect 8260 34048 8266 34060
rect 8260 34020 9076 34048
rect 8260 34008 8266 34020
rect 5997 33983 6055 33989
rect 5997 33949 6009 33983
rect 6043 33949 6055 33983
rect 5997 33943 6055 33949
rect 6086 33940 6092 33992
rect 6144 33980 6150 33992
rect 6273 33983 6331 33989
rect 6144 33952 6189 33980
rect 6144 33940 6150 33952
rect 6273 33949 6285 33983
rect 6319 33949 6331 33983
rect 6273 33943 6331 33949
rect 4890 33912 4896 33924
rect 4172 33884 4896 33912
rect 4890 33872 4896 33884
rect 4948 33872 4954 33924
rect 6288 33912 6316 33943
rect 7098 33940 7104 33992
rect 7156 33980 7162 33992
rect 7745 33983 7803 33989
rect 7745 33980 7757 33983
rect 7156 33952 7757 33980
rect 7156 33940 7162 33952
rect 7745 33949 7757 33952
rect 7791 33949 7803 33983
rect 7745 33943 7803 33949
rect 7834 33980 7892 33986
rect 7834 33946 7846 33980
rect 7880 33946 7892 33980
rect 7834 33940 7892 33946
rect 7926 33940 7932 33992
rect 7984 33989 7990 33992
rect 7984 33980 7992 33989
rect 8113 33983 8171 33989
rect 7984 33952 8029 33980
rect 7984 33943 7992 33952
rect 8113 33949 8125 33983
rect 8159 33949 8171 33983
rect 8938 33980 8944 33992
rect 8899 33952 8944 33980
rect 8113 33943 8171 33949
rect 7984 33940 7990 33943
rect 6196 33884 6316 33912
rect 7849 33912 7877 33940
rect 8018 33912 8024 33924
rect 7849 33884 8024 33912
rect 6196 33856 6224 33884
rect 8018 33872 8024 33884
rect 8076 33872 8082 33924
rect 3326 33804 3332 33856
rect 3384 33844 3390 33856
rect 6178 33844 6184 33856
rect 3384 33816 6184 33844
rect 3384 33804 3390 33816
rect 6178 33804 6184 33816
rect 6236 33804 6242 33856
rect 8128 33844 8156 33943
rect 8938 33940 8944 33952
rect 8996 33940 9002 33992
rect 9048 33989 9076 34020
rect 9232 33989 9260 34088
rect 13722 34076 13728 34088
rect 13780 34076 13786 34128
rect 16850 34116 16856 34128
rect 14292 34088 16856 34116
rect 9858 34008 9864 34060
rect 9916 34048 9922 34060
rect 10410 34048 10416 34060
rect 9916 34020 10416 34048
rect 9916 34008 9922 34020
rect 10410 34008 10416 34020
rect 10468 34048 10474 34060
rect 11701 34051 11759 34057
rect 10468 34020 10824 34048
rect 10468 34008 10474 34020
rect 9034 33983 9092 33989
rect 9034 33949 9046 33983
rect 9080 33949 9092 33983
rect 9034 33943 9092 33949
rect 9217 33983 9275 33989
rect 9217 33949 9229 33983
rect 9263 33949 9275 33983
rect 9217 33943 9275 33949
rect 9447 33983 9505 33989
rect 9447 33949 9459 33983
rect 9493 33980 9505 33983
rect 10134 33980 10140 33992
rect 9493 33952 10140 33980
rect 9493 33949 9505 33952
rect 9447 33943 9505 33949
rect 10134 33940 10140 33952
rect 10192 33940 10198 33992
rect 10226 33940 10232 33992
rect 10284 33980 10290 33992
rect 10505 33983 10563 33989
rect 10505 33980 10517 33983
rect 10284 33952 10517 33980
rect 10284 33940 10290 33952
rect 10505 33949 10517 33952
rect 10551 33949 10563 33983
rect 10686 33980 10692 33992
rect 10647 33952 10692 33980
rect 10505 33943 10563 33949
rect 10686 33940 10692 33952
rect 10744 33940 10750 33992
rect 10796 33989 10824 34020
rect 11701 34017 11713 34051
rect 11747 34048 11759 34051
rect 14292 34048 14320 34088
rect 16850 34076 16856 34088
rect 16908 34076 16914 34128
rect 17957 34119 18015 34125
rect 17957 34085 17969 34119
rect 18003 34085 18015 34119
rect 17957 34079 18015 34085
rect 24504 34088 25636 34116
rect 11747 34020 14320 34048
rect 14369 34051 14427 34057
rect 11747 34017 11759 34020
rect 11701 34011 11759 34017
rect 14369 34017 14381 34051
rect 14415 34048 14427 34051
rect 14642 34048 14648 34060
rect 14415 34020 14648 34048
rect 14415 34017 14427 34020
rect 14369 34011 14427 34017
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33949 10839 33983
rect 10781 33943 10839 33949
rect 10873 33983 10931 33989
rect 10873 33949 10885 33983
rect 10919 33980 10931 33983
rect 11716 33980 11744 34011
rect 14642 34008 14648 34020
rect 14700 34008 14706 34060
rect 10919 33952 11744 33980
rect 10919 33949 10931 33952
rect 10873 33943 10931 33949
rect 13722 33940 13728 33992
rect 13780 33980 13786 33992
rect 14093 33983 14151 33989
rect 13780 33952 14044 33980
rect 13780 33940 13786 33952
rect 8570 33872 8576 33924
rect 8628 33912 8634 33924
rect 9309 33915 9367 33921
rect 9309 33912 9321 33915
rect 8628 33884 9321 33912
rect 8628 33872 8634 33884
rect 9309 33881 9321 33884
rect 9355 33881 9367 33915
rect 9309 33875 9367 33881
rect 9416 33884 9720 33912
rect 8294 33844 8300 33856
rect 8128 33816 8300 33844
rect 8294 33804 8300 33816
rect 8352 33844 8358 33856
rect 9416 33844 9444 33884
rect 9582 33844 9588 33856
rect 8352 33816 9444 33844
rect 9543 33816 9588 33844
rect 8352 33804 8358 33816
rect 9582 33804 9588 33816
rect 9640 33804 9646 33856
rect 9692 33844 9720 33884
rect 10594 33872 10600 33924
rect 10652 33912 10658 33924
rect 13357 33915 13415 33921
rect 13357 33912 13369 33915
rect 10652 33884 13369 33912
rect 10652 33872 10658 33884
rect 13357 33881 13369 33884
rect 13403 33881 13415 33915
rect 13357 33875 13415 33881
rect 13541 33915 13599 33921
rect 13541 33881 13553 33915
rect 13587 33912 13599 33915
rect 13906 33912 13912 33924
rect 13587 33884 13912 33912
rect 13587 33881 13599 33884
rect 13541 33875 13599 33881
rect 13906 33872 13912 33884
rect 13964 33872 13970 33924
rect 14016 33912 14044 33952
rect 14093 33949 14105 33983
rect 14139 33980 14151 33983
rect 14182 33980 14188 33992
rect 14139 33952 14188 33980
rect 14139 33949 14151 33952
rect 14093 33943 14151 33949
rect 14182 33940 14188 33952
rect 14240 33940 14246 33992
rect 17310 33980 17316 33992
rect 17271 33952 17316 33980
rect 17310 33940 17316 33952
rect 17368 33940 17374 33992
rect 17494 33989 17500 33992
rect 17461 33983 17500 33989
rect 17461 33949 17473 33983
rect 17461 33943 17500 33949
rect 17494 33940 17500 33943
rect 17552 33940 17558 33992
rect 17770 33940 17776 33992
rect 17828 33989 17834 33992
rect 17828 33980 17836 33989
rect 17972 33980 18000 34079
rect 20714 34048 20720 34060
rect 20675 34020 20720 34048
rect 20714 34008 20720 34020
rect 20772 34008 20778 34060
rect 22370 34008 22376 34060
rect 22428 34048 22434 34060
rect 22646 34048 22652 34060
rect 22428 34020 22652 34048
rect 22428 34008 22434 34020
rect 22646 34008 22652 34020
rect 22704 34048 22710 34060
rect 22704 34020 23612 34048
rect 22704 34008 22710 34020
rect 20162 33980 20168 33992
rect 17828 33952 17873 33980
rect 17972 33952 20168 33980
rect 17828 33943 17836 33952
rect 17828 33940 17834 33943
rect 20162 33940 20168 33952
rect 20220 33940 20226 33992
rect 23382 33980 23388 33992
rect 22756 33952 23388 33980
rect 16025 33915 16083 33921
rect 16025 33912 16037 33915
rect 14016 33884 16037 33912
rect 16025 33881 16037 33884
rect 16071 33881 16083 33915
rect 16025 33875 16083 33881
rect 16209 33915 16267 33921
rect 16209 33881 16221 33915
rect 16255 33912 16267 33915
rect 16574 33912 16580 33924
rect 16255 33884 16580 33912
rect 16255 33881 16267 33884
rect 16209 33875 16267 33881
rect 16574 33872 16580 33884
rect 16632 33912 16638 33924
rect 17589 33915 17647 33921
rect 17589 33912 17601 33915
rect 16632 33884 17601 33912
rect 16632 33872 16638 33884
rect 17589 33881 17601 33884
rect 17635 33881 17647 33915
rect 17589 33875 17647 33881
rect 17681 33915 17739 33921
rect 17681 33881 17693 33915
rect 17727 33912 17739 33915
rect 19426 33912 19432 33924
rect 17727 33884 19432 33912
rect 17727 33881 17739 33884
rect 17681 33875 17739 33881
rect 19242 33844 19248 33856
rect 9692 33816 19248 33844
rect 19242 33804 19248 33816
rect 19300 33804 19306 33856
rect 19352 33853 19380 33884
rect 19426 33872 19432 33884
rect 19484 33872 19490 33924
rect 19978 33872 19984 33924
rect 20036 33912 20042 33924
rect 20450 33915 20508 33921
rect 20450 33912 20462 33915
rect 20036 33884 20462 33912
rect 20036 33872 20042 33884
rect 20450 33881 20462 33884
rect 20496 33881 20508 33915
rect 20450 33875 20508 33881
rect 22756 33856 22784 33952
rect 23382 33940 23388 33952
rect 23440 33940 23446 33992
rect 23584 33989 23612 34020
rect 23569 33983 23627 33989
rect 23569 33949 23581 33983
rect 23615 33949 23627 33983
rect 23569 33943 23627 33949
rect 23753 33983 23811 33989
rect 23753 33949 23765 33983
rect 23799 33980 23811 33983
rect 24302 33980 24308 33992
rect 23799 33952 24308 33980
rect 23799 33949 23811 33952
rect 23753 33943 23811 33949
rect 24302 33940 24308 33952
rect 24360 33940 24366 33992
rect 23014 33872 23020 33924
rect 23072 33912 23078 33924
rect 23477 33915 23535 33921
rect 23477 33912 23489 33915
rect 23072 33884 23489 33912
rect 23072 33872 23078 33884
rect 23477 33881 23489 33884
rect 23523 33881 23535 33915
rect 23477 33875 23535 33881
rect 24210 33872 24216 33924
rect 24268 33912 24274 33924
rect 24504 33921 24532 34088
rect 24946 34008 24952 34060
rect 25004 34048 25010 34060
rect 25004 34020 25347 34048
rect 25004 34008 25010 34020
rect 24578 33940 24584 33992
rect 24636 33980 24642 33992
rect 25041 33983 25099 33989
rect 25041 33980 25053 33983
rect 24636 33952 25053 33980
rect 24636 33940 24642 33952
rect 25041 33949 25053 33952
rect 25087 33949 25099 33983
rect 25201 33980 25207 33992
rect 25162 33952 25207 33980
rect 25041 33943 25099 33949
rect 25201 33940 25207 33952
rect 25259 33940 25265 33992
rect 25319 33989 25347 34020
rect 25304 33983 25362 33989
rect 25304 33949 25316 33983
rect 25350 33949 25362 33983
rect 25304 33943 25362 33949
rect 25455 33983 25513 33989
rect 25455 33949 25467 33983
rect 25501 33980 25513 33983
rect 25608 33980 25636 34088
rect 27522 34048 27528 34060
rect 27483 34020 27528 34048
rect 27522 34008 27528 34020
rect 27580 34008 27586 34060
rect 30282 34048 30288 34060
rect 30243 34020 30288 34048
rect 30282 34008 30288 34020
rect 30340 34008 30346 34060
rect 35360 34048 35388 34144
rect 35360 34020 36308 34048
rect 35894 33980 35900 33992
rect 25501 33952 25636 33980
rect 35855 33952 35900 33980
rect 25501 33949 25513 33952
rect 25455 33943 25513 33949
rect 35894 33940 35900 33952
rect 35952 33940 35958 33992
rect 36078 33980 36084 33992
rect 36039 33952 36084 33980
rect 36078 33940 36084 33952
rect 36136 33940 36142 33992
rect 36280 33989 36308 34020
rect 36173 33983 36231 33989
rect 36173 33949 36185 33983
rect 36219 33949 36231 33983
rect 36173 33943 36231 33949
rect 36265 33983 36323 33989
rect 36265 33949 36277 33983
rect 36311 33949 36323 33983
rect 36265 33943 36323 33949
rect 24489 33915 24547 33921
rect 24489 33912 24501 33915
rect 24268 33884 24501 33912
rect 24268 33872 24274 33884
rect 24489 33881 24501 33884
rect 24535 33881 24547 33915
rect 24489 33875 24547 33881
rect 25685 33915 25743 33921
rect 25685 33881 25697 33915
rect 25731 33912 25743 33915
rect 27258 33915 27316 33921
rect 27258 33912 27270 33915
rect 25731 33884 27270 33912
rect 25731 33881 25743 33884
rect 25685 33875 25743 33881
rect 27258 33881 27270 33884
rect 27304 33881 27316 33915
rect 27258 33875 27316 33881
rect 29638 33872 29644 33924
rect 29696 33912 29702 33924
rect 30530 33915 30588 33921
rect 30530 33912 30542 33915
rect 29696 33884 30542 33912
rect 29696 33872 29702 33884
rect 30530 33881 30542 33884
rect 30576 33881 30588 33915
rect 30530 33875 30588 33881
rect 31110 33872 31116 33924
rect 31168 33912 31174 33924
rect 32125 33915 32183 33921
rect 32125 33912 32137 33915
rect 31168 33884 32137 33912
rect 31168 33872 31174 33884
rect 32125 33881 32137 33884
rect 32171 33881 32183 33915
rect 32125 33875 32183 33881
rect 32309 33915 32367 33921
rect 32309 33881 32321 33915
rect 32355 33881 32367 33915
rect 36188 33912 36216 33943
rect 36446 33912 36452 33924
rect 36188 33884 36452 33912
rect 32309 33875 32367 33881
rect 19337 33847 19395 33853
rect 19337 33813 19349 33847
rect 19383 33813 19395 33847
rect 19337 33807 19395 33813
rect 22189 33847 22247 33853
rect 22189 33813 22201 33847
rect 22235 33844 22247 33847
rect 22370 33844 22376 33856
rect 22235 33816 22376 33844
rect 22235 33813 22247 33816
rect 22189 33807 22247 33813
rect 22370 33804 22376 33816
rect 22428 33804 22434 33856
rect 22738 33844 22744 33856
rect 22699 33816 22744 33844
rect 22738 33804 22744 33816
rect 22796 33804 22802 33856
rect 23198 33844 23204 33856
rect 23159 33816 23204 33844
rect 23198 33804 23204 33816
rect 23256 33804 23262 33856
rect 23566 33804 23572 33856
rect 23624 33844 23630 33856
rect 24854 33844 24860 33856
rect 23624 33816 24860 33844
rect 23624 33804 23630 33816
rect 24854 33804 24860 33816
rect 24912 33804 24918 33856
rect 25038 33804 25044 33856
rect 25096 33844 25102 33856
rect 26145 33847 26203 33853
rect 26145 33844 26157 33847
rect 25096 33816 26157 33844
rect 25096 33804 25102 33816
rect 26145 33813 26157 33816
rect 26191 33813 26203 33847
rect 26145 33807 26203 33813
rect 31478 33804 31484 33856
rect 31536 33844 31542 33856
rect 31665 33847 31723 33853
rect 31665 33844 31677 33847
rect 31536 33816 31677 33844
rect 31536 33804 31542 33816
rect 31665 33813 31677 33816
rect 31711 33844 31723 33847
rect 32324 33844 32352 33875
rect 36446 33872 36452 33884
rect 36504 33872 36510 33924
rect 32490 33844 32496 33856
rect 31711 33816 32352 33844
rect 32451 33816 32496 33844
rect 31711 33813 31723 33816
rect 31665 33807 31723 33813
rect 32490 33804 32496 33816
rect 32548 33804 32554 33856
rect 33410 33844 33416 33856
rect 33371 33816 33416 33844
rect 33410 33804 33416 33816
rect 33468 33804 33474 33856
rect 36541 33847 36599 33853
rect 36541 33813 36553 33847
rect 36587 33844 36599 33847
rect 38194 33844 38200 33856
rect 36587 33816 38200 33844
rect 36587 33813 36599 33816
rect 36541 33807 36599 33813
rect 38194 33804 38200 33816
rect 38252 33804 38258 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 4246 33600 4252 33652
rect 4304 33640 4310 33652
rect 4801 33643 4859 33649
rect 4801 33640 4813 33643
rect 4304 33612 4813 33640
rect 4304 33600 4310 33612
rect 4801 33609 4813 33612
rect 4847 33609 4859 33643
rect 4801 33603 4859 33609
rect 4890 33600 4896 33652
rect 4948 33640 4954 33652
rect 6638 33640 6644 33652
rect 4948 33612 6644 33640
rect 4948 33600 4954 33612
rect 6638 33600 6644 33612
rect 6696 33640 6702 33652
rect 8294 33640 8300 33652
rect 6696 33612 8064 33640
rect 8255 33612 8300 33640
rect 6696 33600 6702 33612
rect 8036 33584 8064 33612
rect 8294 33600 8300 33612
rect 8352 33600 8358 33652
rect 9309 33643 9367 33649
rect 9309 33609 9321 33643
rect 9355 33640 9367 33643
rect 10318 33640 10324 33652
rect 9355 33612 10324 33640
rect 9355 33609 9367 33612
rect 9309 33603 9367 33609
rect 10318 33600 10324 33612
rect 10376 33600 10382 33652
rect 14185 33643 14243 33649
rect 14185 33609 14197 33643
rect 14231 33640 14243 33643
rect 14826 33640 14832 33652
rect 14231 33612 14832 33640
rect 14231 33609 14243 33612
rect 14185 33603 14243 33609
rect 14826 33600 14832 33612
rect 14884 33600 14890 33652
rect 19334 33600 19340 33652
rect 19392 33600 19398 33652
rect 19705 33643 19763 33649
rect 19705 33609 19717 33643
rect 19751 33640 19763 33643
rect 19978 33640 19984 33652
rect 19751 33612 19984 33640
rect 19751 33609 19763 33612
rect 19705 33603 19763 33609
rect 19978 33600 19984 33612
rect 20036 33600 20042 33652
rect 24029 33643 24087 33649
rect 24029 33609 24041 33643
rect 24075 33640 24087 33643
rect 24118 33640 24124 33652
rect 24075 33612 24124 33640
rect 24075 33609 24087 33612
rect 24029 33603 24087 33609
rect 24118 33600 24124 33612
rect 24176 33600 24182 33652
rect 24394 33600 24400 33652
rect 24452 33640 24458 33652
rect 24762 33640 24768 33652
rect 24452 33612 24768 33640
rect 24452 33600 24458 33612
rect 24762 33600 24768 33612
rect 24820 33640 24826 33652
rect 24946 33640 24952 33652
rect 24820 33612 24952 33640
rect 24820 33600 24826 33612
rect 24946 33600 24952 33612
rect 25004 33600 25010 33652
rect 29086 33640 29092 33652
rect 29047 33612 29092 33640
rect 29086 33600 29092 33612
rect 29144 33600 29150 33652
rect 29638 33640 29644 33652
rect 29599 33612 29644 33640
rect 29638 33600 29644 33612
rect 29696 33600 29702 33652
rect 29730 33600 29736 33652
rect 29788 33640 29794 33652
rect 30975 33643 31033 33649
rect 30975 33640 30987 33643
rect 29788 33612 30987 33640
rect 29788 33600 29794 33612
rect 4157 33575 4215 33581
rect 4157 33541 4169 33575
rect 4203 33572 4215 33575
rect 4706 33572 4712 33584
rect 4203 33544 4712 33572
rect 4203 33541 4215 33544
rect 4157 33535 4215 33541
rect 4706 33532 4712 33544
rect 4764 33532 4770 33584
rect 4982 33572 4988 33584
rect 4943 33544 4988 33572
rect 4982 33532 4988 33544
rect 5040 33532 5046 33584
rect 5169 33575 5227 33581
rect 5169 33541 5181 33575
rect 5215 33572 5227 33575
rect 6730 33572 6736 33584
rect 5215 33544 6736 33572
rect 5215 33541 5227 33544
rect 5169 33535 5227 33541
rect 4341 33507 4399 33513
rect 4341 33473 4353 33507
rect 4387 33504 4399 33507
rect 5184 33504 5212 33535
rect 6730 33532 6736 33544
rect 6788 33532 6794 33584
rect 8018 33532 8024 33584
rect 8076 33572 8082 33584
rect 9769 33575 9827 33581
rect 9769 33572 9781 33575
rect 8076 33544 9781 33572
rect 8076 33532 8082 33544
rect 9769 33541 9781 33544
rect 9815 33541 9827 33575
rect 9769 33535 9827 33541
rect 10134 33532 10140 33584
rect 10192 33572 10198 33584
rect 15194 33572 15200 33584
rect 10192 33544 15200 33572
rect 10192 33532 10198 33544
rect 15194 33532 15200 33544
rect 15252 33572 15258 33584
rect 15289 33575 15347 33581
rect 15289 33572 15301 33575
rect 15252 33544 15301 33572
rect 15252 33532 15258 33544
rect 15289 33541 15301 33544
rect 15335 33541 15347 33575
rect 15289 33535 15347 33541
rect 15473 33575 15531 33581
rect 15473 33541 15485 33575
rect 15519 33572 15531 33575
rect 16942 33572 16948 33584
rect 15519 33544 16948 33572
rect 15519 33541 15531 33544
rect 15473 33535 15531 33541
rect 16942 33532 16948 33544
rect 17000 33572 17006 33584
rect 17770 33572 17776 33584
rect 17000 33544 17776 33572
rect 17000 33532 17006 33544
rect 17770 33532 17776 33544
rect 17828 33532 17834 33584
rect 19352 33572 19380 33600
rect 19260 33544 19380 33572
rect 9122 33504 9128 33516
rect 4387 33476 5212 33504
rect 9083 33476 9128 33504
rect 4387 33473 4399 33476
rect 4341 33467 4399 33473
rect 9122 33464 9128 33476
rect 9180 33464 9186 33516
rect 9953 33507 10011 33513
rect 9953 33473 9965 33507
rect 9999 33473 10011 33507
rect 10594 33504 10600 33516
rect 10555 33476 10600 33504
rect 9953 33467 10011 33473
rect 4982 33436 4988 33448
rect 4908 33408 4988 33436
rect 4908 33312 4936 33408
rect 4982 33396 4988 33408
rect 5040 33396 5046 33448
rect 9968 33436 9996 33467
rect 10594 33464 10600 33476
rect 10652 33464 10658 33516
rect 14001 33507 14059 33513
rect 14001 33473 14013 33507
rect 14047 33504 14059 33507
rect 15010 33504 15016 33516
rect 14047 33476 15016 33504
rect 14047 33473 14059 33476
rect 14001 33467 14059 33473
rect 15010 33464 15016 33476
rect 15068 33464 15074 33516
rect 19058 33504 19064 33516
rect 19019 33476 19064 33504
rect 19058 33464 19064 33476
rect 19116 33464 19122 33516
rect 19260 33513 19288 33544
rect 23014 33532 23020 33584
rect 23072 33572 23078 33584
rect 23385 33575 23443 33581
rect 23385 33572 23397 33575
rect 23072 33544 23397 33572
rect 23072 33532 23078 33544
rect 23385 33541 23397 33544
rect 23431 33541 23443 33575
rect 23566 33572 23572 33584
rect 23527 33544 23572 33572
rect 23385 33535 23443 33541
rect 23566 33532 23572 33544
rect 23624 33532 23630 33584
rect 23934 33532 23940 33584
rect 23992 33572 23998 33584
rect 23992 33544 24302 33572
rect 23992 33532 23998 33544
rect 19245 33507 19303 33513
rect 19245 33473 19257 33507
rect 19291 33473 19303 33507
rect 19245 33467 19303 33473
rect 19337 33507 19395 33513
rect 19337 33473 19349 33507
rect 19383 33473 19395 33507
rect 19337 33467 19395 33473
rect 19429 33507 19487 33513
rect 19429 33473 19441 33507
rect 19475 33504 19487 33507
rect 20254 33504 20260 33516
rect 19475 33476 20260 33504
rect 19475 33473 19487 33476
rect 19429 33467 19487 33473
rect 17126 33436 17132 33448
rect 9968 33408 17132 33436
rect 17126 33396 17132 33408
rect 17184 33436 17190 33448
rect 17589 33439 17647 33445
rect 17589 33436 17601 33439
rect 17184 33408 17601 33436
rect 17184 33396 17190 33408
rect 17589 33405 17601 33408
rect 17635 33405 17647 33439
rect 17589 33399 17647 33405
rect 17865 33439 17923 33445
rect 17865 33405 17877 33439
rect 17911 33436 17923 33439
rect 19352 33436 19380 33467
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 21913 33507 21971 33513
rect 21913 33473 21925 33507
rect 21959 33504 21971 33507
rect 22649 33507 22707 33513
rect 22649 33504 22661 33507
rect 21959 33476 22661 33504
rect 21959 33473 21971 33476
rect 21913 33467 21971 33473
rect 22649 33473 22661 33476
rect 22695 33504 22707 33507
rect 22922 33504 22928 33516
rect 22695 33476 22928 33504
rect 22695 33473 22707 33476
rect 22649 33467 22707 33473
rect 22922 33464 22928 33476
rect 22980 33464 22986 33516
rect 24274 33513 24302 33544
rect 24578 33532 24584 33584
rect 24636 33572 24642 33584
rect 24636 33544 24808 33572
rect 24636 33532 24642 33544
rect 24259 33507 24317 33513
rect 24259 33473 24271 33507
rect 24305 33473 24317 33507
rect 24259 33467 24317 33473
rect 24381 33467 24387 33519
rect 24439 33513 24445 33519
rect 24439 33507 24455 33513
rect 24443 33473 24455 33507
rect 24439 33467 24455 33473
rect 24489 33507 24547 33513
rect 24489 33473 24501 33507
rect 24535 33504 24547 33507
rect 24685 33507 24743 33513
rect 24535 33476 24624 33504
rect 24535 33473 24547 33476
rect 24489 33467 24547 33473
rect 20070 33436 20076 33448
rect 17911 33408 20076 33436
rect 17911 33405 17923 33408
rect 17865 33399 17923 33405
rect 20070 33396 20076 33408
rect 20128 33396 20134 33448
rect 6178 33328 6184 33380
rect 6236 33368 6242 33380
rect 10686 33368 10692 33380
rect 6236 33340 10692 33368
rect 6236 33328 6242 33340
rect 10686 33328 10692 33340
rect 10744 33368 10750 33380
rect 20272 33377 20300 33464
rect 23201 33439 23259 33445
rect 23201 33405 23213 33439
rect 23247 33436 23259 33439
rect 24596 33436 24624 33476
rect 24685 33473 24697 33507
rect 24731 33504 24743 33507
rect 24780 33504 24808 33544
rect 25130 33504 25136 33516
rect 24731 33476 24808 33504
rect 25091 33476 25136 33504
rect 24731 33473 24743 33476
rect 24685 33467 24743 33473
rect 25130 33464 25136 33476
rect 25188 33464 25194 33516
rect 29104 33504 29132 33600
rect 30024 33513 30052 33612
rect 30975 33609 30987 33612
rect 31021 33609 31033 33643
rect 30975 33603 31033 33609
rect 31202 33600 31208 33652
rect 31260 33640 31266 33652
rect 33410 33640 33416 33652
rect 31260 33612 33416 33640
rect 31260 33600 31266 33612
rect 33410 33600 33416 33612
rect 33468 33640 33474 33652
rect 35253 33643 35311 33649
rect 35253 33640 35265 33643
rect 33468 33612 35265 33640
rect 33468 33600 33474 33612
rect 35253 33609 35265 33612
rect 35299 33640 35311 33643
rect 35299 33612 36124 33640
rect 35299 33609 35311 33612
rect 35253 33603 35311 33609
rect 32490 33572 32496 33584
rect 30116 33544 32496 33572
rect 30116 33513 30144 33544
rect 32490 33532 32496 33544
rect 32548 33532 32554 33584
rect 35894 33572 35900 33584
rect 35820 33544 35900 33572
rect 29917 33507 29975 33513
rect 29917 33504 29929 33507
rect 29104 33476 29929 33504
rect 29917 33473 29929 33476
rect 29963 33473 29975 33507
rect 29917 33467 29975 33473
rect 30009 33507 30067 33513
rect 30009 33473 30021 33507
rect 30055 33473 30067 33507
rect 30009 33467 30067 33473
rect 30101 33507 30159 33513
rect 30101 33473 30113 33507
rect 30147 33473 30159 33507
rect 30101 33467 30159 33473
rect 30285 33507 30343 33513
rect 30285 33473 30297 33507
rect 30331 33504 30343 33507
rect 30558 33504 30564 33516
rect 30331 33476 30564 33504
rect 30331 33473 30343 33476
rect 30285 33467 30343 33473
rect 30558 33464 30564 33476
rect 30616 33504 30622 33516
rect 35820 33513 35848 33544
rect 35894 33532 35900 33544
rect 35952 33532 35958 33584
rect 36096 33572 36124 33612
rect 36449 33575 36507 33581
rect 36096 33544 36216 33572
rect 35805 33507 35863 33513
rect 35805 33504 35817 33507
rect 30616 33476 35817 33504
rect 30616 33464 30622 33476
rect 35805 33473 35817 33476
rect 35851 33473 35863 33507
rect 35986 33504 35992 33516
rect 35947 33476 35992 33504
rect 35805 33467 35863 33473
rect 35986 33464 35992 33476
rect 36044 33464 36050 33516
rect 36188 33513 36216 33544
rect 36449 33541 36461 33575
rect 36495 33572 36507 33575
rect 38390 33575 38448 33581
rect 38390 33572 38402 33575
rect 36495 33544 38402 33572
rect 36495 33541 36507 33544
rect 36449 33535 36507 33541
rect 38390 33541 38402 33544
rect 38436 33541 38448 33575
rect 38390 33535 38448 33541
rect 36081 33507 36139 33513
rect 36081 33473 36093 33507
rect 36127 33473 36139 33507
rect 36081 33467 36139 33473
rect 36173 33507 36231 33513
rect 36173 33473 36185 33507
rect 36219 33473 36231 33507
rect 36173 33467 36231 33473
rect 23247 33408 24624 33436
rect 30745 33439 30803 33445
rect 23247 33405 23259 33408
rect 23201 33399 23259 33405
rect 30745 33405 30757 33439
rect 30791 33405 30803 33439
rect 36096 33436 36124 33467
rect 38562 33464 38568 33516
rect 38620 33504 38626 33516
rect 38657 33507 38715 33513
rect 38657 33504 38669 33507
rect 38620 33476 38669 33504
rect 38620 33464 38626 33476
rect 38657 33473 38669 33476
rect 38703 33473 38715 33507
rect 38657 33467 38715 33473
rect 36446 33436 36452 33448
rect 36096 33408 36452 33436
rect 30745 33399 30803 33405
rect 10781 33371 10839 33377
rect 10781 33368 10793 33371
rect 10744 33340 10793 33368
rect 10744 33328 10750 33340
rect 10781 33337 10793 33340
rect 10827 33337 10839 33371
rect 10781 33331 10839 33337
rect 20257 33371 20315 33377
rect 20257 33337 20269 33371
rect 20303 33368 20315 33371
rect 25222 33368 25228 33380
rect 20303 33340 25228 33368
rect 20303 33337 20315 33340
rect 20257 33331 20315 33337
rect 25222 33328 25228 33340
rect 25280 33328 25286 33380
rect 30760 33368 30788 33399
rect 36446 33396 36452 33408
rect 36504 33396 36510 33448
rect 31846 33368 31852 33380
rect 30760 33340 31852 33368
rect 31846 33328 31852 33340
rect 31904 33328 31910 33380
rect 58158 33368 58164 33380
rect 58119 33340 58164 33368
rect 58158 33328 58164 33340
rect 58216 33328 58222 33380
rect 3973 33303 4031 33309
rect 3973 33269 3985 33303
rect 4019 33300 4031 33303
rect 4614 33300 4620 33312
rect 4019 33272 4620 33300
rect 4019 33269 4031 33272
rect 3973 33263 4031 33269
rect 4614 33260 4620 33272
rect 4672 33260 4678 33312
rect 4890 33260 4896 33312
rect 4948 33260 4954 33312
rect 22465 33303 22523 33309
rect 22465 33269 22477 33303
rect 22511 33300 22523 33303
rect 24486 33300 24492 33312
rect 22511 33272 24492 33300
rect 22511 33269 22523 33272
rect 22465 33263 22523 33269
rect 24486 33260 24492 33272
rect 24544 33260 24550 33312
rect 25130 33260 25136 33312
rect 25188 33300 25194 33312
rect 31202 33300 31208 33312
rect 25188 33272 31208 33300
rect 25188 33260 25194 33272
rect 31202 33260 31208 33272
rect 31260 33260 31266 33312
rect 37274 33300 37280 33312
rect 37235 33272 37280 33300
rect 37274 33260 37280 33272
rect 37332 33260 37338 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 6730 33056 6736 33108
rect 6788 33096 6794 33108
rect 7193 33099 7251 33105
rect 7193 33096 7205 33099
rect 6788 33068 7205 33096
rect 6788 33056 6794 33068
rect 7193 33065 7205 33068
rect 7239 33065 7251 33099
rect 7193 33059 7251 33065
rect 7466 33056 7472 33108
rect 7524 33096 7530 33108
rect 9030 33096 9036 33108
rect 7524 33068 9036 33096
rect 7524 33056 7530 33068
rect 9030 33056 9036 33068
rect 9088 33096 9094 33108
rect 17402 33096 17408 33108
rect 9088 33068 17408 33096
rect 9088 33056 9094 33068
rect 17402 33056 17408 33068
rect 17460 33056 17466 33108
rect 17773 33099 17831 33105
rect 17773 33065 17785 33099
rect 17819 33096 17831 33099
rect 19150 33096 19156 33108
rect 17819 33068 19156 33096
rect 17819 33065 17831 33068
rect 17773 33059 17831 33065
rect 19150 33056 19156 33068
rect 19208 33056 19214 33108
rect 20346 33096 20352 33108
rect 19444 33068 20352 33096
rect 4798 33028 4804 33040
rect 4172 33000 4804 33028
rect 4172 32901 4200 33000
rect 4798 32988 4804 33000
rect 4856 32988 4862 33040
rect 7650 32988 7656 33040
rect 7708 33028 7714 33040
rect 8113 33031 8171 33037
rect 8113 33028 8125 33031
rect 7708 33000 8125 33028
rect 7708 32988 7714 33000
rect 8113 32997 8125 33000
rect 8159 32997 8171 33031
rect 8113 32991 8171 32997
rect 11992 33000 12940 33028
rect 4614 32960 4620 32972
rect 4264 32932 4620 32960
rect 4264 32901 4292 32932
rect 4614 32920 4620 32932
rect 4672 32920 4678 32972
rect 4985 32963 5043 32969
rect 4985 32929 4997 32963
rect 5031 32960 5043 32963
rect 5074 32960 5080 32972
rect 5031 32932 5080 32960
rect 5031 32929 5043 32932
rect 4985 32923 5043 32929
rect 4065 32895 4123 32901
rect 4065 32861 4077 32895
rect 4111 32861 4123 32895
rect 4065 32855 4123 32861
rect 4157 32895 4215 32901
rect 4157 32861 4169 32895
rect 4203 32861 4215 32895
rect 4157 32855 4215 32861
rect 4249 32895 4307 32901
rect 4249 32861 4261 32895
rect 4295 32861 4307 32895
rect 4249 32855 4307 32861
rect 4433 32895 4491 32901
rect 4433 32861 4445 32895
rect 4479 32892 4491 32895
rect 5000 32892 5028 32923
rect 5074 32920 5080 32932
rect 5132 32960 5138 32972
rect 7006 32960 7012 32972
rect 5132 32932 7012 32960
rect 5132 32920 5138 32932
rect 7006 32920 7012 32932
rect 7064 32920 7070 32972
rect 9585 32963 9643 32969
rect 9585 32929 9597 32963
rect 9631 32960 9643 32963
rect 10042 32960 10048 32972
rect 9631 32932 10048 32960
rect 9631 32929 9643 32932
rect 9585 32923 9643 32929
rect 4479 32864 5028 32892
rect 6365 32895 6423 32901
rect 4479 32861 4491 32864
rect 4433 32855 4491 32861
rect 6365 32861 6377 32895
rect 6411 32892 6423 32895
rect 6730 32892 6736 32904
rect 6411 32864 6736 32892
rect 6411 32861 6423 32864
rect 6365 32855 6423 32861
rect 4080 32824 4108 32855
rect 6730 32852 6736 32864
rect 6788 32852 6794 32904
rect 7374 32892 7380 32904
rect 7335 32864 7380 32892
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 8297 32895 8355 32901
rect 8297 32861 8309 32895
rect 8343 32892 8355 32895
rect 9600 32892 9628 32923
rect 10042 32920 10048 32932
rect 10100 32920 10106 32972
rect 9858 32892 9864 32904
rect 8343 32864 9628 32892
rect 9819 32864 9864 32892
rect 8343 32861 8355 32864
rect 8297 32855 8355 32861
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 9950 32852 9956 32904
rect 10008 32892 10014 32904
rect 11701 32895 11759 32901
rect 11701 32892 11713 32895
rect 10008 32864 11713 32892
rect 10008 32852 10014 32864
rect 11701 32861 11713 32864
rect 11747 32861 11759 32895
rect 11701 32855 11759 32861
rect 11992 32836 12020 33000
rect 12802 32960 12808 32972
rect 12406 32932 12808 32960
rect 12069 32895 12127 32901
rect 12069 32861 12081 32895
rect 12115 32892 12127 32895
rect 12406 32892 12434 32932
rect 12802 32920 12808 32932
rect 12860 32920 12866 32972
rect 12912 32901 12940 33000
rect 16850 32988 16856 33040
rect 16908 33028 16914 33040
rect 19444 33028 19472 33068
rect 20346 33056 20352 33068
rect 20404 33096 20410 33108
rect 22002 33096 22008 33108
rect 20404 33068 22008 33096
rect 20404 33056 20410 33068
rect 22002 33056 22008 33068
rect 22060 33096 22066 33108
rect 22557 33099 22615 33105
rect 22557 33096 22569 33099
rect 22060 33068 22569 33096
rect 22060 33056 22066 33068
rect 22557 33065 22569 33068
rect 22603 33065 22615 33099
rect 22557 33059 22615 33065
rect 23658 33056 23664 33108
rect 23716 33096 23722 33108
rect 23753 33099 23811 33105
rect 23753 33096 23765 33099
rect 23716 33068 23765 33096
rect 23716 33056 23722 33068
rect 23753 33065 23765 33068
rect 23799 33065 23811 33099
rect 23753 33059 23811 33065
rect 16908 33000 19472 33028
rect 16908 32988 16914 33000
rect 23768 32960 23796 33059
rect 23934 33056 23940 33108
rect 23992 33096 23998 33108
rect 25130 33096 25136 33108
rect 23992 33068 25136 33096
rect 23992 33056 23998 33068
rect 25130 33056 25136 33068
rect 25188 33056 25194 33108
rect 27338 33056 27344 33108
rect 27396 33096 27402 33108
rect 29641 33099 29699 33105
rect 29641 33096 29653 33099
rect 27396 33068 29653 33096
rect 27396 33056 27402 33068
rect 29641 33065 29653 33068
rect 29687 33096 29699 33099
rect 32030 33096 32036 33108
rect 29687 33068 32036 33096
rect 29687 33065 29699 33068
rect 29641 33059 29699 33065
rect 32030 33056 32036 33068
rect 32088 33056 32094 33108
rect 35437 33099 35495 33105
rect 35437 33065 35449 33099
rect 35483 33096 35495 33099
rect 35986 33096 35992 33108
rect 35483 33068 35992 33096
rect 35483 33065 35495 33068
rect 35437 33059 35495 33065
rect 35986 33056 35992 33068
rect 36044 33056 36050 33108
rect 31110 33028 31116 33040
rect 31071 33000 31116 33028
rect 31110 32988 31116 33000
rect 31168 32988 31174 33040
rect 35342 33028 35348 33040
rect 34808 33000 35348 33028
rect 34808 32972 34836 33000
rect 35342 32988 35348 33000
rect 35400 32988 35406 33040
rect 35802 32988 35808 33040
rect 35860 33028 35866 33040
rect 37093 33031 37151 33037
rect 37093 33028 37105 33031
rect 35860 33000 37105 33028
rect 35860 32988 35866 33000
rect 37093 32997 37105 33000
rect 37139 32997 37151 33031
rect 37093 32991 37151 32997
rect 24397 32963 24455 32969
rect 24397 32960 24409 32963
rect 23768 32932 24409 32960
rect 24397 32929 24409 32932
rect 24443 32929 24455 32963
rect 24397 32923 24455 32929
rect 25222 32920 25228 32972
rect 25280 32960 25286 32972
rect 34790 32960 34796 32972
rect 25280 32932 34796 32960
rect 25280 32920 25286 32932
rect 34790 32920 34796 32932
rect 34848 32920 34854 32972
rect 37274 32960 37280 32972
rect 35268 32932 37280 32960
rect 12115 32864 12434 32892
rect 12897 32895 12955 32901
rect 12115 32861 12127 32864
rect 12069 32855 12127 32861
rect 12897 32861 12909 32895
rect 12943 32861 12955 32895
rect 12897 32855 12955 32861
rect 12986 32852 12992 32904
rect 13044 32892 13050 32904
rect 14093 32895 14151 32901
rect 14093 32892 14105 32895
rect 13044 32864 14105 32892
rect 13044 32852 13050 32864
rect 14093 32861 14105 32864
rect 14139 32892 14151 32895
rect 16114 32892 16120 32904
rect 14139 32864 16120 32892
rect 14139 32861 14151 32864
rect 14093 32855 14151 32861
rect 16114 32852 16120 32864
rect 16172 32852 16178 32904
rect 17586 32892 17592 32904
rect 17547 32864 17592 32892
rect 17586 32852 17592 32864
rect 17644 32852 17650 32904
rect 20806 32852 20812 32904
rect 20864 32892 20870 32904
rect 21637 32895 21695 32901
rect 21637 32892 21649 32895
rect 20864 32864 21649 32892
rect 20864 32852 20870 32864
rect 21637 32861 21649 32864
rect 21683 32861 21695 32895
rect 21637 32855 21695 32861
rect 24486 32852 24492 32904
rect 24544 32892 24550 32904
rect 24673 32895 24731 32901
rect 24673 32892 24685 32895
rect 24544 32864 24685 32892
rect 24544 32852 24550 32864
rect 24673 32861 24685 32864
rect 24719 32861 24731 32895
rect 24673 32855 24731 32861
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32892 28871 32895
rect 30466 32892 30472 32904
rect 28859 32864 30472 32892
rect 28859 32861 28871 32864
rect 28813 32855 28871 32861
rect 30466 32852 30472 32864
rect 30524 32852 30530 32904
rect 30558 32852 30564 32904
rect 30616 32892 30622 32904
rect 30929 32895 30987 32901
rect 30929 32892 30941 32895
rect 30616 32864 30941 32892
rect 30616 32852 30622 32864
rect 30929 32861 30941 32864
rect 30975 32861 30987 32895
rect 30929 32855 30987 32861
rect 32582 32852 32588 32904
rect 32640 32892 32646 32904
rect 32677 32895 32735 32901
rect 32677 32892 32689 32895
rect 32640 32864 32689 32892
rect 32640 32852 32646 32864
rect 32677 32861 32689 32864
rect 32723 32861 32735 32895
rect 33042 32892 33048 32904
rect 33003 32864 33048 32892
rect 32677 32855 32735 32861
rect 33042 32852 33048 32864
rect 33100 32852 33106 32904
rect 33134 32852 33140 32904
rect 33192 32892 33198 32904
rect 35268 32901 35296 32932
rect 37274 32920 37280 32932
rect 37332 32920 37338 32972
rect 38473 32963 38531 32969
rect 38473 32929 38485 32963
rect 38519 32960 38531 32963
rect 38562 32960 38568 32972
rect 38519 32932 38568 32960
rect 38519 32929 38531 32932
rect 38473 32923 38531 32929
rect 38562 32920 38568 32932
rect 38620 32920 38626 32972
rect 35253 32895 35311 32901
rect 35253 32892 35265 32895
rect 33192 32864 35265 32892
rect 33192 32852 33198 32864
rect 35253 32861 35265 32864
rect 35299 32861 35311 32895
rect 35253 32855 35311 32861
rect 35894 32852 35900 32904
rect 35952 32892 35958 32904
rect 36078 32892 36084 32904
rect 35952 32864 35997 32892
rect 36039 32864 36084 32892
rect 35952 32852 35958 32864
rect 36078 32852 36084 32864
rect 36136 32852 36142 32904
rect 36173 32895 36231 32901
rect 36173 32861 36185 32895
rect 36219 32861 36231 32895
rect 36173 32855 36231 32861
rect 5166 32824 5172 32836
rect 4080 32796 5172 32824
rect 5166 32784 5172 32796
rect 5224 32784 5230 32836
rect 6549 32827 6607 32833
rect 6549 32793 6561 32827
rect 6595 32824 6607 32827
rect 7098 32824 7104 32836
rect 6595 32796 7104 32824
rect 6595 32793 6607 32796
rect 6549 32787 6607 32793
rect 7098 32784 7104 32796
rect 7156 32784 7162 32836
rect 11885 32827 11943 32833
rect 11885 32793 11897 32827
rect 11931 32793 11943 32827
rect 11885 32787 11943 32793
rect 3786 32756 3792 32768
rect 3747 32728 3792 32756
rect 3786 32716 3792 32728
rect 3844 32716 3850 32768
rect 6733 32759 6791 32765
rect 6733 32725 6745 32759
rect 6779 32756 6791 32759
rect 6914 32756 6920 32768
rect 6779 32728 6920 32756
rect 6779 32725 6791 32728
rect 6733 32719 6791 32725
rect 6914 32716 6920 32728
rect 6972 32716 6978 32768
rect 11900 32756 11928 32787
rect 11974 32784 11980 32836
rect 12032 32824 12038 32836
rect 12526 32824 12532 32836
rect 12032 32796 12077 32824
rect 12176 32796 12532 32824
rect 12032 32784 12038 32796
rect 12176 32756 12204 32796
rect 12526 32784 12532 32796
rect 12584 32784 12590 32836
rect 12618 32784 12624 32836
rect 12676 32824 12682 32836
rect 12713 32827 12771 32833
rect 12713 32824 12725 32827
rect 12676 32796 12725 32824
rect 12676 32784 12682 32796
rect 12713 32793 12725 32796
rect 12759 32793 12771 32827
rect 14360 32827 14418 32833
rect 12713 32787 12771 32793
rect 12912 32796 13216 32824
rect 11900 32728 12204 32756
rect 12253 32759 12311 32765
rect 12253 32725 12265 32759
rect 12299 32756 12311 32759
rect 12912 32756 12940 32796
rect 13078 32756 13084 32768
rect 12299 32728 12940 32756
rect 13039 32728 13084 32756
rect 12299 32725 12311 32728
rect 12253 32719 12311 32725
rect 13078 32716 13084 32728
rect 13136 32716 13142 32768
rect 13188 32756 13216 32796
rect 14360 32793 14372 32827
rect 14406 32824 14418 32827
rect 14550 32824 14556 32836
rect 14406 32796 14556 32824
rect 14406 32793 14418 32796
rect 14360 32787 14418 32793
rect 14550 32784 14556 32796
rect 14608 32784 14614 32836
rect 21392 32827 21450 32833
rect 21392 32793 21404 32827
rect 21438 32824 21450 32827
rect 21818 32824 21824 32836
rect 21438 32796 21824 32824
rect 21438 32793 21450 32796
rect 21392 32787 21450 32793
rect 21818 32784 21824 32796
rect 21876 32784 21882 32836
rect 28534 32784 28540 32836
rect 28592 32824 28598 32836
rect 28629 32827 28687 32833
rect 28629 32824 28641 32827
rect 28592 32796 28641 32824
rect 28592 32784 28598 32796
rect 28629 32793 28641 32796
rect 28675 32793 28687 32827
rect 28629 32787 28687 32793
rect 32769 32827 32827 32833
rect 32769 32793 32781 32827
rect 32815 32793 32827 32827
rect 32769 32787 32827 32793
rect 15102 32756 15108 32768
rect 13188 32728 15108 32756
rect 15102 32716 15108 32728
rect 15160 32716 15166 32768
rect 15470 32756 15476 32768
rect 15431 32728 15476 32756
rect 15470 32716 15476 32728
rect 15528 32716 15534 32768
rect 15562 32716 15568 32768
rect 15620 32756 15626 32768
rect 17770 32756 17776 32768
rect 15620 32728 17776 32756
rect 15620 32716 15626 32728
rect 17770 32716 17776 32728
rect 17828 32716 17834 32768
rect 20257 32759 20315 32765
rect 20257 32725 20269 32759
rect 20303 32756 20315 32759
rect 21082 32756 21088 32768
rect 20303 32728 21088 32756
rect 20303 32725 20315 32728
rect 20257 32719 20315 32725
rect 21082 32716 21088 32728
rect 21140 32716 21146 32768
rect 23566 32716 23572 32768
rect 23624 32756 23630 32768
rect 27706 32756 27712 32768
rect 23624 32728 27712 32756
rect 23624 32716 23630 32728
rect 27706 32716 27712 32728
rect 27764 32716 27770 32768
rect 28445 32759 28503 32765
rect 28445 32725 28457 32759
rect 28491 32756 28503 32759
rect 28718 32756 28724 32768
rect 28491 32728 28724 32756
rect 28491 32725 28503 32728
rect 28445 32719 28503 32725
rect 28718 32716 28724 32728
rect 28776 32716 28782 32768
rect 31662 32716 31668 32768
rect 31720 32756 31726 32768
rect 31938 32756 31944 32768
rect 31720 32728 31944 32756
rect 31720 32716 31726 32728
rect 31938 32716 31944 32728
rect 31996 32716 32002 32768
rect 32122 32716 32128 32768
rect 32180 32756 32186 32768
rect 32493 32759 32551 32765
rect 32493 32756 32505 32759
rect 32180 32728 32505 32756
rect 32180 32716 32186 32728
rect 32493 32725 32505 32728
rect 32539 32725 32551 32759
rect 32784 32756 32812 32787
rect 32858 32784 32864 32836
rect 32916 32824 32922 32836
rect 35066 32824 35072 32836
rect 32916 32796 32961 32824
rect 35027 32796 35072 32824
rect 32916 32784 32922 32796
rect 35066 32784 35072 32796
rect 35124 32784 35130 32836
rect 36188 32824 36216 32855
rect 36262 32852 36268 32904
rect 36320 32892 36326 32904
rect 36320 32864 36365 32892
rect 36320 32852 36326 32864
rect 38194 32852 38200 32904
rect 38252 32901 38258 32904
rect 38252 32892 38264 32901
rect 38252 32864 38297 32892
rect 38252 32855 38264 32864
rect 38252 32852 38258 32855
rect 36446 32824 36452 32836
rect 36188 32796 36452 32824
rect 36446 32784 36452 32796
rect 36504 32784 36510 32836
rect 35802 32756 35808 32768
rect 32784 32728 35808 32756
rect 32493 32719 32551 32725
rect 35802 32716 35808 32728
rect 35860 32716 35866 32768
rect 36538 32756 36544 32768
rect 36499 32728 36544 32756
rect 36538 32716 36544 32728
rect 36596 32716 36602 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 4617 32555 4675 32561
rect 4617 32521 4629 32555
rect 4663 32552 4675 32555
rect 5166 32552 5172 32564
rect 4663 32524 5172 32552
rect 4663 32521 4675 32524
rect 4617 32515 4675 32521
rect 5166 32512 5172 32524
rect 5224 32552 5230 32564
rect 6086 32552 6092 32564
rect 5224 32524 6092 32552
rect 5224 32512 5230 32524
rect 6086 32512 6092 32524
rect 6144 32512 6150 32564
rect 6454 32512 6460 32564
rect 6512 32552 6518 32564
rect 7282 32552 7288 32564
rect 6512 32524 7288 32552
rect 6512 32512 6518 32524
rect 7282 32512 7288 32524
rect 7340 32512 7346 32564
rect 7561 32555 7619 32561
rect 7561 32521 7573 32555
rect 7607 32552 7619 32555
rect 11609 32555 11667 32561
rect 7607 32524 10088 32552
rect 7607 32521 7619 32524
rect 7561 32515 7619 32521
rect 6178 32484 6184 32496
rect 2516 32456 6184 32484
rect 2130 32308 2136 32360
rect 2188 32348 2194 32360
rect 2516 32357 2544 32456
rect 6178 32444 6184 32456
rect 6236 32444 6242 32496
rect 7466 32484 7472 32496
rect 6656 32456 7472 32484
rect 2768 32419 2826 32425
rect 2768 32385 2780 32419
rect 2814 32416 2826 32419
rect 3786 32416 3792 32428
rect 2814 32388 3792 32416
rect 2814 32385 2826 32388
rect 2768 32379 2826 32385
rect 3786 32376 3792 32388
rect 3844 32376 3850 32428
rect 5534 32376 5540 32428
rect 5592 32416 5598 32428
rect 6656 32425 6684 32456
rect 7466 32444 7472 32456
rect 7524 32444 7530 32496
rect 5813 32419 5871 32425
rect 5813 32416 5825 32419
rect 5592 32388 5825 32416
rect 5592 32376 5598 32388
rect 5813 32385 5825 32388
rect 5859 32416 5871 32419
rect 6641 32419 6699 32425
rect 6641 32416 6653 32419
rect 5859 32388 6653 32416
rect 5859 32385 5871 32388
rect 5813 32379 5871 32385
rect 6641 32385 6653 32388
rect 6687 32385 6699 32419
rect 6641 32379 6699 32385
rect 6730 32419 6788 32425
rect 6730 32385 6742 32419
rect 6776 32385 6788 32419
rect 6730 32379 6788 32385
rect 6825 32419 6883 32425
rect 6825 32385 6837 32419
rect 6871 32416 6883 32419
rect 6914 32416 6920 32428
rect 6871 32388 6920 32416
rect 6871 32385 6883 32388
rect 6825 32379 6883 32385
rect 2501 32351 2559 32357
rect 2501 32348 2513 32351
rect 2188 32320 2513 32348
rect 2188 32308 2194 32320
rect 2501 32317 2513 32320
rect 2547 32317 2559 32351
rect 2501 32311 2559 32317
rect 5442 32308 5448 32360
rect 5500 32348 5506 32360
rect 6454 32348 6460 32360
rect 5500 32320 6460 32348
rect 5500 32308 5506 32320
rect 6454 32308 6460 32320
rect 6512 32308 6518 32360
rect 3881 32283 3939 32289
rect 3881 32249 3893 32283
rect 3927 32280 3939 32283
rect 4706 32280 4712 32292
rect 3927 32252 4712 32280
rect 3927 32249 3939 32252
rect 3881 32243 3939 32249
rect 4706 32240 4712 32252
rect 4764 32280 4770 32292
rect 6546 32280 6552 32292
rect 4764 32252 6552 32280
rect 4764 32240 4770 32252
rect 6546 32240 6552 32252
rect 6604 32240 6610 32292
rect 6365 32215 6423 32221
rect 6365 32181 6377 32215
rect 6411 32212 6423 32215
rect 6454 32212 6460 32224
rect 6411 32184 6460 32212
rect 6411 32181 6423 32184
rect 6365 32175 6423 32181
rect 6454 32172 6460 32184
rect 6512 32172 6518 32224
rect 6638 32172 6644 32224
rect 6696 32212 6702 32224
rect 6748 32212 6776 32379
rect 6914 32376 6920 32388
rect 6972 32376 6978 32428
rect 7006 32376 7012 32428
rect 7064 32416 7070 32428
rect 7576 32416 7604 32515
rect 9950 32484 9956 32496
rect 9911 32456 9956 32484
rect 9950 32444 9956 32456
rect 10008 32444 10014 32496
rect 10060 32484 10088 32524
rect 11609 32521 11621 32555
rect 11655 32552 11667 32555
rect 11974 32552 11980 32564
rect 11655 32524 11980 32552
rect 11655 32521 11667 32524
rect 11609 32515 11667 32521
rect 11974 32512 11980 32524
rect 12032 32512 12038 32564
rect 12406 32524 23796 32552
rect 12406 32484 12434 32524
rect 14550 32484 14556 32496
rect 10060 32456 12434 32484
rect 14511 32456 14556 32484
rect 14550 32444 14556 32456
rect 14608 32444 14614 32496
rect 15010 32484 15016 32496
rect 14971 32456 15016 32484
rect 15010 32444 15016 32456
rect 15068 32444 15074 32496
rect 15197 32487 15255 32493
rect 15197 32453 15209 32487
rect 15243 32484 15255 32487
rect 15470 32484 15476 32496
rect 15243 32456 15476 32484
rect 15243 32453 15255 32456
rect 15197 32447 15255 32453
rect 15470 32444 15476 32456
rect 15528 32484 15534 32496
rect 17037 32487 17095 32493
rect 15528 32456 16804 32484
rect 15528 32444 15534 32456
rect 7064 32388 7604 32416
rect 9033 32419 9091 32425
rect 7064 32376 7070 32388
rect 9033 32385 9045 32419
rect 9079 32416 9091 32419
rect 9122 32416 9128 32428
rect 9079 32388 9128 32416
rect 9079 32385 9091 32388
rect 9033 32379 9091 32385
rect 9122 32376 9128 32388
rect 9180 32416 9186 32428
rect 9398 32416 9404 32428
rect 9180 32388 9404 32416
rect 9180 32376 9186 32388
rect 9398 32376 9404 32388
rect 9456 32416 9462 32428
rect 9769 32419 9827 32425
rect 9769 32416 9781 32419
rect 9456 32388 9781 32416
rect 9456 32376 9462 32388
rect 9769 32385 9781 32388
rect 9815 32385 9827 32419
rect 12710 32416 12716 32428
rect 12768 32425 12774 32428
rect 12680 32388 12716 32416
rect 9769 32379 9827 32385
rect 12710 32376 12716 32388
rect 12768 32379 12780 32425
rect 12986 32416 12992 32428
rect 12947 32388 12992 32416
rect 12768 32376 12774 32379
rect 12986 32376 12992 32388
rect 13044 32376 13050 32428
rect 13906 32416 13912 32428
rect 13867 32388 13912 32416
rect 13906 32376 13912 32388
rect 13964 32376 13970 32428
rect 14093 32419 14151 32425
rect 14093 32385 14105 32419
rect 14139 32385 14151 32419
rect 14093 32379 14151 32385
rect 7282 32308 7288 32360
rect 7340 32348 7346 32360
rect 8757 32351 8815 32357
rect 8757 32348 8769 32351
rect 7340 32320 8769 32348
rect 7340 32308 7346 32320
rect 8757 32317 8769 32320
rect 8803 32317 8815 32351
rect 14108 32348 14136 32379
rect 14182 32376 14188 32428
rect 14240 32416 14246 32428
rect 14366 32425 14372 32428
rect 14323 32419 14372 32425
rect 14240 32388 14285 32416
rect 14240 32376 14246 32388
rect 14323 32385 14335 32419
rect 14369 32385 14372 32419
rect 14323 32379 14372 32385
rect 14366 32376 14372 32379
rect 14424 32376 14430 32428
rect 15102 32376 15108 32428
rect 15160 32416 15166 32428
rect 16776 32425 16804 32456
rect 17037 32453 17049 32487
rect 17083 32484 17095 32487
rect 17494 32484 17500 32496
rect 17083 32456 17500 32484
rect 17083 32453 17095 32456
rect 17037 32447 17095 32453
rect 17494 32444 17500 32456
rect 17552 32444 17558 32496
rect 21082 32484 21088 32496
rect 21043 32456 21088 32484
rect 21082 32444 21088 32456
rect 21140 32484 21146 32496
rect 21634 32484 21640 32496
rect 21140 32456 21640 32484
rect 21140 32444 21146 32456
rect 21634 32444 21640 32456
rect 21692 32444 21698 32496
rect 21818 32484 21824 32496
rect 21779 32456 21824 32484
rect 21818 32444 21824 32456
rect 21876 32444 21882 32496
rect 16669 32419 16727 32425
rect 16669 32416 16681 32419
rect 15160 32388 16681 32416
rect 15160 32376 15166 32388
rect 16669 32385 16681 32388
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 16762 32419 16820 32425
rect 16762 32385 16774 32419
rect 16808 32385 16820 32419
rect 16762 32379 16820 32385
rect 16945 32419 17003 32425
rect 16945 32385 16957 32419
rect 16991 32385 17003 32419
rect 16945 32379 17003 32385
rect 17134 32419 17192 32425
rect 17134 32385 17146 32419
rect 17180 32416 17192 32419
rect 20898 32416 20904 32428
rect 17180 32388 17264 32416
rect 20859 32388 20904 32416
rect 17180 32385 17192 32388
rect 17134 32379 17192 32385
rect 15381 32351 15439 32357
rect 15381 32348 15393 32351
rect 14108 32320 15393 32348
rect 8757 32311 8815 32317
rect 15381 32317 15393 32320
rect 15427 32317 15439 32351
rect 15381 32311 15439 32317
rect 16574 32308 16580 32360
rect 16632 32348 16638 32360
rect 16960 32348 16988 32379
rect 16632 32320 16988 32348
rect 16632 32308 16638 32320
rect 16942 32240 16948 32292
rect 17000 32280 17006 32292
rect 17236 32280 17264 32388
rect 20898 32376 20904 32388
rect 20956 32376 20962 32428
rect 22002 32376 22008 32428
rect 22060 32425 22066 32428
rect 22060 32419 22109 32425
rect 22060 32385 22063 32419
rect 22097 32385 22109 32419
rect 22186 32416 22192 32428
rect 22147 32388 22192 32416
rect 22060 32379 22109 32385
rect 22060 32376 22066 32379
rect 22186 32376 22192 32388
rect 22244 32376 22250 32428
rect 22281 32419 22339 32425
rect 22281 32385 22293 32419
rect 22327 32385 22339 32419
rect 22462 32416 22468 32428
rect 22423 32388 22468 32416
rect 22281 32379 22339 32385
rect 21269 32351 21327 32357
rect 21269 32317 21281 32351
rect 21315 32348 21327 32351
rect 22296 32348 22324 32379
rect 22462 32376 22468 32388
rect 22520 32376 22526 32428
rect 22922 32416 22928 32428
rect 22883 32388 22928 32416
rect 22922 32376 22928 32388
rect 22980 32376 22986 32428
rect 23566 32348 23572 32360
rect 21315 32320 22324 32348
rect 22940 32320 23572 32348
rect 21315 32317 21327 32320
rect 21269 32311 21327 32317
rect 17000 32252 17264 32280
rect 17000 32240 17006 32252
rect 17402 32240 17408 32292
rect 17460 32280 17466 32292
rect 22940 32280 22968 32320
rect 23566 32308 23572 32320
rect 23624 32308 23630 32360
rect 23106 32280 23112 32292
rect 17460 32252 22968 32280
rect 23067 32252 23112 32280
rect 17460 32240 17466 32252
rect 23106 32240 23112 32252
rect 23164 32240 23170 32292
rect 23768 32280 23796 32524
rect 24486 32512 24492 32564
rect 24544 32512 24550 32564
rect 28534 32512 28540 32564
rect 28592 32552 28598 32564
rect 28810 32552 28816 32564
rect 28592 32524 28816 32552
rect 28592 32512 28598 32524
rect 28810 32512 28816 32524
rect 28868 32552 28874 32564
rect 30929 32555 30987 32561
rect 30929 32552 30941 32555
rect 28868 32524 30941 32552
rect 28868 32512 28874 32524
rect 30929 32521 30941 32524
rect 30975 32521 30987 32555
rect 30929 32515 30987 32521
rect 31938 32512 31944 32564
rect 31996 32552 32002 32564
rect 35253 32555 35311 32561
rect 35253 32552 35265 32555
rect 31996 32524 35265 32552
rect 31996 32512 32002 32524
rect 35253 32521 35265 32524
rect 35299 32552 35311 32555
rect 35299 32524 36032 32552
rect 35299 32521 35311 32524
rect 35253 32515 35311 32521
rect 24504 32484 24532 32512
rect 24136 32456 24532 32484
rect 24136 32425 24164 32456
rect 24670 32444 24676 32496
rect 24728 32484 24734 32496
rect 24854 32484 24860 32496
rect 24728 32456 24860 32484
rect 24728 32444 24734 32456
rect 24854 32444 24860 32456
rect 24912 32444 24918 32496
rect 27338 32484 27344 32496
rect 27299 32456 27344 32484
rect 27338 32444 27344 32456
rect 27396 32444 27402 32496
rect 32677 32487 32735 32493
rect 32677 32453 32689 32487
rect 32723 32484 32735 32487
rect 33134 32484 33140 32496
rect 32723 32456 33140 32484
rect 32723 32453 32735 32456
rect 32677 32447 32735 32453
rect 33134 32444 33140 32456
rect 33192 32444 33198 32496
rect 35066 32444 35072 32496
rect 35124 32484 35130 32496
rect 35342 32484 35348 32496
rect 35124 32456 35348 32484
rect 35124 32444 35130 32456
rect 35342 32444 35348 32456
rect 35400 32484 35406 32496
rect 35805 32487 35863 32493
rect 35805 32484 35817 32487
rect 35400 32456 35817 32484
rect 35400 32444 35406 32456
rect 35805 32453 35817 32456
rect 35851 32453 35863 32487
rect 36004 32484 36032 32524
rect 36078 32512 36084 32564
rect 36136 32552 36142 32564
rect 36173 32555 36231 32561
rect 36173 32552 36185 32555
rect 36136 32524 36185 32552
rect 36136 32512 36142 32524
rect 36173 32521 36185 32524
rect 36219 32521 36231 32555
rect 36173 32515 36231 32521
rect 36262 32484 36268 32496
rect 36004 32456 36268 32484
rect 35805 32447 35863 32453
rect 36262 32444 36268 32456
rect 36320 32444 36326 32496
rect 24121 32419 24179 32425
rect 24121 32385 24133 32419
rect 24167 32385 24179 32419
rect 24284 32419 24342 32425
rect 24284 32416 24296 32419
rect 24121 32379 24179 32385
rect 24228 32388 24296 32416
rect 23842 32308 23848 32360
rect 23900 32348 23906 32360
rect 24228 32348 24256 32388
rect 24284 32385 24296 32388
rect 24330 32385 24342 32419
rect 24284 32379 24342 32385
rect 24384 32419 24442 32425
rect 24384 32385 24396 32419
rect 24430 32385 24442 32419
rect 24384 32379 24442 32385
rect 24535 32419 24593 32425
rect 24535 32385 24547 32419
rect 24581 32416 24593 32419
rect 25222 32416 25228 32428
rect 24581 32388 25228 32416
rect 24581 32385 24593 32388
rect 24535 32379 24593 32385
rect 23900 32320 24256 32348
rect 24399 32348 24427 32379
rect 25222 32376 25228 32388
rect 25280 32376 25286 32428
rect 28258 32376 28264 32428
rect 28316 32416 28322 32428
rect 29805 32419 29863 32425
rect 29805 32416 29817 32419
rect 28316 32388 29817 32416
rect 28316 32376 28322 32388
rect 29805 32385 29817 32388
rect 29851 32385 29863 32419
rect 29805 32379 29863 32385
rect 31754 32376 31760 32428
rect 31812 32416 31818 32428
rect 31938 32416 31944 32428
rect 31812 32388 31944 32416
rect 31812 32376 31818 32388
rect 31938 32376 31944 32388
rect 31996 32376 32002 32428
rect 32582 32416 32588 32428
rect 32543 32388 32588 32416
rect 32582 32376 32588 32388
rect 32640 32376 32646 32428
rect 32766 32376 32772 32428
rect 32824 32416 32830 32428
rect 32953 32419 33011 32425
rect 32824 32388 32869 32416
rect 32824 32376 32830 32388
rect 32953 32385 32965 32419
rect 32999 32416 33011 32419
rect 34514 32416 34520 32428
rect 32999 32388 34520 32416
rect 32999 32385 33011 32388
rect 32953 32379 33011 32385
rect 34514 32376 34520 32388
rect 34572 32376 34578 32428
rect 35989 32419 36047 32425
rect 35989 32385 36001 32419
rect 36035 32416 36047 32419
rect 36078 32416 36084 32428
rect 36035 32388 36084 32416
rect 36035 32385 36047 32388
rect 35989 32379 36047 32385
rect 36078 32376 36084 32388
rect 36136 32376 36142 32428
rect 24854 32348 24860 32360
rect 24399 32320 24860 32348
rect 23900 32308 23906 32320
rect 24854 32308 24860 32320
rect 24912 32308 24918 32360
rect 29549 32351 29607 32357
rect 29549 32348 29561 32351
rect 28644 32320 29561 32348
rect 28534 32280 28540 32292
rect 23768 32252 28540 32280
rect 28534 32240 28540 32252
rect 28592 32240 28598 32292
rect 10134 32212 10140 32224
rect 6696 32184 6776 32212
rect 10095 32184 10140 32212
rect 6696 32172 6702 32184
rect 10134 32172 10140 32184
rect 10192 32172 10198 32224
rect 17313 32215 17371 32221
rect 17313 32181 17325 32215
rect 17359 32212 17371 32215
rect 17678 32212 17684 32224
rect 17359 32184 17684 32212
rect 17359 32181 17371 32184
rect 17313 32175 17371 32181
rect 17678 32172 17684 32184
rect 17736 32172 17742 32224
rect 17770 32172 17776 32224
rect 17828 32212 17834 32224
rect 23124 32212 23152 32240
rect 23934 32212 23940 32224
rect 17828 32184 23940 32212
rect 17828 32172 17834 32184
rect 23934 32172 23940 32184
rect 23992 32172 23998 32224
rect 24762 32212 24768 32224
rect 24723 32184 24768 32212
rect 24762 32172 24768 32184
rect 24820 32172 24826 32224
rect 26786 32172 26792 32224
rect 26844 32212 26850 32224
rect 28644 32221 28672 32320
rect 29549 32317 29561 32320
rect 29595 32317 29607 32351
rect 29549 32311 29607 32317
rect 28629 32215 28687 32221
rect 28629 32212 28641 32215
rect 26844 32184 28641 32212
rect 26844 32172 26850 32184
rect 28629 32181 28641 32184
rect 28675 32181 28687 32215
rect 28629 32175 28687 32181
rect 32214 32172 32220 32224
rect 32272 32212 32278 32224
rect 32401 32215 32459 32221
rect 32401 32212 32413 32215
rect 32272 32184 32413 32212
rect 32272 32172 32278 32184
rect 32401 32181 32413 32184
rect 32447 32181 32459 32215
rect 58158 32212 58164 32224
rect 58119 32184 58164 32212
rect 32401 32175 32459 32181
rect 58158 32172 58164 32184
rect 58216 32172 58222 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 6822 31968 6828 32020
rect 6880 32008 6886 32020
rect 7009 32011 7067 32017
rect 7009 32008 7021 32011
rect 6880 31980 7021 32008
rect 6880 31968 6886 31980
rect 7009 31977 7021 31980
rect 7055 31977 7067 32011
rect 7009 31971 7067 31977
rect 7024 31872 7052 31971
rect 7374 31968 7380 32020
rect 7432 32008 7438 32020
rect 7432 31980 9904 32008
rect 7432 31968 7438 31980
rect 9876 31940 9904 31980
rect 9950 31968 9956 32020
rect 10008 32008 10014 32020
rect 10321 32011 10379 32017
rect 10321 32008 10333 32011
rect 10008 31980 10333 32008
rect 10008 31968 10014 31980
rect 10321 31977 10333 31980
rect 10367 31977 10379 32011
rect 10321 31971 10379 31977
rect 12529 32011 12587 32017
rect 12529 31977 12541 32011
rect 12575 32008 12587 32011
rect 12710 32008 12716 32020
rect 12575 31980 12716 32008
rect 12575 31977 12587 31980
rect 12529 31971 12587 31977
rect 12710 31968 12716 31980
rect 12768 31968 12774 32020
rect 16758 32008 16764 32020
rect 16132 31980 16764 32008
rect 16132 31940 16160 31980
rect 16758 31968 16764 31980
rect 16816 31968 16822 32020
rect 17494 32008 17500 32020
rect 17455 31980 17500 32008
rect 17494 31968 17500 31980
rect 17552 31968 17558 32020
rect 19981 32011 20039 32017
rect 19981 31977 19993 32011
rect 20027 32008 20039 32011
rect 20898 32008 20904 32020
rect 20027 31980 20904 32008
rect 20027 31977 20039 31980
rect 19981 31971 20039 31977
rect 20898 31968 20904 31980
rect 20956 32008 20962 32020
rect 22833 32011 22891 32017
rect 20956 31980 22094 32008
rect 20956 31968 20962 31980
rect 9876 31912 16160 31940
rect 8938 31872 8944 31884
rect 7024 31844 8944 31872
rect 8938 31832 8944 31844
rect 8996 31832 9002 31884
rect 16114 31872 16120 31884
rect 16075 31844 16120 31872
rect 16114 31832 16120 31844
rect 16172 31832 16178 31884
rect 1857 31807 1915 31813
rect 1857 31773 1869 31807
rect 1903 31804 1915 31807
rect 1946 31804 1952 31816
rect 1903 31776 1952 31804
rect 1903 31773 1915 31776
rect 1857 31767 1915 31773
rect 1946 31764 1952 31776
rect 2004 31764 2010 31816
rect 5718 31804 5724 31816
rect 5631 31776 5724 31804
rect 5718 31764 5724 31776
rect 5776 31804 5782 31816
rect 8021 31807 8079 31813
rect 8021 31804 8033 31807
rect 5776 31776 8033 31804
rect 5776 31764 5782 31776
rect 8021 31773 8033 31776
rect 8067 31804 8079 31807
rect 11054 31804 11060 31816
rect 8067 31776 11060 31804
rect 8067 31773 8079 31776
rect 8021 31767 8079 31773
rect 11054 31764 11060 31776
rect 11112 31764 11118 31816
rect 12710 31764 12716 31816
rect 12768 31804 12774 31816
rect 12805 31807 12863 31813
rect 12805 31804 12817 31807
rect 12768 31776 12817 31804
rect 12768 31764 12774 31776
rect 12805 31773 12817 31776
rect 12851 31773 12863 31807
rect 12805 31767 12863 31773
rect 12894 31801 12952 31807
rect 12894 31767 12906 31801
rect 12940 31767 12952 31801
rect 12894 31761 12952 31767
rect 12986 31764 12992 31816
rect 13044 31804 13050 31816
rect 13044 31776 13089 31804
rect 13044 31764 13050 31776
rect 13170 31764 13176 31816
rect 13228 31804 13234 31816
rect 16384 31807 16442 31813
rect 13228 31776 13273 31804
rect 13228 31764 13234 31776
rect 16384 31773 16396 31807
rect 16430 31804 16442 31807
rect 16666 31804 16672 31816
rect 16430 31776 16672 31804
rect 16430 31773 16442 31776
rect 16384 31767 16442 31773
rect 16666 31764 16672 31776
rect 16724 31764 16730 31816
rect 16758 31764 16764 31816
rect 16816 31804 16822 31816
rect 17512 31804 17540 31968
rect 22066 31872 22094 31980
rect 22833 31977 22845 32011
rect 22879 32008 22891 32011
rect 22922 32008 22928 32020
rect 22879 31980 22928 32008
rect 22879 31977 22891 31980
rect 22833 31971 22891 31977
rect 22922 31968 22928 31980
rect 22980 32008 22986 32020
rect 27154 32008 27160 32020
rect 22980 31980 27160 32008
rect 22980 31968 22986 31980
rect 27154 31968 27160 31980
rect 27212 31968 27218 32020
rect 27706 32008 27712 32020
rect 27667 31980 27712 32008
rect 27706 31968 27712 31980
rect 27764 31968 27770 32020
rect 28258 32008 28264 32020
rect 28219 31980 28264 32008
rect 28258 31968 28264 31980
rect 28316 31968 28322 32020
rect 28534 31968 28540 32020
rect 28592 32008 28598 32020
rect 30101 32011 30159 32017
rect 30101 32008 30113 32011
rect 28592 31980 30113 32008
rect 28592 31968 28598 31980
rect 30101 31977 30113 31980
rect 30147 32008 30159 32011
rect 30374 32008 30380 32020
rect 30147 31980 30380 32008
rect 30147 31977 30159 31980
rect 30101 31971 30159 31977
rect 30374 31968 30380 31980
rect 30432 31968 30438 32020
rect 31662 32008 31668 32020
rect 30484 31980 31668 32008
rect 26329 31943 26387 31949
rect 26329 31909 26341 31943
rect 26375 31940 26387 31943
rect 30484 31940 30512 31980
rect 31662 31968 31668 31980
rect 31720 31968 31726 32020
rect 35986 32008 35992 32020
rect 35947 31980 35992 32008
rect 35986 31968 35992 31980
rect 36044 31968 36050 32020
rect 36078 31968 36084 32020
rect 36136 32008 36142 32020
rect 37001 32011 37059 32017
rect 37001 32008 37013 32011
rect 36136 31980 37013 32008
rect 36136 31968 36142 31980
rect 37001 31977 37013 31980
rect 37047 31977 37059 32011
rect 37001 31971 37059 31977
rect 26375 31912 30512 31940
rect 31205 31943 31263 31949
rect 26375 31909 26387 31912
rect 26329 31903 26387 31909
rect 31205 31909 31217 31943
rect 31251 31940 31263 31943
rect 31294 31940 31300 31952
rect 31251 31912 31300 31940
rect 31251 31909 31263 31912
rect 31205 31903 31263 31909
rect 31294 31900 31300 31912
rect 31352 31900 31358 31952
rect 31754 31900 31760 31952
rect 31812 31940 31818 31952
rect 32217 31943 32275 31949
rect 32217 31940 32229 31943
rect 31812 31912 32229 31940
rect 31812 31900 31818 31912
rect 32217 31909 32229 31912
rect 32263 31909 32275 31943
rect 32217 31903 32275 31909
rect 22830 31872 22836 31884
rect 22066 31844 22836 31872
rect 22830 31832 22836 31844
rect 22888 31832 22894 31884
rect 25777 31875 25835 31881
rect 25777 31841 25789 31875
rect 25823 31872 25835 31875
rect 26234 31872 26240 31884
rect 25823 31844 26240 31872
rect 25823 31841 25835 31844
rect 25777 31835 25835 31841
rect 26234 31832 26240 31844
rect 26292 31872 26298 31884
rect 26786 31872 26792 31884
rect 26292 31844 26792 31872
rect 26292 31832 26298 31844
rect 26786 31832 26792 31844
rect 26844 31832 26850 31884
rect 30098 31872 30104 31884
rect 28644 31844 30104 31872
rect 18141 31807 18199 31813
rect 18141 31804 18153 31807
rect 16816 31776 17448 31804
rect 17512 31776 18153 31804
rect 16816 31764 16822 31776
rect 2124 31739 2182 31745
rect 2124 31705 2136 31739
rect 2170 31736 2182 31739
rect 2590 31736 2596 31748
rect 2170 31708 2596 31736
rect 2170 31705 2182 31708
rect 2124 31699 2182 31705
rect 2590 31696 2596 31708
rect 2648 31696 2654 31748
rect 9208 31739 9266 31745
rect 9208 31705 9220 31739
rect 9254 31736 9266 31739
rect 9674 31736 9680 31748
rect 9254 31708 9680 31736
rect 9254 31705 9266 31708
rect 9208 31699 9266 31705
rect 9674 31696 9680 31708
rect 9732 31696 9738 31748
rect 3237 31671 3295 31677
rect 3237 31637 3249 31671
rect 3283 31668 3295 31671
rect 3878 31668 3884 31680
rect 3283 31640 3884 31668
rect 3283 31637 3295 31640
rect 3237 31631 3295 31637
rect 3878 31628 3884 31640
rect 3936 31628 3942 31680
rect 12909 31668 12937 31761
rect 16574 31696 16580 31748
rect 16632 31736 16638 31748
rect 16850 31736 16856 31748
rect 16632 31708 16856 31736
rect 16632 31696 16638 31708
rect 16850 31696 16856 31708
rect 16908 31696 16914 31748
rect 17420 31736 17448 31776
rect 18141 31773 18153 31776
rect 18187 31773 18199 31807
rect 18141 31767 18199 31773
rect 19426 31764 19432 31816
rect 19484 31804 19490 31816
rect 19797 31807 19855 31813
rect 19797 31804 19809 31807
rect 19484 31776 19809 31804
rect 19484 31764 19490 31776
rect 19797 31773 19809 31776
rect 19843 31804 19855 31807
rect 20441 31807 20499 31813
rect 20441 31804 20453 31807
rect 19843 31776 20453 31804
rect 19843 31773 19855 31776
rect 19797 31767 19855 31773
rect 20441 31773 20453 31776
rect 20487 31773 20499 31807
rect 20441 31767 20499 31773
rect 24762 31764 24768 31816
rect 24820 31804 24826 31816
rect 25510 31807 25568 31813
rect 25510 31804 25522 31807
rect 24820 31776 25522 31804
rect 24820 31764 24826 31776
rect 25510 31773 25522 31776
rect 25556 31773 25568 31807
rect 26510 31804 26516 31816
rect 26471 31776 26516 31804
rect 25510 31767 25568 31773
rect 26510 31764 26516 31776
rect 26568 31764 26574 31816
rect 27706 31764 27712 31816
rect 27764 31804 27770 31816
rect 28644 31813 28672 31844
rect 30098 31832 30104 31844
rect 30156 31832 30162 31884
rect 32582 31872 32588 31884
rect 31404 31844 32588 31872
rect 28537 31807 28595 31813
rect 28537 31804 28549 31807
rect 27764 31776 28549 31804
rect 27764 31764 27770 31776
rect 28537 31773 28549 31776
rect 28583 31773 28595 31807
rect 28537 31767 28595 31773
rect 28629 31807 28687 31813
rect 28629 31773 28641 31807
rect 28675 31773 28687 31807
rect 28629 31767 28687 31773
rect 28718 31764 28724 31816
rect 28776 31804 28782 31816
rect 31404 31813 31432 31844
rect 28905 31807 28963 31813
rect 28776 31776 28821 31804
rect 28776 31764 28782 31776
rect 28905 31773 28917 31807
rect 28951 31804 28963 31807
rect 31389 31807 31447 31813
rect 28951 31776 28985 31804
rect 28951 31773 28963 31776
rect 28905 31767 28963 31773
rect 31389 31773 31401 31807
rect 31435 31773 31447 31807
rect 31389 31767 31447 31773
rect 17586 31736 17592 31748
rect 17420 31708 17592 31736
rect 17586 31696 17592 31708
rect 17644 31736 17650 31748
rect 17957 31739 18015 31745
rect 17957 31736 17969 31739
rect 17644 31708 17969 31736
rect 17644 31696 17650 31708
rect 17957 31705 17969 31708
rect 18003 31705 18015 31739
rect 17957 31699 18015 31705
rect 22922 31696 22928 31748
rect 22980 31736 22986 31748
rect 22980 31708 26556 31736
rect 22980 31696 22986 31708
rect 26528 31680 26556 31708
rect 28442 31696 28448 31748
rect 28500 31736 28506 31748
rect 28920 31736 28948 31767
rect 31478 31764 31484 31816
rect 31536 31804 31542 31816
rect 31757 31807 31815 31813
rect 31536 31776 31581 31804
rect 31536 31764 31542 31776
rect 31757 31773 31769 31807
rect 31803 31804 31815 31807
rect 31938 31804 31944 31816
rect 31803 31776 31944 31804
rect 31803 31773 31815 31776
rect 31757 31767 31815 31773
rect 31938 31764 31944 31776
rect 31996 31764 32002 31816
rect 32306 31764 32312 31816
rect 32364 31804 32370 31816
rect 32416 31813 32444 31844
rect 32582 31832 32588 31844
rect 32640 31832 32646 31884
rect 32674 31832 32680 31884
rect 32732 31872 32738 31884
rect 32732 31844 32812 31872
rect 32732 31832 32738 31844
rect 32401 31807 32459 31813
rect 32401 31804 32413 31807
rect 32364 31776 32413 31804
rect 32364 31764 32370 31776
rect 32401 31773 32413 31776
rect 32447 31773 32459 31807
rect 32401 31767 32459 31773
rect 32490 31764 32496 31816
rect 32548 31804 32554 31816
rect 32784 31813 32812 31844
rect 32769 31807 32827 31813
rect 32548 31776 32593 31804
rect 32548 31764 32554 31776
rect 32769 31773 32781 31807
rect 32815 31773 32827 31807
rect 35802 31804 35808 31816
rect 35763 31776 35808 31804
rect 32769 31767 32827 31773
rect 35802 31764 35808 31776
rect 35860 31764 35866 31816
rect 36538 31764 36544 31816
rect 36596 31804 36602 31816
rect 38114 31807 38172 31813
rect 38114 31804 38126 31807
rect 36596 31776 38126 31804
rect 36596 31764 36602 31776
rect 38114 31773 38126 31776
rect 38160 31773 38172 31807
rect 38114 31767 38172 31773
rect 38381 31807 38439 31813
rect 38381 31773 38393 31807
rect 38427 31804 38439 31807
rect 38562 31804 38568 31816
rect 38427 31776 38568 31804
rect 38427 31773 38439 31776
rect 38381 31767 38439 31773
rect 38562 31764 38568 31776
rect 38620 31764 38626 31816
rect 28500 31708 28948 31736
rect 28500 31696 28506 31708
rect 29822 31696 29828 31748
rect 29880 31736 29886 31748
rect 30009 31739 30067 31745
rect 30009 31736 30021 31739
rect 29880 31708 30021 31736
rect 29880 31696 29886 31708
rect 30009 31705 30021 31708
rect 30055 31705 30067 31739
rect 30009 31699 30067 31705
rect 31573 31739 31631 31745
rect 31573 31705 31585 31739
rect 31619 31736 31631 31739
rect 32585 31739 32643 31745
rect 32585 31736 32597 31739
rect 31619 31708 32597 31736
rect 31619 31705 31631 31708
rect 31573 31699 31631 31705
rect 32585 31705 32597 31708
rect 32631 31736 32643 31739
rect 32674 31736 32680 31748
rect 32631 31708 32680 31736
rect 32631 31705 32643 31708
rect 32585 31699 32643 31705
rect 32674 31696 32680 31708
rect 32732 31696 32738 31748
rect 35342 31696 35348 31748
rect 35400 31736 35406 31748
rect 35621 31739 35679 31745
rect 35621 31736 35633 31739
rect 35400 31708 35633 31736
rect 35400 31696 35406 31708
rect 35621 31705 35633 31708
rect 35667 31705 35679 31739
rect 35621 31699 35679 31705
rect 13262 31668 13268 31680
rect 12909 31640 13268 31668
rect 13262 31628 13268 31640
rect 13320 31628 13326 31680
rect 14185 31671 14243 31677
rect 14185 31637 14197 31671
rect 14231 31668 14243 31671
rect 14366 31668 14372 31680
rect 14231 31640 14372 31668
rect 14231 31637 14243 31640
rect 14185 31631 14243 31637
rect 14366 31628 14372 31640
rect 14424 31668 14430 31680
rect 17310 31668 17316 31680
rect 14424 31640 17316 31668
rect 14424 31628 14430 31640
rect 17310 31628 17316 31640
rect 17368 31628 17374 31680
rect 18322 31668 18328 31680
rect 18283 31640 18328 31668
rect 18322 31628 18328 31640
rect 18380 31628 18386 31680
rect 24394 31668 24400 31680
rect 24355 31640 24400 31668
rect 24394 31628 24400 31640
rect 24452 31628 24458 31680
rect 26510 31628 26516 31680
rect 26568 31668 26574 31680
rect 31110 31668 31116 31680
rect 26568 31640 31116 31668
rect 26568 31628 26574 31640
rect 31110 31628 31116 31640
rect 31168 31628 31174 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 2958 31424 2964 31476
rect 3016 31464 3022 31476
rect 3418 31464 3424 31476
rect 3016 31436 3424 31464
rect 3016 31424 3022 31436
rect 3418 31424 3424 31436
rect 3476 31424 3482 31476
rect 3786 31424 3792 31476
rect 3844 31464 3850 31476
rect 4062 31464 4068 31476
rect 3844 31436 4068 31464
rect 3844 31424 3850 31436
rect 4062 31424 4068 31436
rect 4120 31424 4126 31476
rect 9674 31464 9680 31476
rect 9635 31436 9680 31464
rect 9674 31424 9680 31436
rect 9732 31424 9738 31476
rect 13170 31424 13176 31476
rect 13228 31464 13234 31476
rect 13449 31467 13507 31473
rect 13449 31464 13461 31467
rect 13228 31436 13461 31464
rect 13228 31424 13234 31436
rect 13449 31433 13461 31436
rect 13495 31433 13507 31467
rect 16666 31464 16672 31476
rect 16627 31436 16672 31464
rect 13449 31427 13507 31433
rect 16666 31424 16672 31436
rect 16724 31424 16730 31476
rect 17126 31464 17132 31476
rect 17052 31436 17132 31464
rect 6454 31356 6460 31408
rect 6512 31396 6518 31408
rect 6610 31399 6668 31405
rect 6610 31396 6622 31399
rect 6512 31368 6622 31396
rect 6512 31356 6518 31368
rect 6610 31365 6622 31368
rect 6656 31365 6668 31399
rect 6610 31359 6668 31365
rect 12710 31356 12716 31408
rect 12768 31396 12774 31408
rect 14001 31399 14059 31405
rect 14001 31396 14013 31399
rect 12768 31368 14013 31396
rect 12768 31356 12774 31368
rect 14001 31365 14013 31368
rect 14047 31396 14059 31399
rect 14047 31368 16574 31396
rect 14047 31365 14059 31368
rect 14001 31359 14059 31365
rect 2130 31328 2136 31340
rect 2091 31300 2136 31328
rect 2130 31288 2136 31300
rect 2188 31288 2194 31340
rect 2400 31331 2458 31337
rect 2400 31297 2412 31331
rect 2446 31328 2458 31331
rect 2682 31328 2688 31340
rect 2446 31300 2688 31328
rect 2446 31297 2458 31300
rect 2400 31291 2458 31297
rect 2682 31288 2688 31300
rect 2740 31288 2746 31340
rect 9858 31288 9864 31340
rect 9916 31337 9922 31340
rect 9916 31331 9965 31337
rect 9916 31297 9919 31331
rect 9953 31297 9965 31331
rect 9916 31291 9965 31297
rect 9916 31288 9922 31291
rect 10023 31288 10029 31340
rect 10081 31337 10087 31340
rect 10081 31331 10100 31337
rect 10088 31297 10100 31331
rect 10081 31291 10100 31297
rect 10081 31288 10087 31291
rect 10134 31288 10140 31340
rect 10192 31337 10198 31340
rect 10192 31328 10200 31337
rect 10321 31331 10379 31337
rect 10192 31300 10237 31328
rect 10192 31291 10200 31300
rect 10321 31297 10333 31331
rect 10367 31297 10379 31331
rect 10321 31291 10379 31297
rect 10192 31288 10198 31291
rect 6178 31220 6184 31272
rect 6236 31260 6242 31272
rect 6365 31263 6423 31269
rect 6365 31260 6377 31263
rect 6236 31232 6377 31260
rect 6236 31220 6242 31232
rect 6365 31229 6377 31232
rect 6411 31229 6423 31263
rect 6365 31223 6423 31229
rect 10226 31220 10232 31272
rect 10284 31260 10290 31272
rect 10336 31260 10364 31291
rect 10502 31288 10508 31340
rect 10560 31328 10566 31340
rect 10873 31331 10931 31337
rect 10873 31328 10885 31331
rect 10560 31300 10885 31328
rect 10560 31288 10566 31300
rect 10873 31297 10885 31300
rect 10919 31328 10931 31331
rect 14366 31328 14372 31340
rect 10919 31300 14372 31328
rect 10919 31297 10931 31300
rect 10873 31291 10931 31297
rect 14366 31288 14372 31300
rect 14424 31288 14430 31340
rect 16546 31328 16574 31368
rect 17052 31337 17080 31436
rect 17126 31424 17132 31436
rect 17184 31424 17190 31476
rect 21910 31424 21916 31476
rect 21968 31464 21974 31476
rect 22005 31467 22063 31473
rect 22005 31464 22017 31467
rect 21968 31436 22017 31464
rect 21968 31424 21974 31436
rect 22005 31433 22017 31436
rect 22051 31433 22063 31467
rect 22005 31427 22063 31433
rect 23842 31424 23848 31476
rect 23900 31464 23906 31476
rect 24213 31467 24271 31473
rect 24213 31464 24225 31467
rect 23900 31436 24225 31464
rect 23900 31424 23906 31436
rect 24213 31433 24225 31436
rect 24259 31433 24271 31467
rect 25498 31464 25504 31476
rect 24213 31427 24271 31433
rect 24320 31436 25504 31464
rect 18322 31396 18328 31408
rect 17144 31368 18328 31396
rect 17144 31337 17172 31368
rect 18322 31356 18328 31368
rect 18380 31356 18386 31408
rect 22186 31396 22192 31408
rect 20180 31368 22192 31396
rect 16945 31331 17003 31337
rect 16945 31328 16957 31331
rect 16546 31300 16957 31328
rect 16945 31297 16957 31300
rect 16991 31297 17003 31331
rect 16945 31291 17003 31297
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31297 17095 31331
rect 17037 31291 17095 31297
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31328 17371 31331
rect 17954 31328 17960 31340
rect 17359 31300 17960 31328
rect 17359 31297 17371 31300
rect 17313 31291 17371 31297
rect 10284 31232 10364 31260
rect 16960 31260 16988 31291
rect 17954 31288 17960 31300
rect 18012 31328 18018 31340
rect 19058 31328 19064 31340
rect 18012 31300 19064 31328
rect 18012 31288 18018 31300
rect 19058 31288 19064 31300
rect 19116 31288 19122 31340
rect 20180 31337 20208 31368
rect 22186 31356 22192 31368
rect 22244 31356 22250 31408
rect 24320 31396 24348 31436
rect 25498 31424 25504 31436
rect 25556 31424 25562 31476
rect 26145 31467 26203 31473
rect 26145 31433 26157 31467
rect 26191 31464 26203 31467
rect 26510 31464 26516 31476
rect 26191 31436 26516 31464
rect 26191 31433 26203 31436
rect 26145 31427 26203 31433
rect 26510 31424 26516 31436
rect 26568 31424 26574 31476
rect 28994 31424 29000 31476
rect 29052 31424 29058 31476
rect 30374 31424 30380 31476
rect 30432 31464 30438 31476
rect 30653 31467 30711 31473
rect 30653 31464 30665 31467
rect 30432 31436 30665 31464
rect 30432 31424 30438 31436
rect 30653 31433 30665 31436
rect 30699 31433 30711 31467
rect 30653 31427 30711 31433
rect 23492 31368 24348 31396
rect 24581 31399 24639 31405
rect 20165 31331 20223 31337
rect 19269 31300 20116 31328
rect 19269 31260 19297 31300
rect 19889 31263 19947 31269
rect 19889 31260 19901 31263
rect 16960 31232 19297 31260
rect 19352 31232 19901 31260
rect 10284 31220 10290 31232
rect 9858 31152 9864 31204
rect 9916 31192 9922 31204
rect 10502 31192 10508 31204
rect 9916 31164 10508 31192
rect 9916 31152 9922 31164
rect 10502 31152 10508 31164
rect 10560 31152 10566 31204
rect 11698 31152 11704 31204
rect 11756 31192 11762 31204
rect 14182 31192 14188 31204
rect 11756 31164 14188 31192
rect 11756 31152 11762 31164
rect 14182 31152 14188 31164
rect 14240 31152 14246 31204
rect 17420 31136 17448 31232
rect 19352 31136 19380 31232
rect 19889 31229 19901 31232
rect 19935 31229 19947 31263
rect 20088 31260 20116 31300
rect 20165 31297 20177 31331
rect 20211 31297 20223 31331
rect 20165 31291 20223 31297
rect 21269 31331 21327 31337
rect 21269 31297 21281 31331
rect 21315 31328 21327 31331
rect 21821 31331 21879 31337
rect 21821 31328 21833 31331
rect 21315 31300 21833 31328
rect 21315 31297 21327 31300
rect 21269 31291 21327 31297
rect 21821 31297 21833 31300
rect 21867 31328 21879 31331
rect 22922 31328 22928 31340
rect 21867 31300 22928 31328
rect 21867 31297 21879 31300
rect 21821 31291 21879 31297
rect 22922 31288 22928 31300
rect 22980 31288 22986 31340
rect 23492 31337 23520 31368
rect 24581 31365 24593 31399
rect 24627 31396 24639 31399
rect 24670 31396 24676 31408
rect 24627 31368 24676 31396
rect 24627 31365 24639 31368
rect 24581 31359 24639 31365
rect 24670 31356 24676 31368
rect 24728 31356 24734 31408
rect 28721 31399 28779 31405
rect 28721 31365 28733 31399
rect 28767 31396 28779 31399
rect 29012 31396 29040 31424
rect 28767 31368 29040 31396
rect 32585 31399 32643 31405
rect 28767 31365 28779 31368
rect 28721 31359 28779 31365
rect 32585 31365 32597 31399
rect 32631 31396 32643 31399
rect 36078 31396 36084 31408
rect 32631 31368 36084 31396
rect 32631 31365 32643 31368
rect 32585 31359 32643 31365
rect 36078 31356 36084 31368
rect 36136 31356 36142 31408
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31328 23075 31331
rect 23477 31331 23535 31337
rect 23477 31328 23489 31331
rect 23063 31300 23489 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 23477 31297 23489 31300
rect 23523 31297 23535 31331
rect 24394 31328 24400 31340
rect 24355 31300 24400 31328
rect 23477 31291 23535 31297
rect 24394 31288 24400 31300
rect 24452 31288 24458 31340
rect 28534 31288 28540 31340
rect 28592 31328 28598 31340
rect 28629 31331 28687 31337
rect 28629 31328 28641 31331
rect 28592 31300 28641 31328
rect 28592 31288 28598 31300
rect 28629 31297 28641 31300
rect 28675 31297 28687 31331
rect 28629 31291 28687 31297
rect 28813 31331 28871 31337
rect 28813 31297 28825 31331
rect 28859 31297 28871 31331
rect 28813 31291 28871 31297
rect 28997 31331 29055 31337
rect 28997 31297 29009 31331
rect 29043 31328 29055 31331
rect 29270 31328 29276 31340
rect 29043 31300 29276 31328
rect 29043 31297 29055 31300
rect 28997 31291 29055 31297
rect 24946 31260 24952 31272
rect 20088 31232 24952 31260
rect 19889 31223 19947 31229
rect 24946 31220 24952 31232
rect 25004 31260 25010 31272
rect 25041 31263 25099 31269
rect 25041 31260 25053 31263
rect 25004 31232 25053 31260
rect 25004 31220 25010 31232
rect 25041 31229 25053 31232
rect 25087 31260 25099 31263
rect 26050 31260 26056 31272
rect 25087 31232 26056 31260
rect 25087 31229 25099 31232
rect 25041 31223 25099 31229
rect 26050 31220 26056 31232
rect 26108 31220 26114 31272
rect 28718 31220 28724 31272
rect 28776 31260 28782 31272
rect 28828 31260 28856 31291
rect 29270 31288 29276 31300
rect 29328 31288 29334 31340
rect 32306 31288 32312 31340
rect 32364 31328 32370 31340
rect 32493 31331 32551 31337
rect 32493 31328 32505 31331
rect 32364 31300 32505 31328
rect 32364 31288 32370 31300
rect 32493 31297 32505 31300
rect 32539 31297 32551 31331
rect 32674 31328 32680 31340
rect 32635 31300 32680 31328
rect 32493 31291 32551 31297
rect 32674 31288 32680 31300
rect 32732 31288 32738 31340
rect 32861 31331 32919 31337
rect 32861 31297 32873 31331
rect 32907 31328 32919 31331
rect 33226 31328 33232 31340
rect 32907 31300 33232 31328
rect 32907 31297 32919 31300
rect 32861 31291 32919 31297
rect 33226 31288 33232 31300
rect 33284 31288 33290 31340
rect 28776 31232 28856 31260
rect 28776 31220 28782 31232
rect 22833 31195 22891 31201
rect 22833 31161 22845 31195
rect 22879 31192 22891 31195
rect 25130 31192 25136 31204
rect 22879 31164 25136 31192
rect 22879 31161 22891 31164
rect 22833 31155 22891 31161
rect 25130 31152 25136 31164
rect 25188 31152 25194 31204
rect 25682 31152 25688 31204
rect 25740 31192 25746 31204
rect 28445 31195 28503 31201
rect 28445 31192 28457 31195
rect 25740 31164 28457 31192
rect 25740 31152 25746 31164
rect 28445 31161 28457 31164
rect 28491 31161 28503 31195
rect 28445 31155 28503 31161
rect 3510 31124 3516 31136
rect 3471 31096 3516 31124
rect 3510 31084 3516 31096
rect 3568 31084 3574 31136
rect 4062 31124 4068 31136
rect 4023 31096 4068 31124
rect 4062 31084 4068 31096
rect 4120 31084 4126 31136
rect 7098 31084 7104 31136
rect 7156 31124 7162 31136
rect 7742 31124 7748 31136
rect 7156 31096 7748 31124
rect 7156 31084 7162 31096
rect 7742 31084 7748 31096
rect 7800 31084 7806 31136
rect 12250 31124 12256 31136
rect 12211 31096 12256 31124
rect 12250 31084 12256 31096
rect 12308 31084 12314 31136
rect 12434 31084 12440 31136
rect 12492 31124 12498 31136
rect 12805 31127 12863 31133
rect 12805 31124 12817 31127
rect 12492 31096 12817 31124
rect 12492 31084 12498 31096
rect 12805 31093 12817 31096
rect 12851 31093 12863 31127
rect 12805 31087 12863 31093
rect 17402 31084 17408 31136
rect 17460 31124 17466 31136
rect 17773 31127 17831 31133
rect 17773 31124 17785 31127
rect 17460 31096 17785 31124
rect 17460 31084 17466 31096
rect 17773 31093 17785 31096
rect 17819 31093 17831 31127
rect 19334 31124 19340 31136
rect 19295 31096 19340 31124
rect 17773 31087 17831 31093
rect 19334 31084 19340 31096
rect 19392 31084 19398 31136
rect 23842 31084 23848 31136
rect 23900 31124 23906 31136
rect 24026 31124 24032 31136
rect 23900 31096 24032 31124
rect 23900 31084 23906 31096
rect 24026 31084 24032 31096
rect 24084 31084 24090 31136
rect 28994 31084 29000 31136
rect 29052 31124 29058 31136
rect 29733 31127 29791 31133
rect 29733 31124 29745 31127
rect 29052 31096 29745 31124
rect 29052 31084 29058 31096
rect 29733 31093 29745 31096
rect 29779 31124 29791 31127
rect 29822 31124 29828 31136
rect 29779 31096 29828 31124
rect 29779 31093 29791 31096
rect 29733 31087 29791 31093
rect 29822 31084 29828 31096
rect 29880 31084 29886 31136
rect 32309 31127 32367 31133
rect 32309 31093 32321 31127
rect 32355 31124 32367 31127
rect 32858 31124 32864 31136
rect 32355 31096 32864 31124
rect 32355 31093 32367 31096
rect 32309 31087 32367 31093
rect 32858 31084 32864 31096
rect 32916 31084 32922 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 2590 30920 2596 30932
rect 2551 30892 2596 30920
rect 2590 30880 2596 30892
rect 2648 30880 2654 30932
rect 7098 30880 7104 30932
rect 7156 30920 7162 30932
rect 7561 30923 7619 30929
rect 7561 30920 7573 30923
rect 7156 30892 7573 30920
rect 7156 30880 7162 30892
rect 7561 30889 7573 30892
rect 7607 30920 7619 30923
rect 8202 30920 8208 30932
rect 7607 30892 8208 30920
rect 7607 30889 7619 30892
rect 7561 30883 7619 30889
rect 8202 30880 8208 30892
rect 8260 30880 8266 30932
rect 23845 30923 23903 30929
rect 23845 30889 23857 30923
rect 23891 30920 23903 30923
rect 24670 30920 24676 30932
rect 23891 30892 24676 30920
rect 23891 30889 23903 30892
rect 23845 30883 23903 30889
rect 24670 30880 24676 30892
rect 24728 30880 24734 30932
rect 26050 30880 26056 30932
rect 26108 30920 26114 30932
rect 33686 30920 33692 30932
rect 26108 30892 33692 30920
rect 26108 30880 26114 30892
rect 33686 30880 33692 30892
rect 33744 30880 33750 30932
rect 4062 30852 4068 30864
rect 2792 30824 4068 30852
rect 2792 30648 2820 30824
rect 4062 30812 4068 30824
rect 4120 30812 4126 30864
rect 17313 30855 17371 30861
rect 17313 30821 17325 30855
rect 17359 30821 17371 30855
rect 24394 30852 24400 30864
rect 17313 30815 17371 30821
rect 22066 30824 24400 30852
rect 15473 30787 15531 30793
rect 15473 30753 15485 30787
rect 15519 30784 15531 30787
rect 16114 30784 16120 30796
rect 15519 30756 16120 30784
rect 15519 30753 15531 30756
rect 15473 30747 15531 30753
rect 16114 30744 16120 30756
rect 16172 30784 16178 30796
rect 17328 30784 17356 30815
rect 17770 30784 17776 30796
rect 16172 30756 17776 30784
rect 16172 30744 16178 30756
rect 17770 30744 17776 30756
rect 17828 30784 17834 30796
rect 19245 30787 19303 30793
rect 19245 30784 19257 30787
rect 17828 30756 19257 30784
rect 17828 30744 17834 30756
rect 19245 30753 19257 30756
rect 19291 30753 19303 30787
rect 22066 30784 22094 30824
rect 24394 30812 24400 30824
rect 24452 30812 24458 30864
rect 22925 30787 22983 30793
rect 22925 30784 22937 30787
rect 19245 30747 19303 30753
rect 21376 30756 22094 30784
rect 22480 30756 22937 30784
rect 2869 30719 2927 30725
rect 2869 30685 2881 30719
rect 2915 30685 2927 30719
rect 2869 30679 2927 30685
rect 2958 30713 3016 30719
rect 2958 30679 2970 30713
rect 3004 30679 3016 30713
rect 2875 30648 2903 30679
rect 2958 30673 3016 30679
rect 3053 30716 3111 30722
rect 3053 30682 3065 30716
rect 3099 30682 3111 30716
rect 3053 30676 3111 30682
rect 3237 30719 3295 30725
rect 3237 30685 3249 30719
rect 3283 30716 3295 30719
rect 3326 30716 3332 30728
rect 3283 30688 3332 30716
rect 3283 30685 3295 30688
rect 3237 30679 3295 30685
rect 3326 30676 3332 30688
rect 3384 30676 3390 30728
rect 3878 30676 3884 30728
rect 3936 30716 3942 30728
rect 3973 30719 4031 30725
rect 3973 30716 3985 30719
rect 3936 30688 3985 30716
rect 3936 30676 3942 30688
rect 3973 30685 3985 30688
rect 4019 30685 4031 30719
rect 3973 30679 4031 30685
rect 4157 30719 4215 30725
rect 4157 30685 4169 30719
rect 4203 30716 4215 30719
rect 4614 30716 4620 30728
rect 4203 30688 4620 30716
rect 4203 30685 4215 30688
rect 4157 30679 4215 30685
rect 4614 30676 4620 30688
rect 4672 30716 4678 30728
rect 5442 30716 5448 30728
rect 4672 30688 5448 30716
rect 4672 30676 4678 30688
rect 5442 30676 5448 30688
rect 5500 30676 5506 30728
rect 6178 30716 6184 30728
rect 6091 30688 6184 30716
rect 6178 30676 6184 30688
rect 6236 30716 6242 30728
rect 6822 30716 6828 30728
rect 6236 30688 6828 30716
rect 6236 30676 6242 30688
rect 6822 30676 6828 30688
rect 6880 30676 6886 30728
rect 9674 30716 9680 30728
rect 9635 30688 9680 30716
rect 9674 30676 9680 30688
rect 9732 30676 9738 30728
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30716 9919 30719
rect 10778 30716 10784 30728
rect 9907 30688 10784 30716
rect 9907 30685 9919 30688
rect 9861 30679 9919 30685
rect 10778 30676 10784 30688
rect 10836 30676 10842 30728
rect 11072 30688 15332 30716
rect 2792 30620 2903 30648
rect 2985 30592 3013 30673
rect 3068 30648 3096 30676
rect 6454 30657 6460 30660
rect 3789 30651 3847 30657
rect 3789 30648 3801 30651
rect 3068 30620 3801 30648
rect 3789 30617 3801 30620
rect 3835 30617 3847 30651
rect 3789 30611 3847 30617
rect 6448 30611 6460 30657
rect 6512 30648 6518 30660
rect 6512 30620 6548 30648
rect 6454 30608 6460 30611
rect 6512 30608 6518 30620
rect 11072 30592 11100 30688
rect 12161 30651 12219 30657
rect 12161 30617 12173 30651
rect 12207 30648 12219 30651
rect 12250 30648 12256 30660
rect 12207 30620 12256 30648
rect 12207 30617 12219 30620
rect 12161 30611 12219 30617
rect 12250 30608 12256 30620
rect 12308 30608 12314 30660
rect 12710 30608 12716 30660
rect 12768 30648 12774 30660
rect 13173 30651 13231 30657
rect 13173 30648 13185 30651
rect 12768 30620 13185 30648
rect 12768 30608 12774 30620
rect 13173 30617 13185 30620
rect 13219 30617 13231 30651
rect 13354 30648 13360 30660
rect 13315 30620 13360 30648
rect 13173 30611 13231 30617
rect 13354 30608 13360 30620
rect 13412 30648 13418 30660
rect 15194 30648 15200 30660
rect 15252 30657 15258 30660
rect 13412 30620 14136 30648
rect 15164 30620 15200 30648
rect 13412 30608 13418 30620
rect 2958 30540 2964 30592
rect 3016 30540 3022 30592
rect 9398 30540 9404 30592
rect 9456 30580 9462 30592
rect 9493 30583 9551 30589
rect 9493 30580 9505 30583
rect 9456 30552 9505 30580
rect 9456 30540 9462 30552
rect 9493 30549 9505 30552
rect 9539 30549 9551 30583
rect 9493 30543 9551 30549
rect 10873 30583 10931 30589
rect 10873 30549 10885 30583
rect 10919 30580 10931 30583
rect 11054 30580 11060 30592
rect 10919 30552 11060 30580
rect 10919 30549 10931 30552
rect 10873 30543 10931 30549
rect 11054 30540 11060 30552
rect 11112 30540 11118 30592
rect 12621 30583 12679 30589
rect 12621 30549 12633 30583
rect 12667 30580 12679 30583
rect 12986 30580 12992 30592
rect 12667 30552 12992 30580
rect 12667 30549 12679 30552
rect 12621 30543 12679 30549
rect 12986 30540 12992 30552
rect 13044 30540 13050 30592
rect 13541 30583 13599 30589
rect 13541 30549 13553 30583
rect 13587 30580 13599 30583
rect 13722 30580 13728 30592
rect 13587 30552 13728 30580
rect 13587 30549 13599 30552
rect 13541 30543 13599 30549
rect 13722 30540 13728 30552
rect 13780 30540 13786 30592
rect 14108 30589 14136 30620
rect 15194 30608 15200 30620
rect 15252 30611 15264 30657
rect 15304 30648 15332 30688
rect 20898 30676 20904 30728
rect 20956 30716 20962 30728
rect 21376 30725 21404 30756
rect 21269 30719 21327 30725
rect 21269 30716 21281 30719
rect 20956 30688 21281 30716
rect 20956 30676 20962 30688
rect 21269 30685 21281 30688
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 21361 30719 21419 30725
rect 21361 30685 21373 30719
rect 21407 30685 21419 30719
rect 21634 30716 21640 30728
rect 21595 30688 21640 30716
rect 21361 30679 21419 30685
rect 21634 30676 21640 30688
rect 21692 30676 21698 30728
rect 21818 30676 21824 30728
rect 21876 30716 21882 30728
rect 22480 30716 22508 30756
rect 22925 30753 22937 30756
rect 22971 30753 22983 30787
rect 22925 30747 22983 30753
rect 24946 30744 24952 30796
rect 25004 30744 25010 30796
rect 30926 30744 30932 30796
rect 30984 30784 30990 30796
rect 30984 30756 31340 30784
rect 30984 30744 30990 30756
rect 21876 30688 22508 30716
rect 21876 30676 21882 30688
rect 22554 30676 22560 30728
rect 22612 30716 22618 30728
rect 22649 30719 22707 30725
rect 22649 30716 22661 30719
rect 22612 30688 22661 30716
rect 22612 30676 22618 30688
rect 22649 30685 22661 30688
rect 22695 30685 22707 30719
rect 23658 30716 23664 30728
rect 23619 30688 23664 30716
rect 22649 30679 22707 30685
rect 23658 30676 23664 30688
rect 23716 30676 23722 30728
rect 24486 30716 24492 30728
rect 24447 30688 24492 30716
rect 24486 30676 24492 30688
rect 24544 30676 24550 30728
rect 24670 30716 24676 30728
rect 24631 30688 24676 30716
rect 24670 30676 24676 30688
rect 24728 30676 24734 30728
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30685 24823 30719
rect 24765 30679 24823 30685
rect 24857 30719 24915 30725
rect 24857 30685 24869 30719
rect 24903 30713 24915 30719
rect 24964 30713 24992 30744
rect 24903 30685 24992 30713
rect 24857 30679 24915 30685
rect 15838 30648 15844 30660
rect 15304 30620 15844 30648
rect 15252 30608 15258 30611
rect 15838 30608 15844 30620
rect 15896 30648 15902 30660
rect 16025 30651 16083 30657
rect 16025 30648 16037 30651
rect 15896 30620 16037 30648
rect 15896 30608 15902 30620
rect 16025 30617 16037 30620
rect 16071 30617 16083 30651
rect 16025 30611 16083 30617
rect 19512 30651 19570 30657
rect 19512 30617 19524 30651
rect 19558 30648 19570 30651
rect 19978 30648 19984 30660
rect 19558 30620 19984 30648
rect 19558 30617 19570 30620
rect 19512 30611 19570 30617
rect 19978 30608 19984 30620
rect 20036 30608 20042 30660
rect 21453 30651 21511 30657
rect 21453 30617 21465 30651
rect 21499 30648 21511 30651
rect 22002 30648 22008 30660
rect 21499 30620 22008 30648
rect 21499 30617 21511 30620
rect 21453 30611 21511 30617
rect 22002 30608 22008 30620
rect 22060 30608 22066 30660
rect 24780 30648 24808 30679
rect 25222 30676 25228 30728
rect 25280 30716 25286 30728
rect 25280 30688 26832 30716
rect 25280 30676 25286 30688
rect 24596 30620 24808 30648
rect 25133 30651 25191 30657
rect 24596 30592 24624 30620
rect 25133 30617 25145 30651
rect 25179 30648 25191 30651
rect 26706 30651 26764 30657
rect 26706 30648 26718 30651
rect 25179 30620 26718 30648
rect 25179 30617 25191 30620
rect 25133 30611 25191 30617
rect 26706 30617 26718 30620
rect 26752 30617 26764 30651
rect 26706 30611 26764 30617
rect 14093 30583 14151 30589
rect 14093 30549 14105 30583
rect 14139 30549 14151 30583
rect 20622 30580 20628 30592
rect 20583 30552 20628 30580
rect 14093 30543 14151 30549
rect 20622 30540 20628 30552
rect 20680 30540 20686 30592
rect 20990 30540 20996 30592
rect 21048 30580 21054 30592
rect 21085 30583 21143 30589
rect 21085 30580 21097 30583
rect 21048 30552 21097 30580
rect 21048 30540 21054 30552
rect 21085 30549 21097 30552
rect 21131 30549 21143 30583
rect 21085 30543 21143 30549
rect 24578 30540 24584 30592
rect 24636 30540 24642 30592
rect 25590 30580 25596 30592
rect 25551 30552 25596 30580
rect 25590 30540 25596 30552
rect 25648 30540 25654 30592
rect 26804 30580 26832 30688
rect 26878 30676 26884 30728
rect 26936 30716 26942 30728
rect 26973 30719 27031 30725
rect 26973 30716 26985 30719
rect 26936 30688 26985 30716
rect 26936 30676 26942 30688
rect 26973 30685 26985 30688
rect 27019 30685 27031 30719
rect 28534 30716 28540 30728
rect 28495 30688 28540 30716
rect 26973 30679 27031 30685
rect 28534 30676 28540 30688
rect 28592 30676 28598 30728
rect 28902 30716 28908 30728
rect 28863 30688 28908 30716
rect 28902 30676 28908 30688
rect 28960 30676 28966 30728
rect 30374 30676 30380 30728
rect 30432 30716 30438 30728
rect 31021 30719 31079 30725
rect 31021 30716 31033 30719
rect 30432 30688 31033 30716
rect 30432 30676 30438 30688
rect 31021 30685 31033 30688
rect 31067 30685 31079 30719
rect 31202 30716 31208 30728
rect 31163 30688 31208 30716
rect 31021 30679 31079 30685
rect 31202 30676 31208 30688
rect 31260 30676 31266 30728
rect 31312 30725 31340 30756
rect 32306 30744 32312 30796
rect 32364 30784 32370 30796
rect 32401 30787 32459 30793
rect 32401 30784 32413 30787
rect 32364 30756 32413 30784
rect 32364 30744 32370 30756
rect 32401 30753 32413 30756
rect 32447 30753 32459 30787
rect 32401 30747 32459 30753
rect 31297 30719 31355 30725
rect 31297 30685 31309 30719
rect 31343 30685 31355 30719
rect 31297 30679 31355 30685
rect 31389 30719 31447 30725
rect 31389 30685 31401 30719
rect 31435 30716 31447 30719
rect 31478 30716 31484 30728
rect 31435 30688 31484 30716
rect 31435 30685 31447 30688
rect 31389 30679 31447 30685
rect 28166 30608 28172 30660
rect 28224 30648 28230 30660
rect 28629 30651 28687 30657
rect 28629 30648 28641 30651
rect 28224 30620 28641 30648
rect 28224 30608 28230 30620
rect 28629 30617 28641 30620
rect 28675 30617 28687 30651
rect 28629 30611 28687 30617
rect 28718 30608 28724 30660
rect 28776 30648 28782 30660
rect 30561 30651 30619 30657
rect 28776 30620 28821 30648
rect 28776 30608 28782 30620
rect 30561 30617 30573 30651
rect 30607 30648 30619 30651
rect 31404 30648 31432 30679
rect 31478 30676 31484 30688
rect 31536 30676 31542 30728
rect 32125 30719 32183 30725
rect 32125 30685 32137 30719
rect 32171 30716 32183 30719
rect 32490 30716 32496 30728
rect 32171 30688 32496 30716
rect 32171 30685 32183 30688
rect 32125 30679 32183 30685
rect 32490 30676 32496 30688
rect 32548 30676 32554 30728
rect 34514 30676 34520 30728
rect 34572 30716 34578 30728
rect 34701 30719 34759 30725
rect 34701 30716 34713 30719
rect 34572 30688 34713 30716
rect 34572 30676 34578 30688
rect 34701 30685 34713 30688
rect 34747 30685 34759 30719
rect 34701 30679 34759 30685
rect 37093 30719 37151 30725
rect 37093 30685 37105 30719
rect 37139 30716 37151 30719
rect 38562 30716 38568 30728
rect 37139 30688 38568 30716
rect 37139 30685 37151 30688
rect 37093 30679 37151 30685
rect 38562 30676 38568 30688
rect 38620 30676 38626 30728
rect 58158 30716 58164 30728
rect 58119 30688 58164 30716
rect 58158 30676 58164 30688
rect 58216 30676 58222 30728
rect 30607 30620 31432 30648
rect 30607 30617 30619 30620
rect 30561 30611 30619 30617
rect 31570 30608 31576 30660
rect 31628 30648 31634 30660
rect 33781 30651 33839 30657
rect 33781 30648 33793 30651
rect 31628 30620 33793 30648
rect 31628 30608 31634 30620
rect 33781 30617 33793 30620
rect 33827 30617 33839 30651
rect 33962 30648 33968 30660
rect 33923 30620 33968 30648
rect 33781 30611 33839 30617
rect 33962 30608 33968 30620
rect 34020 30648 34026 30660
rect 34020 30620 35756 30648
rect 34020 30608 34026 30620
rect 28353 30583 28411 30589
rect 28353 30580 28365 30583
rect 26804 30552 28365 30580
rect 28353 30549 28365 30552
rect 28399 30549 28411 30583
rect 28353 30543 28411 30549
rect 31665 30583 31723 30589
rect 31665 30549 31677 30583
rect 31711 30580 31723 30583
rect 31846 30580 31852 30592
rect 31711 30552 31852 30580
rect 31711 30549 31723 30552
rect 31665 30543 31723 30549
rect 31846 30540 31852 30552
rect 31904 30540 31910 30592
rect 34149 30583 34207 30589
rect 34149 30549 34161 30583
rect 34195 30580 34207 30583
rect 34330 30580 34336 30592
rect 34195 30552 34336 30580
rect 34195 30549 34207 30552
rect 34149 30543 34207 30549
rect 34330 30540 34336 30552
rect 34388 30540 34394 30592
rect 34885 30583 34943 30589
rect 34885 30549 34897 30583
rect 34931 30580 34943 30583
rect 35342 30580 35348 30592
rect 34931 30552 35348 30580
rect 34931 30549 34943 30552
rect 34885 30543 34943 30549
rect 35342 30540 35348 30552
rect 35400 30540 35406 30592
rect 35728 30589 35756 30620
rect 35894 30608 35900 30660
rect 35952 30648 35958 30660
rect 36826 30651 36884 30657
rect 36826 30648 36838 30651
rect 35952 30620 36838 30648
rect 35952 30608 35958 30620
rect 36826 30617 36838 30620
rect 36872 30617 36884 30651
rect 36826 30611 36884 30617
rect 35713 30583 35771 30589
rect 35713 30549 35725 30583
rect 35759 30549 35771 30583
rect 35713 30543 35771 30549
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 2682 30376 2688 30388
rect 2643 30348 2688 30376
rect 2682 30336 2688 30348
rect 2740 30336 2746 30388
rect 2958 30336 2964 30388
rect 3016 30376 3022 30388
rect 3234 30376 3240 30388
rect 3016 30348 3096 30376
rect 3016 30336 3022 30348
rect 3068 30249 3096 30348
rect 3160 30348 3240 30376
rect 3160 30255 3188 30348
rect 3234 30336 3240 30348
rect 3292 30336 3298 30388
rect 6365 30379 6423 30385
rect 6365 30345 6377 30379
rect 6411 30376 6423 30379
rect 6454 30376 6460 30388
rect 6411 30348 6460 30376
rect 6411 30345 6423 30348
rect 6365 30339 6423 30345
rect 6454 30336 6460 30348
rect 6512 30336 6518 30388
rect 10778 30376 10784 30388
rect 10739 30348 10784 30376
rect 10778 30336 10784 30348
rect 10836 30336 10842 30388
rect 12989 30379 13047 30385
rect 12989 30345 13001 30379
rect 13035 30376 13047 30379
rect 13262 30376 13268 30388
rect 13035 30348 13268 30376
rect 13035 30345 13047 30348
rect 12989 30339 13047 30345
rect 13262 30336 13268 30348
rect 13320 30336 13326 30388
rect 15838 30376 15844 30388
rect 15799 30348 15844 30376
rect 15838 30336 15844 30348
rect 15896 30336 15902 30388
rect 28353 30379 28411 30385
rect 28353 30345 28365 30379
rect 28399 30345 28411 30379
rect 28353 30339 28411 30345
rect 30745 30379 30803 30385
rect 30745 30345 30757 30379
rect 30791 30376 30803 30379
rect 30926 30376 30932 30388
rect 30791 30348 30932 30376
rect 30791 30345 30803 30348
rect 30745 30339 30803 30345
rect 3970 30268 3976 30320
rect 4028 30308 4034 30320
rect 4341 30311 4399 30317
rect 4341 30308 4353 30311
rect 4028 30280 4353 30308
rect 4028 30268 4034 30280
rect 4341 30277 4353 30280
rect 4387 30277 4399 30311
rect 4341 30271 4399 30277
rect 11977 30311 12035 30317
rect 11977 30277 11989 30311
rect 12023 30308 12035 30311
rect 12618 30308 12624 30320
rect 12023 30280 12624 30308
rect 12023 30277 12035 30280
rect 11977 30271 12035 30277
rect 12618 30268 12624 30280
rect 12676 30268 12682 30320
rect 13280 30308 13308 30336
rect 14185 30311 14243 30317
rect 13280 30280 13860 30308
rect 3145 30249 3203 30255
rect 2961 30243 3019 30249
rect 2961 30209 2973 30243
rect 3007 30209 3019 30243
rect 2961 30203 3019 30209
rect 3053 30243 3111 30249
rect 3053 30209 3065 30243
rect 3099 30209 3111 30243
rect 3145 30215 3157 30249
rect 3191 30215 3203 30249
rect 3145 30209 3203 30215
rect 3053 30203 3111 30209
rect 2985 30104 3013 30203
rect 3326 30200 3332 30252
rect 3384 30240 3390 30252
rect 3384 30212 3429 30240
rect 3384 30200 3390 30212
rect 3878 30200 3884 30252
rect 3936 30240 3942 30252
rect 4065 30243 4123 30249
rect 4065 30240 4077 30243
rect 3936 30212 4077 30240
rect 3936 30200 3942 30212
rect 4065 30209 4077 30212
rect 4111 30209 4123 30243
rect 4065 30203 4123 30209
rect 4249 30243 4307 30249
rect 4249 30209 4261 30243
rect 4295 30209 4307 30243
rect 4249 30203 4307 30209
rect 4433 30243 4491 30249
rect 4433 30209 4445 30243
rect 4479 30240 4491 30243
rect 5074 30240 5080 30252
rect 4479 30212 5080 30240
rect 4479 30209 4491 30212
rect 4433 30203 4491 30209
rect 4264 30172 4292 30203
rect 5074 30200 5080 30212
rect 5132 30200 5138 30252
rect 5626 30200 5632 30252
rect 5684 30240 5690 30252
rect 5813 30243 5871 30249
rect 5813 30240 5825 30243
rect 5684 30212 5825 30240
rect 5684 30200 5690 30212
rect 5813 30209 5825 30212
rect 5859 30240 5871 30243
rect 6362 30240 6368 30252
rect 5859 30212 6368 30240
rect 5859 30209 5871 30212
rect 5813 30203 5871 30209
rect 6362 30200 6368 30212
rect 6420 30240 6426 30252
rect 6641 30243 6699 30249
rect 6641 30240 6653 30243
rect 6420 30212 6653 30240
rect 6420 30200 6426 30212
rect 6641 30209 6653 30212
rect 6687 30209 6699 30243
rect 6641 30203 6699 30209
rect 6733 30243 6791 30249
rect 6733 30209 6745 30243
rect 6779 30209 6791 30243
rect 6733 30203 6791 30209
rect 6825 30243 6883 30249
rect 6825 30209 6837 30243
rect 6871 30240 6883 30243
rect 6914 30240 6920 30252
rect 6871 30212 6920 30240
rect 6871 30209 6883 30212
rect 6825 30203 6883 30209
rect 4982 30172 4988 30184
rect 4264 30144 4988 30172
rect 4982 30132 4988 30144
rect 5040 30132 5046 30184
rect 6748 30172 6776 30203
rect 6914 30200 6920 30212
rect 6972 30200 6978 30252
rect 7009 30243 7067 30249
rect 7009 30209 7021 30243
rect 7055 30240 7067 30243
rect 7558 30240 7564 30252
rect 7055 30212 7564 30240
rect 7055 30209 7067 30212
rect 7009 30203 7067 30209
rect 7558 30200 7564 30212
rect 7616 30200 7622 30252
rect 9907 30243 9965 30249
rect 9907 30209 9919 30243
rect 9953 30209 9965 30243
rect 10042 30243 10100 30249
rect 10042 30240 10054 30243
rect 9907 30203 9965 30209
rect 10041 30209 10054 30240
rect 10088 30209 10100 30243
rect 10041 30203 10100 30209
rect 7466 30172 7472 30184
rect 6748 30144 7472 30172
rect 7466 30132 7472 30144
rect 7524 30132 7530 30184
rect 3418 30104 3424 30116
rect 2985 30076 3424 30104
rect 3418 30064 3424 30076
rect 3476 30104 3482 30116
rect 5077 30107 5135 30113
rect 5077 30104 5089 30107
rect 3476 30076 5089 30104
rect 3476 30064 3482 30076
rect 5077 30073 5089 30076
rect 5123 30073 5135 30107
rect 5077 30067 5135 30073
rect 9217 30107 9275 30113
rect 9217 30073 9229 30107
rect 9263 30104 9275 30107
rect 9922 30104 9950 30203
rect 10041 30172 10069 30203
rect 10134 30200 10140 30252
rect 10192 30249 10198 30252
rect 10192 30240 10200 30249
rect 10321 30243 10379 30249
rect 10192 30212 10237 30240
rect 10192 30203 10200 30212
rect 10321 30209 10333 30243
rect 10367 30209 10379 30243
rect 12158 30240 12164 30252
rect 12071 30212 12164 30240
rect 10321 30203 10379 30209
rect 10192 30200 10198 30203
rect 10041 30144 10088 30172
rect 10060 30116 10088 30144
rect 10226 30132 10232 30184
rect 10284 30172 10290 30184
rect 10336 30172 10364 30203
rect 12158 30200 12164 30212
rect 12216 30240 12222 30252
rect 12805 30243 12863 30249
rect 12805 30240 12817 30243
rect 12216 30212 12817 30240
rect 12216 30200 12222 30212
rect 12805 30209 12817 30212
rect 12851 30209 12863 30243
rect 12805 30203 12863 30209
rect 12986 30200 12992 30252
rect 13044 30240 13050 30252
rect 13044 30212 13137 30240
rect 13044 30200 13050 30212
rect 13170 30200 13176 30252
rect 13228 30240 13234 30252
rect 13541 30243 13599 30249
rect 13541 30240 13553 30243
rect 13228 30212 13553 30240
rect 13228 30200 13234 30212
rect 13541 30209 13553 30212
rect 13587 30209 13599 30243
rect 13722 30240 13728 30252
rect 13683 30212 13728 30240
rect 13541 30203 13599 30209
rect 13722 30200 13728 30212
rect 13780 30200 13786 30252
rect 13832 30249 13860 30280
rect 14185 30277 14197 30311
rect 14231 30308 14243 30311
rect 15194 30308 15200 30320
rect 14231 30280 15200 30308
rect 14231 30277 14243 30280
rect 14185 30271 14243 30277
rect 15194 30268 15200 30280
rect 15252 30268 15258 30320
rect 16758 30308 16764 30320
rect 16719 30280 16764 30308
rect 16758 30268 16764 30280
rect 16816 30268 16822 30320
rect 19705 30311 19763 30317
rect 19705 30277 19717 30311
rect 19751 30308 19763 30311
rect 20622 30308 20628 30320
rect 19751 30280 20628 30308
rect 19751 30277 19763 30280
rect 19705 30271 19763 30277
rect 20622 30268 20628 30280
rect 20680 30268 20686 30320
rect 22002 30268 22008 30320
rect 22060 30308 22066 30320
rect 22281 30311 22339 30317
rect 22281 30308 22293 30311
rect 22060 30280 22293 30308
rect 22060 30268 22066 30280
rect 22281 30277 22293 30280
rect 22327 30277 22339 30311
rect 22281 30271 22339 30277
rect 22373 30311 22431 30317
rect 22373 30277 22385 30311
rect 22419 30308 22431 30311
rect 25038 30308 25044 30320
rect 22419 30280 25044 30308
rect 22419 30277 22431 30280
rect 22373 30271 22431 30277
rect 25038 30268 25044 30280
rect 25096 30268 25102 30320
rect 26050 30268 26056 30320
rect 26108 30308 26114 30320
rect 28368 30308 28396 30339
rect 30926 30336 30932 30348
rect 30984 30336 30990 30388
rect 31202 30376 31208 30388
rect 31163 30348 31208 30376
rect 31202 30336 31208 30348
rect 31260 30336 31266 30388
rect 28626 30308 28632 30320
rect 26108 30280 28396 30308
rect 28587 30280 28632 30308
rect 26108 30268 26114 30280
rect 28626 30268 28632 30280
rect 28684 30268 28690 30320
rect 28718 30268 28724 30320
rect 28776 30308 28782 30320
rect 28776 30280 29960 30308
rect 28776 30268 28782 30280
rect 29932 30252 29960 30280
rect 30374 30268 30380 30320
rect 30432 30308 30438 30320
rect 31389 30311 31447 30317
rect 30432 30280 30788 30308
rect 30432 30268 30438 30280
rect 13817 30243 13875 30249
rect 13817 30209 13829 30243
rect 13863 30209 13875 30243
rect 13817 30203 13875 30209
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30240 13967 30243
rect 13955 30212 14780 30240
rect 13955 30209 13967 30212
rect 13909 30203 13967 30209
rect 10284 30144 10364 30172
rect 12345 30175 12403 30181
rect 10284 30132 10290 30144
rect 12345 30141 12357 30175
rect 12391 30172 12403 30175
rect 12434 30172 12440 30184
rect 12391 30144 12440 30172
rect 12391 30141 12403 30144
rect 12345 30135 12403 30141
rect 12434 30132 12440 30144
rect 12492 30132 12498 30184
rect 13004 30172 13032 30200
rect 13446 30172 13452 30184
rect 13004 30144 13452 30172
rect 13446 30132 13452 30144
rect 13504 30132 13510 30184
rect 9263 30076 9950 30104
rect 9263 30073 9275 30076
rect 9217 30067 9275 30073
rect 4617 30039 4675 30045
rect 4617 30005 4629 30039
rect 4663 30036 4675 30039
rect 4798 30036 4804 30048
rect 4663 30008 4804 30036
rect 4663 30005 4675 30008
rect 4617 29999 4675 30005
rect 4798 29996 4804 30008
rect 4856 29996 4862 30048
rect 7558 30036 7564 30048
rect 7519 30008 7564 30036
rect 7558 29996 7564 30008
rect 7616 29996 7622 30048
rect 9490 29996 9496 30048
rect 9548 30036 9554 30048
rect 9677 30039 9735 30045
rect 9677 30036 9689 30039
rect 9548 30008 9689 30036
rect 9548 29996 9554 30008
rect 9677 30005 9689 30008
rect 9723 30005 9735 30039
rect 9922 30036 9950 30076
rect 10042 30064 10048 30116
rect 10100 30064 10106 30116
rect 10778 30064 10784 30116
rect 10836 30104 10842 30116
rect 14366 30104 14372 30116
rect 10836 30076 14372 30104
rect 10836 30064 10842 30076
rect 14366 30064 14372 30076
rect 14424 30064 14430 30116
rect 12894 30036 12900 30048
rect 9922 30008 12900 30036
rect 9677 29999 9735 30005
rect 12894 29996 12900 30008
rect 12952 29996 12958 30048
rect 14752 30045 14780 30212
rect 15286 30200 15292 30252
rect 15344 30240 15350 30252
rect 16942 30240 16948 30252
rect 15344 30212 16948 30240
rect 15344 30200 15350 30212
rect 16942 30200 16948 30212
rect 17000 30200 17006 30252
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 19426 30240 19432 30252
rect 19107 30212 19432 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 19426 30200 19432 30212
rect 19484 30240 19490 30252
rect 19886 30240 19892 30252
rect 19484 30212 19892 30240
rect 19484 30200 19490 30212
rect 19886 30200 19892 30212
rect 19944 30200 19950 30252
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 22465 30243 22523 30249
rect 22152 30212 22197 30240
rect 22152 30200 22158 30212
rect 22465 30209 22477 30243
rect 22511 30240 22523 30243
rect 23106 30240 23112 30252
rect 22511 30212 23112 30240
rect 22511 30209 22523 30212
rect 22465 30203 22523 30209
rect 16666 30132 16672 30184
rect 16724 30172 16730 30184
rect 17129 30175 17187 30181
rect 17129 30172 17141 30175
rect 16724 30144 17141 30172
rect 16724 30132 16730 30144
rect 17129 30141 17141 30144
rect 17175 30141 17187 30175
rect 17129 30135 17187 30141
rect 17144 30104 17172 30135
rect 20898 30132 20904 30184
rect 20956 30172 20962 30184
rect 22480 30172 22508 30203
rect 23106 30200 23112 30212
rect 23164 30200 23170 30252
rect 24854 30200 24860 30252
rect 24912 30240 24918 30252
rect 24949 30243 25007 30249
rect 24949 30240 24961 30243
rect 24912 30212 24961 30240
rect 24912 30200 24918 30212
rect 24949 30209 24961 30212
rect 24995 30209 25007 30243
rect 28534 30240 28540 30252
rect 28447 30212 28540 30240
rect 24949 30203 25007 30209
rect 28534 30200 28540 30212
rect 28592 30240 28598 30252
rect 28592 30212 28764 30240
rect 28592 30200 28598 30212
rect 20956 30144 22508 30172
rect 20956 30132 20962 30144
rect 24578 30132 24584 30184
rect 24636 30172 24642 30184
rect 24673 30175 24731 30181
rect 24673 30172 24685 30175
rect 24636 30144 24685 30172
rect 24636 30132 24642 30144
rect 24673 30141 24685 30144
rect 24719 30141 24731 30175
rect 24673 30135 24731 30141
rect 28736 30104 28764 30212
rect 28810 30200 28816 30252
rect 28868 30240 28874 30252
rect 28905 30243 28963 30249
rect 28905 30240 28917 30243
rect 28868 30212 28917 30240
rect 28868 30200 28874 30212
rect 28905 30209 28917 30212
rect 28951 30209 28963 30243
rect 29914 30240 29920 30252
rect 29875 30212 29920 30240
rect 28905 30203 28963 30209
rect 29914 30200 29920 30212
rect 29972 30240 29978 30252
rect 30760 30249 30788 30280
rect 31389 30277 31401 30311
rect 31435 30308 31447 30311
rect 32950 30308 32956 30320
rect 31435 30280 32956 30308
rect 31435 30277 31447 30280
rect 31389 30271 31447 30277
rect 32950 30268 32956 30280
rect 33008 30268 33014 30320
rect 33686 30308 33692 30320
rect 33647 30280 33692 30308
rect 33686 30268 33692 30280
rect 33744 30308 33750 30320
rect 34238 30308 34244 30320
rect 33744 30280 34244 30308
rect 33744 30268 33750 30280
rect 34238 30268 34244 30280
rect 34296 30308 34302 30320
rect 34793 30311 34851 30317
rect 34296 30280 34560 30308
rect 34296 30268 34302 30280
rect 30561 30243 30619 30249
rect 30561 30240 30573 30243
rect 29972 30212 30573 30240
rect 29972 30200 29978 30212
rect 30561 30209 30573 30212
rect 30607 30209 30619 30243
rect 30561 30203 30619 30209
rect 30745 30243 30803 30249
rect 30745 30209 30757 30243
rect 30791 30209 30803 30243
rect 31570 30240 31576 30252
rect 31483 30212 31576 30240
rect 30745 30203 30803 30209
rect 31570 30200 31576 30212
rect 31628 30200 31634 30252
rect 32674 30240 32680 30252
rect 32635 30212 32680 30240
rect 32674 30200 32680 30212
rect 32732 30200 32738 30252
rect 33594 30200 33600 30252
rect 33652 30240 33658 30252
rect 34149 30243 34207 30249
rect 34149 30240 34161 30243
rect 33652 30212 34161 30240
rect 33652 30200 33658 30212
rect 34149 30209 34161 30212
rect 34195 30209 34207 30243
rect 34330 30240 34336 30252
rect 34291 30212 34336 30240
rect 34149 30203 34207 30209
rect 34330 30200 34336 30212
rect 34388 30200 34394 30252
rect 34532 30249 34560 30280
rect 34793 30277 34805 30311
rect 34839 30308 34851 30311
rect 35894 30308 35900 30320
rect 34839 30280 35900 30308
rect 34839 30277 34851 30280
rect 34793 30271 34851 30277
rect 35894 30268 35900 30280
rect 35952 30268 35958 30320
rect 34425 30243 34483 30249
rect 34425 30209 34437 30243
rect 34471 30209 34483 30243
rect 34425 30203 34483 30209
rect 34517 30243 34575 30249
rect 34517 30209 34529 30243
rect 34563 30209 34575 30243
rect 34517 30203 34575 30209
rect 35529 30243 35587 30249
rect 35529 30209 35541 30243
rect 35575 30240 35587 30243
rect 35986 30240 35992 30252
rect 35575 30212 35992 30240
rect 35575 30209 35587 30212
rect 35529 30203 35587 30209
rect 29733 30175 29791 30181
rect 29733 30141 29745 30175
rect 29779 30172 29791 30175
rect 30101 30175 30159 30181
rect 29779 30144 29960 30172
rect 29779 30141 29791 30144
rect 29733 30135 29791 30141
rect 29822 30104 29828 30116
rect 17144 30076 24532 30104
rect 14737 30039 14795 30045
rect 14737 30005 14749 30039
rect 14783 30036 14795 30039
rect 14826 30036 14832 30048
rect 14783 30008 14832 30036
rect 14783 30005 14795 30008
rect 14737 29999 14795 30005
rect 14826 29996 14832 30008
rect 14884 29996 14890 30048
rect 19426 29996 19432 30048
rect 19484 30036 19490 30048
rect 19521 30039 19579 30045
rect 19521 30036 19533 30039
rect 19484 30008 19533 30036
rect 19484 29996 19490 30008
rect 19521 30005 19533 30008
rect 19567 30005 19579 30039
rect 22646 30036 22652 30048
rect 22607 30008 22652 30036
rect 19521 29999 19579 30005
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 24504 30036 24532 30076
rect 28184 30076 28672 30104
rect 28736 30076 29828 30104
rect 28184 30036 28212 30076
rect 24504 30008 28212 30036
rect 28644 30036 28672 30076
rect 29822 30064 29828 30076
rect 29880 30064 29886 30116
rect 29546 30036 29552 30048
rect 28644 30008 29552 30036
rect 29546 29996 29552 30008
rect 29604 30036 29610 30048
rect 29932 30036 29960 30144
rect 30101 30141 30113 30175
rect 30147 30172 30159 30175
rect 31588 30172 31616 30200
rect 30147 30144 31616 30172
rect 32953 30175 33011 30181
rect 30147 30141 30159 30144
rect 30101 30135 30159 30141
rect 32953 30141 32965 30175
rect 32999 30172 33011 30175
rect 33042 30172 33048 30184
rect 32999 30144 33048 30172
rect 32999 30141 33011 30144
rect 32953 30135 33011 30141
rect 33042 30132 33048 30144
rect 33100 30132 33106 30184
rect 30926 30064 30932 30116
rect 30984 30104 30990 30116
rect 34440 30104 34468 30203
rect 35986 30200 35992 30212
rect 36044 30240 36050 30252
rect 36446 30240 36452 30252
rect 36044 30212 36452 30240
rect 36044 30200 36050 30212
rect 36446 30200 36452 30212
rect 36504 30200 36510 30252
rect 37277 30243 37335 30249
rect 37277 30209 37289 30243
rect 37323 30209 37335 30243
rect 37458 30240 37464 30252
rect 37419 30212 37464 30240
rect 37277 30203 37335 30209
rect 35253 30175 35311 30181
rect 35253 30172 35265 30175
rect 30984 30076 34468 30104
rect 34532 30144 35265 30172
rect 30984 30064 30990 30076
rect 29604 30008 29960 30036
rect 29604 29996 29610 30008
rect 31754 29996 31760 30048
rect 31812 30036 31818 30048
rect 34532 30036 34560 30144
rect 35253 30141 35265 30144
rect 35299 30141 35311 30175
rect 35253 30135 35311 30141
rect 35342 30132 35348 30184
rect 35400 30172 35406 30184
rect 37292 30172 37320 30203
rect 37458 30200 37464 30212
rect 37516 30200 37522 30252
rect 35400 30144 37320 30172
rect 35400 30132 35406 30144
rect 31812 30008 34560 30036
rect 31812 29996 31818 30008
rect 35710 29996 35716 30048
rect 35768 30036 35774 30048
rect 37645 30039 37703 30045
rect 37645 30036 37657 30039
rect 35768 30008 37657 30036
rect 35768 29996 35774 30008
rect 37645 30005 37657 30008
rect 37691 30005 37703 30039
rect 37645 29999 37703 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 3234 29832 3240 29844
rect 3195 29804 3240 29832
rect 3234 29792 3240 29804
rect 3292 29792 3298 29844
rect 6914 29832 6920 29844
rect 6875 29804 6920 29832
rect 6914 29792 6920 29804
rect 6972 29792 6978 29844
rect 7576 29804 12434 29832
rect 4614 29764 4620 29776
rect 2985 29736 4620 29764
rect 2774 29588 2780 29640
rect 2832 29628 2838 29640
rect 2869 29631 2927 29637
rect 2869 29628 2881 29631
rect 2832 29600 2881 29628
rect 2832 29588 2838 29600
rect 2869 29597 2881 29600
rect 2915 29628 2927 29631
rect 2985 29628 3013 29736
rect 4614 29724 4620 29736
rect 4672 29724 4678 29776
rect 3142 29656 3148 29708
rect 3200 29696 3206 29708
rect 3200 29668 4384 29696
rect 3200 29656 3206 29668
rect 2915 29600 3013 29628
rect 3053 29631 3111 29637
rect 2915 29597 2927 29600
rect 2869 29591 2927 29597
rect 3053 29597 3065 29631
rect 3099 29628 3111 29631
rect 3510 29628 3516 29640
rect 3099 29600 3516 29628
rect 3099 29597 3111 29600
rect 3053 29591 3111 29597
rect 3510 29588 3516 29600
rect 3568 29628 3574 29640
rect 4356 29637 4384 29668
rect 4065 29631 4123 29637
rect 4065 29628 4077 29631
rect 3568 29600 4077 29628
rect 3568 29588 3574 29600
rect 4065 29597 4077 29600
rect 4111 29597 4123 29631
rect 4065 29591 4123 29597
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29597 4399 29631
rect 4341 29591 4399 29597
rect 4433 29631 4491 29637
rect 4433 29597 4445 29631
rect 4479 29628 4491 29631
rect 5074 29628 5080 29640
rect 4479 29600 5080 29628
rect 4479 29597 4491 29600
rect 4433 29591 4491 29597
rect 5074 29588 5080 29600
rect 5132 29588 5138 29640
rect 6733 29631 6791 29637
rect 6733 29597 6745 29631
rect 6779 29628 6791 29631
rect 7098 29628 7104 29640
rect 6779 29600 7104 29628
rect 6779 29597 6791 29600
rect 6733 29591 6791 29597
rect 7098 29588 7104 29600
rect 7156 29588 7162 29640
rect 7576 29637 7604 29804
rect 12406 29764 12434 29804
rect 13170 29792 13176 29844
rect 13228 29832 13234 29844
rect 13449 29835 13507 29841
rect 13449 29832 13461 29835
rect 13228 29804 13461 29832
rect 13228 29792 13234 29804
rect 13449 29801 13461 29804
rect 13495 29801 13507 29835
rect 13449 29795 13507 29801
rect 19889 29835 19947 29841
rect 19889 29801 19901 29835
rect 19935 29832 19947 29835
rect 19978 29832 19984 29844
rect 19935 29804 19984 29832
rect 19935 29801 19947 29804
rect 19889 29795 19947 29801
rect 19978 29792 19984 29804
rect 20036 29792 20042 29844
rect 29546 29832 29552 29844
rect 20088 29804 22094 29832
rect 15010 29764 15016 29776
rect 12406 29736 15016 29764
rect 15010 29724 15016 29736
rect 15068 29724 15074 29776
rect 15746 29724 15752 29776
rect 15804 29764 15810 29776
rect 20088 29764 20116 29804
rect 15804 29736 20116 29764
rect 20809 29767 20867 29773
rect 15804 29724 15810 29736
rect 20809 29733 20821 29767
rect 20855 29764 20867 29767
rect 21174 29764 21180 29776
rect 20855 29736 21180 29764
rect 20855 29733 20867 29736
rect 20809 29727 20867 29733
rect 21174 29724 21180 29736
rect 21232 29724 21238 29776
rect 21818 29724 21824 29776
rect 21876 29764 21882 29776
rect 21913 29767 21971 29773
rect 21913 29764 21925 29767
rect 21876 29736 21925 29764
rect 21876 29724 21882 29736
rect 21913 29733 21925 29736
rect 21959 29733 21971 29767
rect 21913 29727 21971 29733
rect 8938 29656 8944 29708
rect 8996 29696 9002 29708
rect 9217 29699 9275 29705
rect 9217 29696 9229 29699
rect 8996 29668 9229 29696
rect 8996 29656 9002 29668
rect 9217 29665 9229 29668
rect 9263 29665 9275 29699
rect 9217 29659 9275 29665
rect 11333 29699 11391 29705
rect 11333 29665 11345 29699
rect 11379 29696 11391 29699
rect 12526 29696 12532 29708
rect 11379 29668 12532 29696
rect 11379 29665 11391 29668
rect 11333 29659 11391 29665
rect 12526 29656 12532 29668
rect 12584 29656 12590 29708
rect 12894 29656 12900 29708
rect 12952 29696 12958 29708
rect 18049 29699 18107 29705
rect 18049 29696 18061 29699
rect 12952 29668 18061 29696
rect 12952 29656 12958 29668
rect 18049 29665 18061 29668
rect 18095 29696 18107 29699
rect 18095 29668 19656 29696
rect 18095 29665 18107 29668
rect 18049 29659 18107 29665
rect 9490 29637 9496 29640
rect 7561 29631 7619 29637
rect 7561 29597 7573 29631
rect 7607 29597 7619 29631
rect 9484 29628 9496 29637
rect 9451 29600 9496 29628
rect 7561 29591 7619 29597
rect 9484 29591 9496 29600
rect 9490 29588 9496 29591
rect 9548 29588 9554 29640
rect 11057 29631 11115 29637
rect 11057 29597 11069 29631
rect 11103 29628 11115 29631
rect 11146 29628 11152 29640
rect 11103 29600 11152 29628
rect 11103 29597 11115 29600
rect 11057 29591 11115 29597
rect 11146 29588 11152 29600
rect 11204 29588 11210 29640
rect 12437 29631 12495 29637
rect 12437 29597 12449 29631
rect 12483 29597 12495 29631
rect 12544 29628 12572 29656
rect 12621 29631 12679 29637
rect 12621 29628 12633 29631
rect 12544 29600 12633 29628
rect 12437 29591 12495 29597
rect 12621 29597 12633 29600
rect 12667 29597 12679 29631
rect 12802 29628 12808 29640
rect 12763 29600 12808 29628
rect 12621 29591 12679 29597
rect 4249 29563 4307 29569
rect 4249 29529 4261 29563
rect 4295 29560 4307 29563
rect 4982 29560 4988 29572
rect 4295 29532 4988 29560
rect 4295 29529 4307 29532
rect 4249 29523 4307 29529
rect 4982 29520 4988 29532
rect 5040 29520 5046 29572
rect 6549 29563 6607 29569
rect 6549 29529 6561 29563
rect 6595 29560 6607 29563
rect 7006 29560 7012 29572
rect 6595 29532 7012 29560
rect 6595 29529 6607 29532
rect 6549 29523 6607 29529
rect 7006 29520 7012 29532
rect 7064 29560 7070 29572
rect 7064 29532 7420 29560
rect 7064 29520 7070 29532
rect 4617 29495 4675 29501
rect 4617 29461 4629 29495
rect 4663 29492 4675 29495
rect 4706 29492 4712 29504
rect 4663 29464 4712 29492
rect 4663 29461 4675 29464
rect 4617 29455 4675 29461
rect 4706 29452 4712 29464
rect 4764 29452 4770 29504
rect 7392 29501 7420 29532
rect 7377 29495 7435 29501
rect 7377 29461 7389 29495
rect 7423 29461 7435 29495
rect 7377 29455 7435 29461
rect 9950 29452 9956 29504
rect 10008 29492 10014 29504
rect 10597 29495 10655 29501
rect 10597 29492 10609 29495
rect 10008 29464 10609 29492
rect 10008 29452 10014 29464
rect 10597 29461 10609 29464
rect 10643 29492 10655 29495
rect 12452 29492 12480 29591
rect 12802 29588 12808 29600
rect 12860 29588 12866 29640
rect 15749 29631 15807 29637
rect 15749 29597 15761 29631
rect 15795 29628 15807 29631
rect 16758 29628 16764 29640
rect 15795 29600 16764 29628
rect 15795 29597 15807 29600
rect 15749 29591 15807 29597
rect 16758 29588 16764 29600
rect 16816 29588 16822 29640
rect 17586 29588 17592 29640
rect 17644 29628 17650 29640
rect 19245 29631 19303 29637
rect 19245 29628 19257 29631
rect 17644 29600 19257 29628
rect 17644 29588 17650 29600
rect 19245 29597 19257 29600
rect 19291 29597 19303 29631
rect 19426 29628 19432 29640
rect 19387 29600 19432 29628
rect 19245 29591 19303 29597
rect 19426 29588 19432 29600
rect 19484 29588 19490 29640
rect 19628 29637 19656 29668
rect 20622 29656 20628 29708
rect 20680 29696 20686 29708
rect 22066 29696 22094 29804
rect 25148 29804 27292 29832
rect 29507 29804 29552 29832
rect 23845 29699 23903 29705
rect 23845 29696 23857 29699
rect 20680 29668 21404 29696
rect 22066 29668 23857 29696
rect 20680 29656 20686 29668
rect 19521 29631 19579 29637
rect 19521 29597 19533 29631
rect 19567 29597 19579 29631
rect 19521 29591 19579 29597
rect 19613 29631 19671 29637
rect 19613 29597 19625 29631
rect 19659 29597 19671 29631
rect 19613 29591 19671 29597
rect 12713 29563 12771 29569
rect 12713 29529 12725 29563
rect 12759 29560 12771 29563
rect 13354 29560 13360 29572
rect 12759 29532 13360 29560
rect 12759 29529 12771 29532
rect 12713 29523 12771 29529
rect 13354 29520 13360 29532
rect 13412 29520 13418 29572
rect 15930 29560 15936 29572
rect 15891 29532 15936 29560
rect 15930 29520 15936 29532
rect 15988 29520 15994 29572
rect 19334 29560 19340 29572
rect 18616 29532 19340 29560
rect 10643 29464 12480 29492
rect 12989 29495 13047 29501
rect 10643 29461 10655 29464
rect 10597 29455 10655 29461
rect 12989 29461 13001 29495
rect 13035 29492 13047 29495
rect 14734 29492 14740 29504
rect 13035 29464 14740 29492
rect 13035 29461 13047 29464
rect 12989 29455 13047 29461
rect 14734 29452 14740 29464
rect 14792 29452 14798 29504
rect 16022 29452 16028 29504
rect 16080 29492 16086 29504
rect 16117 29495 16175 29501
rect 16117 29492 16129 29495
rect 16080 29464 16129 29492
rect 16080 29452 16086 29464
rect 16117 29461 16129 29464
rect 16163 29461 16175 29495
rect 16666 29492 16672 29504
rect 16627 29464 16672 29492
rect 16117 29455 16175 29461
rect 16666 29452 16672 29464
rect 16724 29452 16730 29504
rect 18414 29452 18420 29504
rect 18472 29492 18478 29504
rect 18616 29501 18644 29532
rect 19334 29520 19340 29532
rect 19392 29560 19398 29572
rect 19536 29560 19564 29591
rect 20898 29588 20904 29640
rect 20956 29628 20962 29640
rect 21376 29637 21404 29668
rect 23845 29665 23857 29668
rect 23891 29696 23903 29699
rect 25148 29696 25176 29804
rect 27264 29764 27292 29804
rect 29546 29792 29552 29804
rect 29604 29792 29610 29844
rect 32950 29832 32956 29844
rect 32911 29804 32956 29832
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 31478 29764 31484 29776
rect 27264 29736 31484 29764
rect 31478 29724 31484 29736
rect 31536 29724 31542 29776
rect 35986 29696 35992 29708
rect 23891 29668 25176 29696
rect 23891 29665 23903 29668
rect 23845 29659 23903 29665
rect 20993 29631 21051 29637
rect 20993 29628 21005 29631
rect 20956 29600 21005 29628
rect 20956 29588 20962 29600
rect 20993 29597 21005 29600
rect 21039 29597 21051 29631
rect 20993 29591 21051 29597
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29597 21419 29631
rect 21361 29591 21419 29597
rect 21450 29588 21456 29640
rect 21508 29628 21514 29640
rect 21508 29600 22968 29628
rect 21508 29588 21514 29600
rect 21082 29560 21088 29572
rect 19392 29532 19564 29560
rect 21043 29532 21088 29560
rect 19392 29520 19398 29532
rect 21082 29520 21088 29532
rect 21140 29520 21146 29572
rect 21177 29563 21235 29569
rect 21177 29529 21189 29563
rect 21223 29560 21235 29563
rect 22002 29560 22008 29572
rect 21223 29532 22008 29560
rect 21223 29529 21235 29532
rect 21177 29523 21235 29529
rect 18601 29495 18659 29501
rect 18601 29492 18613 29495
rect 18472 29464 18613 29492
rect 18472 29452 18478 29464
rect 18601 29461 18613 29464
rect 18647 29461 18659 29495
rect 18601 29455 18659 29461
rect 20714 29452 20720 29504
rect 20772 29492 20778 29504
rect 21192 29492 21220 29523
rect 22002 29520 22008 29532
rect 22060 29560 22066 29572
rect 22833 29563 22891 29569
rect 22833 29560 22845 29563
rect 22060 29532 22845 29560
rect 22060 29520 22066 29532
rect 22833 29529 22845 29532
rect 22879 29529 22891 29563
rect 22940 29560 22968 29600
rect 24486 29588 24492 29640
rect 24544 29628 24550 29640
rect 24765 29631 24823 29637
rect 24765 29628 24777 29631
rect 24544 29600 24777 29628
rect 24544 29588 24550 29600
rect 24765 29597 24777 29600
rect 24811 29597 24823 29631
rect 24946 29628 24952 29640
rect 24907 29600 24952 29628
rect 24765 29591 24823 29597
rect 24946 29588 24952 29600
rect 25004 29588 25010 29640
rect 25148 29637 25176 29668
rect 35820 29668 35992 29696
rect 25041 29631 25099 29637
rect 25041 29597 25053 29631
rect 25087 29597 25099 29631
rect 25041 29591 25099 29597
rect 25133 29631 25191 29637
rect 25133 29597 25145 29631
rect 25179 29597 25191 29631
rect 27249 29631 27307 29637
rect 27249 29628 27261 29631
rect 25133 29591 25191 29597
rect 26804 29600 27261 29628
rect 24578 29560 24584 29572
rect 22940 29532 24584 29560
rect 22833 29523 22891 29529
rect 24578 29520 24584 29532
rect 24636 29560 24642 29572
rect 25056 29560 25084 29591
rect 26804 29572 26832 29600
rect 27249 29597 27261 29600
rect 27295 29597 27307 29631
rect 31570 29628 31576 29640
rect 31531 29600 31576 29628
rect 27249 29591 27307 29597
rect 31570 29588 31576 29600
rect 31628 29588 31634 29640
rect 31846 29637 31852 29640
rect 31840 29591 31852 29637
rect 31904 29628 31910 29640
rect 31904 29600 31940 29628
rect 31846 29588 31852 29591
rect 31904 29588 31910 29600
rect 35434 29588 35440 29640
rect 35492 29628 35498 29640
rect 35529 29631 35587 29637
rect 35529 29628 35541 29631
rect 35492 29600 35541 29628
rect 35492 29588 35498 29600
rect 35529 29597 35541 29600
rect 35575 29597 35587 29631
rect 35710 29628 35716 29640
rect 35671 29600 35716 29628
rect 35529 29591 35587 29597
rect 35710 29588 35716 29600
rect 35768 29588 35774 29640
rect 35820 29637 35848 29668
rect 35986 29656 35992 29668
rect 36044 29656 36050 29708
rect 35805 29631 35863 29637
rect 35805 29597 35817 29631
rect 35851 29597 35863 29631
rect 35805 29591 35863 29597
rect 35894 29588 35900 29640
rect 35952 29628 35958 29640
rect 35952 29600 35997 29628
rect 35952 29588 35958 29600
rect 38562 29588 38568 29640
rect 38620 29628 38626 29640
rect 38657 29631 38715 29637
rect 38657 29628 38669 29631
rect 38620 29600 38669 29628
rect 38620 29588 38626 29600
rect 38657 29597 38669 29600
rect 38703 29597 38715 29631
rect 58158 29628 58164 29640
rect 58119 29600 58164 29628
rect 38657 29591 38715 29597
rect 58158 29588 58164 29600
rect 58216 29588 58222 29640
rect 24636 29532 25084 29560
rect 25409 29563 25467 29569
rect 24636 29520 24642 29532
rect 25409 29529 25421 29563
rect 25455 29560 25467 29563
rect 25455 29532 26740 29560
rect 25455 29529 25467 29532
rect 25409 29523 25467 29529
rect 20772 29464 21220 29492
rect 20772 29452 20778 29464
rect 22462 29452 22468 29504
rect 22520 29492 22526 29504
rect 22925 29495 22983 29501
rect 22925 29492 22937 29495
rect 22520 29464 22937 29492
rect 22520 29452 22526 29464
rect 22925 29461 22937 29464
rect 22971 29461 22983 29495
rect 25866 29492 25872 29504
rect 25827 29464 25872 29492
rect 22925 29455 22983 29461
rect 25866 29452 25872 29464
rect 25924 29452 25930 29504
rect 26712 29492 26740 29532
rect 26786 29520 26792 29572
rect 26844 29520 26850 29572
rect 26982 29563 27040 29569
rect 26982 29560 26994 29563
rect 26896 29532 26994 29560
rect 26896 29492 26924 29532
rect 26982 29529 26994 29532
rect 27028 29529 27040 29563
rect 26982 29523 27040 29529
rect 33870 29520 33876 29572
rect 33928 29560 33934 29572
rect 36173 29563 36231 29569
rect 33928 29532 36124 29560
rect 33928 29520 33934 29532
rect 30374 29492 30380 29504
rect 26712 29464 26924 29492
rect 30335 29464 30380 29492
rect 30374 29452 30380 29464
rect 30432 29452 30438 29504
rect 34606 29452 34612 29504
rect 34664 29492 34670 29504
rect 34977 29495 35035 29501
rect 34977 29492 34989 29495
rect 34664 29464 34989 29492
rect 34664 29452 34670 29464
rect 34977 29461 34989 29464
rect 35023 29492 35035 29495
rect 35526 29492 35532 29504
rect 35023 29464 35532 29492
rect 35023 29461 35035 29464
rect 34977 29455 35035 29461
rect 35526 29452 35532 29464
rect 35584 29492 35590 29504
rect 35802 29492 35808 29504
rect 35584 29464 35808 29492
rect 35584 29452 35590 29464
rect 35802 29452 35808 29464
rect 35860 29452 35866 29504
rect 36096 29492 36124 29532
rect 36173 29529 36185 29563
rect 36219 29560 36231 29563
rect 38390 29563 38448 29569
rect 38390 29560 38402 29563
rect 36219 29532 38402 29560
rect 36219 29529 36231 29532
rect 36173 29523 36231 29529
rect 38390 29529 38402 29532
rect 38436 29529 38448 29563
rect 38390 29523 38448 29529
rect 37277 29495 37335 29501
rect 37277 29492 37289 29495
rect 36096 29464 37289 29492
rect 37277 29461 37289 29464
rect 37323 29492 37335 29495
rect 37458 29492 37464 29504
rect 37323 29464 37464 29492
rect 37323 29461 37335 29464
rect 37277 29455 37335 29461
rect 37458 29452 37464 29464
rect 37516 29452 37522 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 19153 29291 19211 29297
rect 19153 29257 19165 29291
rect 19199 29257 19211 29291
rect 19153 29251 19211 29257
rect 17126 29220 17132 29232
rect 15856 29192 17132 29220
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29152 9551 29155
rect 11698 29152 11704 29164
rect 9539 29124 11704 29152
rect 9539 29121 9551 29124
rect 9493 29115 9551 29121
rect 11698 29112 11704 29124
rect 11756 29112 11762 29164
rect 11885 29155 11943 29161
rect 11885 29121 11897 29155
rect 11931 29152 11943 29155
rect 12802 29152 12808 29164
rect 11931 29124 12808 29152
rect 11931 29121 11943 29124
rect 11885 29115 11943 29121
rect 12802 29112 12808 29124
rect 12860 29112 12866 29164
rect 14642 29112 14648 29164
rect 14700 29152 14706 29164
rect 14826 29152 14832 29164
rect 14700 29124 14832 29152
rect 14700 29112 14706 29124
rect 14826 29112 14832 29124
rect 14884 29152 14890 29164
rect 15013 29155 15071 29161
rect 15013 29152 15025 29155
rect 14884 29124 15025 29152
rect 14884 29112 14890 29124
rect 15013 29121 15025 29124
rect 15059 29152 15071 29155
rect 15746 29152 15752 29164
rect 15059 29124 15752 29152
rect 15059 29121 15071 29124
rect 15013 29115 15071 29121
rect 15746 29112 15752 29124
rect 15804 29112 15810 29164
rect 15856 29161 15884 29192
rect 17126 29180 17132 29192
rect 17184 29180 17190 29232
rect 17310 29180 17316 29232
rect 17368 29220 17374 29232
rect 18138 29220 18144 29232
rect 17368 29192 18144 29220
rect 17368 29180 17374 29192
rect 18138 29180 18144 29192
rect 18196 29180 18202 29232
rect 19168 29220 19196 29251
rect 24946 29248 24952 29300
rect 25004 29288 25010 29300
rect 25133 29291 25191 29297
rect 25133 29288 25145 29291
rect 25004 29260 25145 29288
rect 25004 29248 25010 29260
rect 25133 29257 25145 29260
rect 25179 29257 25191 29291
rect 25133 29251 25191 29257
rect 30009 29291 30067 29297
rect 30009 29257 30021 29291
rect 30055 29288 30067 29291
rect 31754 29288 31760 29300
rect 30055 29260 31760 29288
rect 30055 29257 30067 29260
rect 30009 29251 30067 29257
rect 31754 29248 31760 29260
rect 31812 29248 31818 29300
rect 34790 29248 34796 29300
rect 34848 29288 34854 29300
rect 34885 29291 34943 29297
rect 34885 29288 34897 29291
rect 34848 29260 34897 29288
rect 34848 29248 34854 29260
rect 34885 29257 34897 29260
rect 34931 29257 34943 29291
rect 34885 29251 34943 29257
rect 19797 29223 19855 29229
rect 19797 29220 19809 29223
rect 19168 29192 19809 29220
rect 19797 29189 19809 29192
rect 19843 29220 19855 29223
rect 20622 29220 20628 29232
rect 19843 29192 20484 29220
rect 20583 29192 20628 29220
rect 19843 29189 19855 29192
rect 19797 29183 19855 29189
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29121 15899 29155
rect 15841 29115 15899 29121
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29152 15991 29155
rect 16022 29152 16028 29164
rect 15979 29124 16028 29152
rect 15979 29121 15991 29124
rect 15933 29115 15991 29121
rect 7466 29044 7472 29096
rect 7524 29084 7530 29096
rect 9217 29087 9275 29093
rect 9217 29084 9229 29087
rect 7524 29056 9229 29084
rect 7524 29044 7530 29056
rect 9217 29053 9229 29056
rect 9263 29053 9275 29087
rect 9217 29047 9275 29053
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 10689 29087 10747 29093
rect 10689 29084 10701 29087
rect 9732 29056 10701 29084
rect 9732 29044 9738 29056
rect 10689 29053 10701 29056
rect 10735 29053 10747 29087
rect 10689 29047 10747 29053
rect 10965 29087 11023 29093
rect 10965 29053 10977 29087
rect 11011 29053 11023 29087
rect 10965 29047 11023 29053
rect 10980 29016 11008 29047
rect 11422 29044 11428 29096
rect 11480 29084 11486 29096
rect 11609 29087 11667 29093
rect 11609 29084 11621 29087
rect 11480 29056 11621 29084
rect 11480 29044 11486 29056
rect 11609 29053 11621 29056
rect 11655 29053 11667 29087
rect 11609 29047 11667 29053
rect 15102 29044 15108 29096
rect 15160 29084 15166 29096
rect 15856 29084 15884 29115
rect 16022 29112 16028 29124
rect 16080 29112 16086 29164
rect 16114 29112 16120 29164
rect 16172 29152 16178 29164
rect 17770 29152 17776 29164
rect 16172 29124 16217 29152
rect 17731 29124 17776 29152
rect 16172 29112 16178 29124
rect 17770 29112 17776 29124
rect 17828 29112 17834 29164
rect 17862 29112 17868 29164
rect 17920 29152 17926 29164
rect 18029 29155 18087 29161
rect 18029 29152 18041 29155
rect 17920 29124 18041 29152
rect 17920 29112 17926 29124
rect 18029 29121 18041 29124
rect 18075 29121 18087 29155
rect 19978 29152 19984 29164
rect 19939 29124 19984 29152
rect 18029 29115 18087 29121
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 20456 29161 20484 29192
rect 20622 29180 20628 29192
rect 20680 29180 20686 29232
rect 21082 29180 21088 29232
rect 21140 29220 21146 29232
rect 25866 29220 25872 29232
rect 21140 29192 25872 29220
rect 21140 29180 21146 29192
rect 20441 29155 20499 29161
rect 20441 29121 20453 29155
rect 20487 29121 20499 29155
rect 20717 29155 20775 29161
rect 20717 29152 20729 29155
rect 20441 29115 20499 29121
rect 20640 29124 20729 29152
rect 15160 29056 15884 29084
rect 15160 29044 15166 29056
rect 11146 29016 11152 29028
rect 10980 28988 11152 29016
rect 11146 28976 11152 28988
rect 11204 29016 11210 29028
rect 11882 29016 11888 29028
rect 11204 28988 11888 29016
rect 11204 28976 11210 28988
rect 11882 28976 11888 28988
rect 11940 28976 11946 29028
rect 12434 28976 12440 29028
rect 12492 29016 12498 29028
rect 17126 29016 17132 29028
rect 12492 28988 17132 29016
rect 12492 28976 12498 28988
rect 17126 28976 17132 28988
rect 17184 28976 17190 29028
rect 20640 29016 20668 29124
rect 20717 29121 20729 29124
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 20809 29155 20867 29161
rect 20809 29121 20821 29155
rect 20855 29152 20867 29155
rect 20898 29152 20904 29164
rect 20855 29124 20904 29152
rect 20855 29121 20867 29124
rect 20809 29115 20867 29121
rect 20898 29112 20904 29124
rect 20956 29112 20962 29164
rect 23658 29112 23664 29164
rect 23716 29152 23722 29164
rect 24762 29152 24768 29164
rect 23716 29124 24768 29152
rect 23716 29112 23722 29124
rect 24762 29112 24768 29124
rect 24820 29112 24826 29164
rect 24964 29161 24992 29192
rect 25866 29180 25872 29192
rect 25924 29180 25930 29232
rect 33870 29220 33876 29232
rect 33831 29192 33876 29220
rect 33870 29180 33876 29192
rect 33928 29180 33934 29232
rect 24949 29155 25007 29161
rect 24949 29121 24961 29155
rect 24995 29121 25007 29155
rect 24949 29115 25007 29121
rect 25498 29112 25504 29164
rect 25556 29152 25562 29164
rect 25593 29155 25651 29161
rect 25593 29152 25605 29155
rect 25556 29124 25605 29152
rect 25556 29112 25562 29124
rect 25593 29121 25605 29124
rect 25639 29121 25651 29155
rect 29822 29152 29828 29164
rect 29783 29124 29828 29152
rect 25593 29115 25651 29121
rect 29822 29112 29828 29124
rect 29880 29112 29886 29164
rect 30009 29155 30067 29161
rect 30009 29121 30021 29155
rect 30055 29152 30067 29155
rect 30374 29152 30380 29164
rect 30055 29124 30380 29152
rect 30055 29121 30067 29124
rect 30009 29115 30067 29121
rect 23382 29044 23388 29096
rect 23440 29084 23446 29096
rect 30024 29084 30052 29115
rect 30374 29112 30380 29124
rect 30432 29152 30438 29164
rect 30469 29155 30527 29161
rect 30469 29152 30481 29155
rect 30432 29124 30481 29152
rect 30432 29112 30438 29124
rect 30469 29121 30481 29124
rect 30515 29121 30527 29155
rect 30469 29115 30527 29121
rect 32490 29112 32496 29164
rect 32548 29152 32554 29164
rect 33781 29155 33839 29161
rect 33781 29152 33793 29155
rect 32548 29124 33793 29152
rect 32548 29112 32554 29124
rect 33781 29121 33793 29124
rect 33827 29121 33839 29155
rect 33781 29115 33839 29121
rect 33965 29155 34023 29161
rect 33965 29121 33977 29155
rect 34011 29121 34023 29155
rect 33965 29115 34023 29121
rect 23440 29056 30052 29084
rect 23440 29044 23446 29056
rect 33042 29044 33048 29096
rect 33100 29084 33106 29096
rect 33980 29084 34008 29115
rect 34054 29112 34060 29164
rect 34112 29152 34118 29164
rect 34149 29155 34207 29161
rect 34149 29152 34161 29155
rect 34112 29124 34161 29152
rect 34112 29112 34118 29124
rect 34149 29121 34161 29124
rect 34195 29121 34207 29155
rect 34149 29115 34207 29121
rect 33100 29056 34008 29084
rect 34900 29084 34928 29251
rect 35986 29220 35992 29232
rect 35728 29192 35992 29220
rect 34974 29112 34980 29164
rect 35032 29152 35038 29164
rect 35434 29152 35440 29164
rect 35032 29124 35440 29152
rect 35032 29112 35038 29124
rect 35434 29112 35440 29124
rect 35492 29112 35498 29164
rect 35618 29152 35624 29164
rect 35579 29124 35624 29152
rect 35618 29112 35624 29124
rect 35676 29112 35682 29164
rect 35728 29161 35756 29192
rect 35986 29180 35992 29192
rect 36044 29180 36050 29232
rect 36081 29223 36139 29229
rect 36081 29189 36093 29223
rect 36127 29220 36139 29223
rect 38390 29223 38448 29229
rect 38390 29220 38402 29223
rect 36127 29192 38402 29220
rect 36127 29189 36139 29192
rect 36081 29183 36139 29189
rect 38390 29189 38402 29192
rect 38436 29189 38448 29223
rect 38390 29183 38448 29189
rect 35713 29155 35771 29161
rect 35713 29121 35725 29155
rect 35759 29121 35771 29155
rect 35713 29115 35771 29121
rect 35805 29155 35863 29161
rect 35805 29121 35817 29155
rect 35851 29121 35863 29155
rect 35805 29115 35863 29121
rect 35820 29084 35848 29115
rect 38562 29112 38568 29164
rect 38620 29152 38626 29164
rect 38657 29155 38715 29161
rect 38657 29152 38669 29155
rect 38620 29124 38669 29152
rect 38620 29112 38626 29124
rect 38657 29121 38669 29124
rect 38703 29121 38715 29155
rect 38657 29115 38715 29121
rect 34900 29056 35848 29084
rect 33100 29044 33106 29056
rect 33796 29028 33824 29056
rect 25590 29016 25596 29028
rect 20640 28988 25596 29016
rect 25590 28976 25596 28988
rect 25648 28976 25654 29028
rect 25774 29016 25780 29028
rect 25735 28988 25780 29016
rect 25774 28976 25780 28988
rect 25832 28976 25838 29028
rect 33778 28976 33784 29028
rect 33836 28976 33842 29028
rect 34238 28976 34244 29028
rect 34296 29016 34302 29028
rect 35434 29016 35440 29028
rect 34296 28988 35440 29016
rect 34296 28976 34302 28988
rect 35434 28976 35440 28988
rect 35492 28976 35498 29028
rect 35894 28976 35900 29028
rect 35952 29016 35958 29028
rect 37277 29019 37335 29025
rect 37277 29016 37289 29019
rect 35952 28988 37289 29016
rect 35952 28976 35958 28988
rect 37277 28985 37289 28988
rect 37323 28985 37335 29019
rect 37277 28979 37335 28985
rect 14366 28948 14372 28960
rect 14327 28920 14372 28948
rect 14366 28908 14372 28920
rect 14424 28908 14430 28960
rect 15470 28948 15476 28960
rect 15431 28920 15476 28948
rect 15470 28908 15476 28920
rect 15528 28908 15534 28960
rect 19610 28948 19616 28960
rect 19571 28920 19616 28948
rect 19610 28908 19616 28920
rect 19668 28908 19674 28960
rect 20530 28908 20536 28960
rect 20588 28948 20594 28960
rect 20993 28951 21051 28957
rect 20993 28948 21005 28951
rect 20588 28920 21005 28948
rect 20588 28908 20594 28920
rect 20993 28917 21005 28920
rect 21039 28917 21051 28951
rect 20993 28911 21051 28917
rect 30098 28908 30104 28960
rect 30156 28948 30162 28960
rect 33597 28951 33655 28957
rect 33597 28948 33609 28951
rect 30156 28920 33609 28948
rect 30156 28908 30162 28920
rect 33597 28917 33609 28920
rect 33643 28917 33655 28951
rect 33597 28911 33655 28917
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 10134 28744 10140 28756
rect 10095 28716 10140 28744
rect 10134 28704 10140 28716
rect 10192 28704 10198 28756
rect 12805 28747 12863 28753
rect 12805 28713 12817 28747
rect 12851 28744 12863 28747
rect 12894 28744 12900 28756
rect 12851 28716 12900 28744
rect 12851 28713 12863 28716
rect 12805 28707 12863 28713
rect 12894 28704 12900 28716
rect 12952 28704 12958 28756
rect 13814 28704 13820 28756
rect 13872 28744 13878 28756
rect 14461 28747 14519 28753
rect 14461 28744 14473 28747
rect 13872 28716 14473 28744
rect 13872 28704 13878 28716
rect 14461 28713 14473 28716
rect 14507 28744 14519 28747
rect 15010 28744 15016 28756
rect 14507 28716 15016 28744
rect 14507 28713 14519 28716
rect 14461 28707 14519 28713
rect 15010 28704 15016 28716
rect 15068 28704 15074 28756
rect 17862 28744 17868 28756
rect 17823 28716 17868 28744
rect 17862 28704 17868 28716
rect 17920 28704 17926 28756
rect 23382 28744 23388 28756
rect 17972 28716 23388 28744
rect 9217 28679 9275 28685
rect 9217 28645 9229 28679
rect 9263 28676 9275 28679
rect 10042 28676 10048 28688
rect 9263 28648 10048 28676
rect 9263 28645 9275 28648
rect 9217 28639 9275 28645
rect 10042 28636 10048 28648
rect 10100 28636 10106 28688
rect 16206 28636 16212 28688
rect 16264 28676 16270 28688
rect 17313 28679 17371 28685
rect 17313 28676 17325 28679
rect 16264 28648 17325 28676
rect 16264 28636 16270 28648
rect 17313 28645 17325 28648
rect 17359 28676 17371 28679
rect 17972 28676 18000 28716
rect 23382 28704 23388 28716
rect 23440 28704 23446 28756
rect 24670 28744 24676 28756
rect 24631 28716 24676 28744
rect 24670 28704 24676 28716
rect 24728 28704 24734 28756
rect 25498 28744 25504 28756
rect 25459 28716 25504 28744
rect 25498 28704 25504 28716
rect 25556 28704 25562 28756
rect 28997 28747 29055 28753
rect 28997 28713 29009 28747
rect 29043 28744 29055 28747
rect 29546 28744 29552 28756
rect 29043 28716 29552 28744
rect 29043 28713 29055 28716
rect 28997 28707 29055 28713
rect 29546 28704 29552 28716
rect 29604 28704 29610 28756
rect 30101 28747 30159 28753
rect 30101 28713 30113 28747
rect 30147 28744 30159 28747
rect 30558 28744 30564 28756
rect 30147 28716 30564 28744
rect 30147 28713 30159 28716
rect 30101 28707 30159 28713
rect 30558 28704 30564 28716
rect 30616 28744 30622 28756
rect 30616 28716 31754 28744
rect 30616 28704 30622 28716
rect 18414 28676 18420 28688
rect 17359 28648 18000 28676
rect 18156 28648 18420 28676
rect 17359 28645 17371 28648
rect 17313 28639 17371 28645
rect 4982 28608 4988 28620
rect 4895 28580 4988 28608
rect 2774 28500 2780 28552
rect 2832 28540 2838 28552
rect 2961 28543 3019 28549
rect 2832 28512 2877 28540
rect 2832 28500 2838 28512
rect 2961 28509 2973 28543
rect 3007 28540 3019 28543
rect 3694 28540 3700 28552
rect 3007 28512 3700 28540
rect 3007 28509 3019 28512
rect 2961 28503 3019 28509
rect 3694 28500 3700 28512
rect 3752 28540 3758 28552
rect 4908 28549 4936 28580
rect 4982 28568 4988 28580
rect 5040 28608 5046 28620
rect 9674 28608 9680 28620
rect 5040 28580 9680 28608
rect 5040 28568 5046 28580
rect 4709 28543 4767 28549
rect 4709 28540 4721 28543
rect 3752 28512 4721 28540
rect 3752 28500 3758 28512
rect 4709 28509 4721 28512
rect 4755 28509 4767 28543
rect 4709 28503 4767 28509
rect 4893 28543 4951 28549
rect 4893 28509 4905 28543
rect 4939 28509 4951 28543
rect 4893 28503 4951 28509
rect 5074 28500 5080 28552
rect 5132 28540 5138 28552
rect 9140 28549 9168 28580
rect 9674 28568 9680 28580
rect 9732 28568 9738 28620
rect 11701 28611 11759 28617
rect 11701 28577 11713 28611
rect 11747 28608 11759 28611
rect 12158 28608 12164 28620
rect 11747 28580 12164 28608
rect 11747 28577 11759 28580
rect 11701 28571 11759 28577
rect 9125 28543 9183 28549
rect 5132 28512 8432 28540
rect 5132 28500 5138 28512
rect 4985 28475 5043 28481
rect 4985 28441 4997 28475
rect 5031 28472 5043 28475
rect 5350 28472 5356 28484
rect 5031 28444 5356 28472
rect 5031 28441 5043 28444
rect 4985 28435 5043 28441
rect 5350 28432 5356 28444
rect 5408 28432 5414 28484
rect 5994 28432 6000 28484
rect 6052 28472 6058 28484
rect 7006 28472 7012 28484
rect 6052 28444 7012 28472
rect 6052 28432 6058 28444
rect 7006 28432 7012 28444
rect 7064 28472 7070 28484
rect 7101 28475 7159 28481
rect 7101 28472 7113 28475
rect 7064 28444 7113 28472
rect 7064 28432 7070 28444
rect 7101 28441 7113 28444
rect 7147 28441 7159 28475
rect 7101 28435 7159 28441
rect 7285 28475 7343 28481
rect 7285 28441 7297 28475
rect 7331 28472 7343 28475
rect 8202 28472 8208 28484
rect 7331 28444 8208 28472
rect 7331 28441 7343 28444
rect 7285 28435 7343 28441
rect 8202 28432 8208 28444
rect 8260 28432 8266 28484
rect 8404 28472 8432 28512
rect 9125 28509 9137 28543
rect 9171 28509 9183 28543
rect 9306 28540 9312 28552
rect 9267 28512 9312 28540
rect 9125 28503 9183 28509
rect 9306 28500 9312 28512
rect 9364 28500 9370 28552
rect 9398 28500 9404 28552
rect 9456 28540 9462 28552
rect 9769 28543 9827 28549
rect 9769 28540 9781 28543
rect 9456 28512 9781 28540
rect 9456 28500 9462 28512
rect 9769 28509 9781 28512
rect 9815 28509 9827 28543
rect 9950 28540 9956 28552
rect 9911 28512 9956 28540
rect 9769 28503 9827 28509
rect 9950 28500 9956 28512
rect 10008 28500 10014 28552
rect 11422 28540 11428 28552
rect 11383 28512 11428 28540
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 11716 28472 11744 28571
rect 12158 28568 12164 28580
rect 12216 28568 12222 28620
rect 14093 28611 14151 28617
rect 14093 28577 14105 28611
rect 14139 28608 14151 28611
rect 14366 28608 14372 28620
rect 14139 28580 14372 28608
rect 14139 28577 14151 28580
rect 14093 28571 14151 28577
rect 14366 28568 14372 28580
rect 14424 28608 14430 28620
rect 14918 28608 14924 28620
rect 14424 28580 14924 28608
rect 14424 28568 14430 28580
rect 14918 28568 14924 28580
rect 14976 28568 14982 28620
rect 18156 28608 18184 28648
rect 18414 28636 18420 28648
rect 18472 28636 18478 28688
rect 19889 28679 19947 28685
rect 19889 28645 19901 28679
rect 19935 28676 19947 28679
rect 20806 28676 20812 28688
rect 19935 28648 20812 28676
rect 19935 28645 19947 28648
rect 19889 28639 19947 28645
rect 20806 28636 20812 28648
rect 20864 28676 20870 28688
rect 21082 28676 21088 28688
rect 20864 28648 21088 28676
rect 20864 28636 20870 28648
rect 21082 28636 21088 28648
rect 21140 28636 21146 28688
rect 23934 28636 23940 28688
rect 23992 28676 23998 28688
rect 25222 28676 25228 28688
rect 23992 28648 25228 28676
rect 23992 28636 23998 28648
rect 25222 28636 25228 28648
rect 25280 28636 25286 28688
rect 25516 28676 25544 28704
rect 29270 28676 29276 28688
rect 25516 28648 29276 28676
rect 29270 28636 29276 28648
rect 29328 28636 29334 28688
rect 19610 28608 19616 28620
rect 18156 28580 18276 28608
rect 14277 28543 14335 28549
rect 14277 28509 14289 28543
rect 14323 28509 14335 28543
rect 14277 28503 14335 28509
rect 8404 28444 11744 28472
rect 13722 28432 13728 28484
rect 13780 28472 13786 28484
rect 14292 28472 14320 28503
rect 14826 28500 14832 28552
rect 14884 28540 14890 28552
rect 15470 28549 15476 28552
rect 15197 28543 15255 28549
rect 15197 28540 15209 28543
rect 14884 28512 15209 28540
rect 14884 28500 14890 28512
rect 15197 28509 15209 28512
rect 15243 28509 15255 28543
rect 15464 28540 15476 28549
rect 15431 28512 15476 28540
rect 15197 28503 15255 28509
rect 15464 28503 15476 28512
rect 15470 28500 15476 28503
rect 15528 28500 15534 28552
rect 17034 28500 17040 28552
rect 17092 28540 17098 28552
rect 17586 28540 17592 28552
rect 17092 28512 17592 28540
rect 17092 28500 17098 28512
rect 17586 28500 17592 28512
rect 17644 28540 17650 28552
rect 18138 28540 18144 28552
rect 17644 28512 18000 28540
rect 18099 28512 18144 28540
rect 17644 28500 17650 28512
rect 15010 28472 15016 28484
rect 13780 28444 15016 28472
rect 13780 28432 13786 28444
rect 15010 28432 15016 28444
rect 15068 28432 15074 28484
rect 17126 28472 17132 28484
rect 17087 28444 17132 28472
rect 17126 28432 17132 28444
rect 17184 28432 17190 28484
rect 17972 28472 18000 28512
rect 18138 28500 18144 28512
rect 18196 28500 18202 28552
rect 18248 28549 18276 28580
rect 18340 28580 19616 28608
rect 18340 28549 18368 28580
rect 19610 28568 19616 28580
rect 19668 28568 19674 28620
rect 22186 28568 22192 28620
rect 22244 28608 22250 28620
rect 22830 28608 22836 28620
rect 22244 28580 22836 28608
rect 22244 28568 22250 28580
rect 22830 28568 22836 28580
rect 22888 28608 22894 28620
rect 23293 28611 23351 28617
rect 23293 28608 23305 28611
rect 22888 28580 23305 28608
rect 22888 28568 22894 28580
rect 23293 28577 23305 28580
rect 23339 28577 23351 28611
rect 26510 28608 26516 28620
rect 23293 28571 23351 28577
rect 24780 28580 26516 28608
rect 18233 28543 18291 28549
rect 18233 28509 18245 28543
rect 18279 28509 18291 28543
rect 18233 28503 18291 28509
rect 18325 28543 18383 28549
rect 18325 28509 18337 28543
rect 18371 28509 18383 28543
rect 18325 28503 18383 28509
rect 18509 28543 18567 28549
rect 18509 28509 18521 28543
rect 18555 28509 18567 28543
rect 18509 28503 18567 28509
rect 19705 28543 19763 28549
rect 19705 28509 19717 28543
rect 19751 28540 19763 28543
rect 20441 28543 20499 28549
rect 20441 28540 20453 28543
rect 19751 28512 20453 28540
rect 19751 28509 19763 28512
rect 19705 28503 19763 28509
rect 20441 28509 20453 28512
rect 20487 28540 20499 28543
rect 21637 28543 21695 28549
rect 21637 28540 21649 28543
rect 20487 28512 21649 28540
rect 20487 28509 20499 28512
rect 20441 28503 20499 28509
rect 21637 28509 21649 28512
rect 21683 28540 21695 28543
rect 23106 28540 23112 28552
rect 21683 28512 22094 28540
rect 23067 28512 23112 28540
rect 21683 28509 21695 28512
rect 21637 28503 21695 28509
rect 18524 28472 18552 28503
rect 17972 28444 18552 28472
rect 22066 28472 22094 28512
rect 23106 28500 23112 28512
rect 23164 28500 23170 28552
rect 24780 28540 24808 28580
rect 26510 28568 26516 28580
rect 26568 28568 26574 28620
rect 29564 28608 29592 28704
rect 31726 28676 31754 28716
rect 32030 28704 32036 28756
rect 32088 28744 32094 28756
rect 32493 28747 32551 28753
rect 32493 28744 32505 28747
rect 32088 28716 32505 28744
rect 32088 28704 32094 28716
rect 32493 28713 32505 28716
rect 32539 28744 32551 28747
rect 32582 28744 32588 28756
rect 32539 28716 32588 28744
rect 32539 28713 32551 28716
rect 32493 28707 32551 28713
rect 32582 28704 32588 28716
rect 32640 28704 32646 28756
rect 34606 28744 34612 28756
rect 33520 28716 34612 28744
rect 33410 28676 33416 28688
rect 31726 28648 33416 28676
rect 33410 28636 33416 28648
rect 33468 28636 33474 28688
rect 29733 28611 29791 28617
rect 29733 28608 29745 28611
rect 29564 28580 29745 28608
rect 29733 28577 29745 28580
rect 29779 28577 29791 28611
rect 33520 28608 33548 28716
rect 34606 28704 34612 28716
rect 34664 28704 34670 28756
rect 35618 28704 35624 28756
rect 35676 28744 35682 28756
rect 35713 28747 35771 28753
rect 35713 28744 35725 28747
rect 35676 28716 35725 28744
rect 35676 28704 35682 28716
rect 35713 28713 35725 28716
rect 35759 28713 35771 28747
rect 35713 28707 35771 28713
rect 33686 28636 33692 28688
rect 33744 28676 33750 28688
rect 34514 28676 34520 28688
rect 33744 28648 34520 28676
rect 33744 28636 33750 28648
rect 34514 28636 34520 28648
rect 34572 28636 34578 28688
rect 29733 28571 29791 28577
rect 30024 28580 33548 28608
rect 33704 28580 35572 28608
rect 24596 28512 24808 28540
rect 24857 28543 24915 28549
rect 22465 28475 22523 28481
rect 22465 28472 22477 28475
rect 22066 28444 22477 28472
rect 22465 28441 22477 28444
rect 22511 28472 22523 28475
rect 24596 28472 24624 28512
rect 24857 28509 24869 28543
rect 24903 28540 24915 28543
rect 25590 28540 25596 28552
rect 24903 28512 25596 28540
rect 24903 28509 24915 28512
rect 24857 28503 24915 28509
rect 25590 28500 25596 28512
rect 25648 28500 25654 28552
rect 29822 28500 29828 28552
rect 29880 28540 29886 28552
rect 29917 28543 29975 28549
rect 29917 28540 29929 28543
rect 29880 28512 29929 28540
rect 29880 28500 29886 28512
rect 29917 28509 29929 28512
rect 29963 28509 29975 28543
rect 29917 28503 29975 28509
rect 22511 28444 24624 28472
rect 22511 28441 22523 28444
rect 22465 28435 22523 28441
rect 24670 28432 24676 28484
rect 24728 28472 24734 28484
rect 25041 28475 25099 28481
rect 25041 28472 25053 28475
rect 24728 28444 25053 28472
rect 24728 28432 24734 28444
rect 25041 28441 25053 28444
rect 25087 28441 25099 28475
rect 25041 28435 25099 28441
rect 3142 28404 3148 28416
rect 3103 28376 3148 28404
rect 3142 28364 3148 28376
rect 3200 28364 3206 28416
rect 5261 28407 5319 28413
rect 5261 28373 5273 28407
rect 5307 28404 5319 28407
rect 6730 28404 6736 28416
rect 5307 28376 6736 28404
rect 5307 28373 5319 28376
rect 5261 28367 5319 28373
rect 6730 28364 6736 28376
rect 6788 28364 6794 28416
rect 7374 28364 7380 28416
rect 7432 28404 7438 28416
rect 7469 28407 7527 28413
rect 7469 28404 7481 28407
rect 7432 28376 7481 28404
rect 7432 28364 7438 28376
rect 7469 28373 7481 28376
rect 7515 28373 7527 28407
rect 7469 28367 7527 28373
rect 9306 28364 9312 28416
rect 9364 28404 9370 28416
rect 9766 28404 9772 28416
rect 9364 28376 9772 28404
rect 9364 28364 9370 28376
rect 9766 28364 9772 28376
rect 9824 28364 9830 28416
rect 13446 28364 13452 28416
rect 13504 28404 13510 28416
rect 14182 28404 14188 28416
rect 13504 28376 14188 28404
rect 13504 28364 13510 28376
rect 14182 28364 14188 28376
rect 14240 28364 14246 28416
rect 15194 28364 15200 28416
rect 15252 28404 15258 28416
rect 15930 28404 15936 28416
rect 15252 28376 15936 28404
rect 15252 28364 15258 28376
rect 15930 28364 15936 28376
rect 15988 28404 15994 28416
rect 16577 28407 16635 28413
rect 16577 28404 16589 28407
rect 15988 28376 16589 28404
rect 15988 28364 15994 28376
rect 16577 28373 16589 28376
rect 16623 28373 16635 28407
rect 16577 28367 16635 28373
rect 22373 28407 22431 28413
rect 22373 28373 22385 28407
rect 22419 28404 22431 28407
rect 24210 28404 24216 28416
rect 22419 28376 24216 28404
rect 22419 28373 22431 28376
rect 22373 28367 22431 28373
rect 24210 28364 24216 28376
rect 24268 28404 24274 28416
rect 30024 28404 30052 28580
rect 32490 28500 32496 28552
rect 32548 28540 32554 28552
rect 33704 28549 33732 28580
rect 33597 28543 33655 28549
rect 33597 28540 33609 28543
rect 32548 28512 33609 28540
rect 32548 28500 32554 28512
rect 33597 28509 33609 28512
rect 33643 28509 33655 28543
rect 33597 28503 33655 28509
rect 33689 28543 33747 28549
rect 33689 28509 33701 28543
rect 33735 28509 33747 28543
rect 33689 28503 33747 28509
rect 33965 28543 34023 28549
rect 33965 28509 33977 28543
rect 34011 28540 34023 28543
rect 34698 28540 34704 28552
rect 34011 28512 34704 28540
rect 34011 28509 34023 28512
rect 33965 28503 34023 28509
rect 34698 28500 34704 28512
rect 34756 28500 34762 28552
rect 35342 28540 35348 28552
rect 35303 28512 35348 28540
rect 35342 28500 35348 28512
rect 35400 28500 35406 28552
rect 35544 28549 35572 28580
rect 35529 28543 35587 28549
rect 35529 28509 35541 28543
rect 35575 28540 35587 28543
rect 35894 28540 35900 28552
rect 35575 28512 35900 28540
rect 35575 28509 35587 28512
rect 35529 28503 35587 28509
rect 35894 28500 35900 28512
rect 35952 28500 35958 28552
rect 30742 28472 30748 28484
rect 30655 28444 30748 28472
rect 30742 28432 30748 28444
rect 30800 28472 30806 28484
rect 31205 28475 31263 28481
rect 31205 28472 31217 28475
rect 30800 28444 31217 28472
rect 30800 28432 30806 28444
rect 31205 28441 31217 28444
rect 31251 28441 31263 28475
rect 33778 28472 33784 28484
rect 33739 28444 33784 28472
rect 31205 28435 31263 28441
rect 33778 28432 33784 28444
rect 33836 28432 33842 28484
rect 24268 28376 30052 28404
rect 33413 28407 33471 28413
rect 24268 28364 24274 28376
rect 33413 28373 33425 28407
rect 33459 28404 33471 28407
rect 33686 28404 33692 28416
rect 33459 28376 33692 28404
rect 33459 28373 33471 28376
rect 33413 28367 33471 28373
rect 33686 28364 33692 28376
rect 33744 28364 33750 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 3694 28200 3700 28212
rect 3655 28172 3700 28200
rect 3694 28160 3700 28172
rect 3752 28160 3758 28212
rect 8202 28200 8208 28212
rect 8163 28172 8208 28200
rect 8202 28160 8208 28172
rect 8260 28160 8266 28212
rect 12526 28200 12532 28212
rect 9646 28172 12532 28200
rect 6546 28092 6552 28144
rect 6604 28132 6610 28144
rect 8220 28132 8248 28160
rect 6604 28104 7877 28132
rect 8220 28104 8800 28132
rect 6604 28092 6610 28104
rect 2590 28073 2596 28076
rect 2584 28027 2596 28073
rect 2648 28064 2654 28076
rect 6822 28064 6828 28076
rect 2648 28036 2684 28064
rect 6783 28036 6828 28064
rect 2590 28024 2596 28027
rect 2648 28024 2654 28036
rect 6822 28024 6828 28036
rect 6880 28024 6886 28076
rect 6914 28024 6920 28076
rect 6972 28064 6978 28076
rect 7081 28067 7139 28073
rect 7081 28064 7093 28067
rect 6972 28036 7093 28064
rect 6972 28024 6978 28036
rect 7081 28033 7093 28036
rect 7127 28033 7139 28067
rect 7081 28027 7139 28033
rect 2314 27996 2320 28008
rect 2275 27968 2320 27996
rect 2314 27956 2320 27968
rect 2372 27956 2378 28008
rect 7849 27996 7877 28104
rect 8662 28064 8668 28076
rect 8623 28036 8668 28064
rect 8662 28024 8668 28036
rect 8720 28024 8726 28076
rect 8772 28073 8800 28104
rect 8758 28067 8816 28073
rect 8758 28033 8770 28067
rect 8804 28033 8816 28067
rect 8938 28064 8944 28076
rect 8899 28036 8944 28064
rect 8758 28027 8816 28033
rect 8938 28024 8944 28036
rect 8996 28024 9002 28076
rect 9033 28067 9091 28073
rect 9033 28033 9045 28067
rect 9079 28033 9091 28067
rect 9033 28027 9091 28033
rect 9048 27996 9076 28027
rect 9122 28024 9128 28076
rect 9180 28073 9186 28076
rect 9180 28064 9188 28073
rect 9646 28064 9674 28172
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 12621 28203 12679 28209
rect 12621 28169 12633 28203
rect 12667 28169 12679 28203
rect 13814 28200 13820 28212
rect 12621 28163 12679 28169
rect 12728 28172 13820 28200
rect 12636 28132 12664 28163
rect 11624 28104 12664 28132
rect 9180 28036 9674 28064
rect 9180 28027 9188 28036
rect 9180 28024 9186 28027
rect 10686 28024 10692 28076
rect 10744 28064 10750 28076
rect 11517 28067 11575 28073
rect 11517 28064 11529 28067
rect 10744 28036 11529 28064
rect 10744 28024 10750 28036
rect 11517 28033 11529 28036
rect 11563 28033 11575 28067
rect 11624 28064 11652 28104
rect 11680 28067 11738 28073
rect 11680 28064 11692 28067
rect 11624 28036 11692 28064
rect 11517 28027 11575 28033
rect 11680 28033 11692 28036
rect 11726 28033 11738 28067
rect 11680 28027 11738 28033
rect 11780 28067 11838 28073
rect 11780 28033 11792 28067
rect 11826 28033 11838 28067
rect 11780 28027 11838 28033
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 12728 28064 12756 28172
rect 13814 28160 13820 28172
rect 13872 28160 13878 28212
rect 14182 28200 14188 28212
rect 14095 28172 14188 28200
rect 14182 28160 14188 28172
rect 14240 28200 14246 28212
rect 16206 28200 16212 28212
rect 14240 28172 16212 28200
rect 14240 28160 14246 28172
rect 16206 28160 16212 28172
rect 16264 28160 16270 28212
rect 16942 28200 16948 28212
rect 16855 28172 16948 28200
rect 16942 28160 16948 28172
rect 17000 28200 17006 28212
rect 17126 28200 17132 28212
rect 17000 28172 17132 28200
rect 17000 28160 17006 28172
rect 17126 28160 17132 28172
rect 17184 28160 17190 28212
rect 23842 28200 23848 28212
rect 22066 28172 23848 28200
rect 12805 28135 12863 28141
rect 12805 28101 12817 28135
rect 12851 28132 12863 28135
rect 13078 28132 13084 28144
rect 12851 28104 13084 28132
rect 12851 28101 12863 28104
rect 12805 28095 12863 28101
rect 13078 28092 13084 28104
rect 13136 28132 13142 28144
rect 15194 28132 15200 28144
rect 13136 28104 14964 28132
rect 15155 28104 15200 28132
rect 13136 28092 13142 28104
rect 12989 28067 13047 28073
rect 12989 28064 13001 28067
rect 11931 28036 12434 28064
rect 12728 28036 13001 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 11795 27996 11823 28027
rect 7849 27968 9076 27996
rect 11716 27968 11823 27996
rect 11716 27940 11744 27968
rect 11698 27888 11704 27940
rect 11756 27888 11762 27940
rect 12406 27928 12434 28036
rect 12989 28033 13001 28036
rect 13035 28033 13047 28067
rect 13446 28064 13452 28076
rect 13407 28036 13452 28064
rect 12989 28027 13047 28033
rect 13446 28024 13452 28036
rect 13504 28024 13510 28076
rect 13633 28067 13691 28073
rect 13633 28033 13645 28067
rect 13679 28033 13691 28067
rect 13633 28027 13691 28033
rect 12526 27956 12532 28008
rect 12584 27996 12590 28008
rect 13648 27996 13676 28027
rect 14734 28024 14740 28076
rect 14792 28064 14798 28076
rect 14936 28073 14964 28104
rect 15194 28092 15200 28104
rect 15252 28092 15258 28144
rect 16114 28092 16120 28144
rect 16172 28132 16178 28144
rect 17954 28132 17960 28144
rect 16172 28104 17960 28132
rect 16172 28092 16178 28104
rect 17954 28092 17960 28104
rect 18012 28132 18018 28144
rect 18601 28135 18659 28141
rect 18601 28132 18613 28135
rect 18012 28104 18613 28132
rect 18012 28092 18018 28104
rect 18601 28101 18613 28104
rect 18647 28101 18659 28135
rect 22066 28132 22094 28172
rect 23842 28160 23848 28172
rect 23900 28200 23906 28212
rect 24029 28203 24087 28209
rect 24029 28200 24041 28203
rect 23900 28172 24041 28200
rect 23900 28160 23906 28172
rect 24029 28169 24041 28172
rect 24075 28169 24087 28203
rect 24029 28163 24087 28169
rect 32600 28172 33640 28200
rect 18601 28095 18659 28101
rect 18708 28104 22094 28132
rect 14829 28067 14887 28073
rect 14829 28064 14841 28067
rect 14792 28036 14841 28064
rect 14792 28024 14798 28036
rect 14829 28033 14841 28036
rect 14875 28033 14887 28067
rect 14829 28027 14887 28033
rect 14922 28067 14980 28073
rect 14922 28033 14934 28067
rect 14968 28033 14980 28067
rect 14922 28027 14980 28033
rect 15010 28024 15016 28076
rect 15068 28064 15074 28076
rect 15105 28067 15163 28073
rect 15105 28064 15117 28067
rect 15068 28036 15117 28064
rect 15068 28024 15074 28036
rect 15105 28033 15117 28036
rect 15151 28033 15163 28067
rect 15105 28027 15163 28033
rect 14366 27996 14372 28008
rect 12584 27968 14372 27996
rect 12584 27956 12590 27968
rect 14366 27956 14372 27968
rect 14424 27956 14430 28008
rect 15120 27996 15148 28027
rect 15286 28024 15292 28076
rect 15344 28073 15350 28076
rect 15344 28064 15352 28073
rect 15344 28036 15389 28064
rect 15344 28027 15352 28036
rect 15344 28024 15350 28027
rect 16298 28024 16304 28076
rect 16356 28064 16362 28076
rect 18708 28064 18736 28104
rect 16356 28036 18736 28064
rect 18785 28067 18843 28073
rect 16356 28024 16362 28036
rect 18785 28033 18797 28067
rect 18831 28064 18843 28067
rect 19334 28064 19340 28076
rect 18831 28036 19340 28064
rect 18831 28033 18843 28036
rect 18785 28027 18843 28033
rect 19334 28024 19340 28036
rect 19392 28024 19398 28076
rect 20714 28064 20720 28076
rect 20675 28036 20720 28064
rect 20714 28024 20720 28036
rect 20772 28024 20778 28076
rect 23566 28064 23572 28076
rect 23308 28036 23572 28064
rect 16850 27996 16856 28008
rect 15120 27968 16856 27996
rect 16850 27956 16856 27968
rect 16908 27956 16914 28008
rect 20438 27996 20444 28008
rect 20399 27968 20444 27996
rect 20438 27956 20444 27968
rect 20496 27956 20502 28008
rect 12894 27928 12900 27940
rect 12406 27900 12900 27928
rect 12894 27888 12900 27900
rect 12952 27888 12958 27940
rect 13541 27931 13599 27937
rect 13541 27897 13553 27931
rect 13587 27928 13599 27931
rect 15102 27928 15108 27940
rect 13587 27900 15108 27928
rect 13587 27897 13599 27900
rect 13541 27891 13599 27897
rect 15102 27888 15108 27900
rect 15160 27888 15166 27940
rect 15473 27931 15531 27937
rect 15473 27897 15485 27931
rect 15519 27928 15531 27931
rect 18322 27928 18328 27940
rect 15519 27900 18328 27928
rect 15519 27897 15531 27900
rect 15473 27891 15531 27897
rect 18322 27888 18328 27900
rect 18380 27888 18386 27940
rect 4249 27863 4307 27869
rect 4249 27829 4261 27863
rect 4295 27860 4307 27863
rect 4614 27860 4620 27872
rect 4295 27832 4620 27860
rect 4295 27829 4307 27832
rect 4249 27823 4307 27829
rect 4614 27820 4620 27832
rect 4672 27820 4678 27872
rect 9214 27820 9220 27872
rect 9272 27860 9278 27872
rect 9309 27863 9367 27869
rect 9309 27860 9321 27863
rect 9272 27832 9321 27860
rect 9272 27820 9278 27832
rect 9309 27829 9321 27832
rect 9355 27829 9367 27863
rect 9766 27860 9772 27872
rect 9727 27832 9772 27860
rect 9309 27823 9367 27829
rect 9766 27820 9772 27832
rect 9824 27820 9830 27872
rect 11974 27820 11980 27872
rect 12032 27860 12038 27872
rect 12161 27863 12219 27869
rect 12161 27860 12173 27863
rect 12032 27832 12173 27860
rect 12032 27820 12038 27832
rect 12161 27829 12173 27832
rect 12207 27829 12219 27863
rect 12161 27823 12219 27829
rect 15378 27820 15384 27872
rect 15436 27860 15442 27872
rect 17681 27863 17739 27869
rect 17681 27860 17693 27863
rect 15436 27832 17693 27860
rect 15436 27820 15442 27832
rect 17681 27829 17693 27832
rect 17727 27860 17739 27863
rect 18414 27860 18420 27872
rect 17727 27832 18420 27860
rect 17727 27829 17739 27832
rect 17681 27823 17739 27829
rect 18414 27820 18420 27832
rect 18472 27820 18478 27872
rect 19521 27863 19579 27869
rect 19521 27829 19533 27863
rect 19567 27860 19579 27863
rect 19978 27860 19984 27872
rect 19567 27832 19984 27860
rect 19567 27829 19579 27832
rect 19521 27823 19579 27829
rect 19978 27820 19984 27832
rect 20036 27820 20042 27872
rect 22002 27860 22008 27872
rect 21963 27832 22008 27860
rect 22002 27820 22008 27832
rect 22060 27820 22066 27872
rect 23014 27820 23020 27872
rect 23072 27860 23078 27872
rect 23308 27869 23336 28036
rect 23566 28024 23572 28036
rect 23624 28064 23630 28076
rect 23937 28067 23995 28073
rect 23937 28064 23949 28067
rect 23624 28036 23949 28064
rect 23624 28024 23630 28036
rect 23937 28033 23949 28036
rect 23983 28033 23995 28067
rect 23937 28027 23995 28033
rect 29825 28067 29883 28073
rect 29825 28033 29837 28067
rect 29871 28064 29883 28067
rect 29914 28064 29920 28076
rect 29871 28036 29920 28064
rect 29871 28033 29883 28036
rect 29825 28027 29883 28033
rect 29914 28024 29920 28036
rect 29972 28024 29978 28076
rect 32490 28024 32496 28076
rect 32548 28064 32554 28076
rect 32600 28073 32628 28172
rect 32677 28135 32735 28141
rect 32677 28101 32689 28135
rect 32723 28132 32735 28135
rect 33410 28132 33416 28144
rect 32723 28104 33416 28132
rect 32723 28101 32735 28104
rect 32677 28095 32735 28101
rect 33410 28092 33416 28104
rect 33468 28092 33474 28144
rect 32585 28067 32643 28073
rect 32585 28064 32597 28067
rect 32548 28036 32597 28064
rect 32548 28024 32554 28036
rect 32585 28033 32597 28036
rect 32631 28033 32643 28067
rect 32585 28027 32643 28033
rect 32769 28067 32827 28073
rect 32769 28033 32781 28067
rect 32815 28033 32827 28067
rect 32950 28064 32956 28076
rect 32911 28036 32956 28064
rect 32769 28027 32827 28033
rect 30101 27999 30159 28005
rect 30101 27996 30113 27999
rect 28736 27968 30113 27996
rect 23293 27863 23351 27869
rect 23293 27860 23305 27863
rect 23072 27832 23305 27860
rect 23072 27820 23078 27832
rect 23293 27829 23305 27832
rect 23339 27829 23351 27863
rect 23293 27823 23351 27829
rect 24302 27820 24308 27872
rect 24360 27860 24366 27872
rect 28736 27869 28764 27968
rect 30101 27965 30113 27968
rect 30147 27996 30159 27999
rect 30558 27996 30564 28008
rect 30147 27968 30564 27996
rect 30147 27965 30159 27968
rect 30101 27959 30159 27965
rect 30558 27956 30564 27968
rect 30616 27956 30622 28008
rect 30837 27999 30895 28005
rect 30837 27965 30849 27999
rect 30883 27996 30895 27999
rect 32784 27996 32812 28027
rect 32950 28024 32956 28036
rect 33008 28024 33014 28076
rect 33612 28073 33640 28172
rect 33689 28135 33747 28141
rect 33689 28101 33701 28135
rect 33735 28132 33747 28135
rect 33735 28104 34744 28132
rect 33735 28101 33747 28104
rect 33689 28095 33747 28101
rect 33597 28067 33655 28073
rect 33597 28033 33609 28067
rect 33643 28033 33655 28067
rect 33597 28027 33655 28033
rect 33778 28024 33784 28076
rect 33836 28064 33842 28076
rect 33965 28067 34023 28073
rect 33836 28036 33929 28064
rect 33836 28024 33842 28036
rect 33965 28033 33977 28067
rect 34011 28064 34023 28067
rect 34054 28064 34060 28076
rect 34011 28036 34060 28064
rect 34011 28033 34023 28036
rect 33965 28027 34023 28033
rect 34054 28024 34060 28036
rect 34112 28024 34118 28076
rect 34514 28064 34520 28076
rect 34475 28036 34520 28064
rect 34514 28024 34520 28036
rect 34572 28024 34578 28076
rect 34716 28073 34744 28104
rect 34701 28067 34759 28073
rect 34701 28033 34713 28067
rect 34747 28064 34759 28067
rect 37274 28064 37280 28076
rect 34747 28036 37280 28064
rect 34747 28033 34759 28036
rect 34701 28027 34759 28033
rect 37274 28024 37280 28036
rect 37332 28024 37338 28076
rect 38654 28064 38660 28076
rect 38396 28036 38660 28064
rect 33796 27996 33824 28024
rect 30883 27968 33824 27996
rect 30883 27965 30895 27968
rect 30837 27959 30895 27965
rect 32582 27888 32588 27940
rect 32640 27928 32646 27940
rect 38396 27937 38424 28036
rect 38654 28024 38660 28036
rect 38712 28064 38718 28076
rect 38933 28067 38991 28073
rect 38933 28064 38945 28067
rect 38712 28036 38945 28064
rect 38712 28024 38718 28036
rect 38933 28033 38945 28036
rect 38979 28033 38991 28067
rect 38933 28027 38991 28033
rect 38381 27931 38439 27937
rect 38381 27928 38393 27931
rect 32640 27900 38393 27928
rect 32640 27888 32646 27900
rect 38381 27897 38393 27900
rect 38427 27897 38439 27931
rect 58158 27928 58164 27940
rect 58119 27900 58164 27928
rect 38381 27891 38439 27897
rect 58158 27888 58164 27900
rect 58216 27888 58222 27940
rect 28721 27863 28779 27869
rect 28721 27860 28733 27863
rect 24360 27832 28733 27860
rect 24360 27820 24366 27832
rect 28721 27829 28733 27832
rect 28767 27829 28779 27863
rect 32398 27860 32404 27872
rect 32359 27832 32404 27860
rect 28721 27823 28779 27829
rect 32398 27820 32404 27832
rect 32456 27820 32462 27872
rect 33413 27863 33471 27869
rect 33413 27829 33425 27863
rect 33459 27860 33471 27863
rect 33502 27860 33508 27872
rect 33459 27832 33508 27860
rect 33459 27829 33471 27832
rect 33413 27823 33471 27829
rect 33502 27820 33508 27832
rect 33560 27820 33566 27872
rect 34790 27820 34796 27872
rect 34848 27860 34854 27872
rect 34885 27863 34943 27869
rect 34885 27860 34897 27863
rect 34848 27832 34897 27860
rect 34848 27820 34854 27832
rect 34885 27829 34897 27832
rect 34931 27829 34943 27863
rect 40218 27860 40224 27872
rect 40179 27832 40224 27860
rect 34885 27823 34943 27829
rect 40218 27820 40224 27832
rect 40276 27820 40282 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 2590 27656 2596 27668
rect 2551 27628 2596 27656
rect 2590 27616 2596 27628
rect 2648 27616 2654 27668
rect 6914 27656 6920 27668
rect 6875 27628 6920 27656
rect 6914 27616 6920 27628
rect 6972 27616 6978 27668
rect 9861 27659 9919 27665
rect 9861 27625 9873 27659
rect 9907 27625 9919 27659
rect 9861 27619 9919 27625
rect 4890 27548 4896 27600
rect 4948 27588 4954 27600
rect 9876 27588 9904 27619
rect 10962 27616 10968 27668
rect 11020 27656 11026 27668
rect 13078 27656 13084 27668
rect 11020 27628 12940 27656
rect 13039 27628 13084 27656
rect 11020 27616 11026 27628
rect 11698 27588 11704 27600
rect 4948 27560 5120 27588
rect 9876 27560 11704 27588
rect 4948 27548 4954 27560
rect 4614 27520 4620 27532
rect 2884 27492 4620 27520
rect 2884 27461 2912 27492
rect 4614 27480 4620 27492
rect 4672 27480 4678 27532
rect 2869 27455 2927 27461
rect 2869 27421 2881 27455
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 2958 27449 3016 27455
rect 2958 27415 2970 27449
rect 3004 27415 3016 27449
rect 2958 27409 3016 27415
rect 3053 27452 3111 27458
rect 3053 27418 3065 27452
rect 3099 27418 3111 27452
rect 3053 27412 3111 27418
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27452 3295 27455
rect 3326 27452 3332 27464
rect 3283 27424 3332 27452
rect 3283 27421 3295 27424
rect 3237 27415 3295 27421
rect 3326 27412 3332 27424
rect 3384 27412 3390 27464
rect 3878 27412 3884 27464
rect 3936 27452 3942 27464
rect 4157 27455 4215 27461
rect 4157 27452 4169 27455
rect 3936 27424 4169 27452
rect 3936 27412 3942 27424
rect 4157 27421 4169 27424
rect 4203 27421 4215 27455
rect 4706 27452 4712 27464
rect 4667 27424 4712 27452
rect 4157 27415 4215 27421
rect 4706 27412 4712 27424
rect 4764 27412 4770 27464
rect 4802 27455 4860 27461
rect 4802 27421 4814 27455
rect 4848 27421 4860 27455
rect 4982 27452 4988 27464
rect 4943 27424 4988 27452
rect 4802 27415 4860 27421
rect 2976 27328 3004 27409
rect 3068 27384 3096 27412
rect 3142 27384 3148 27396
rect 3068 27356 3148 27384
rect 3142 27344 3148 27356
rect 3200 27344 3206 27396
rect 3970 27384 3976 27396
rect 3931 27356 3976 27384
rect 3970 27344 3976 27356
rect 4028 27344 4034 27396
rect 2958 27276 2964 27328
rect 3016 27276 3022 27328
rect 3602 27276 3608 27328
rect 3660 27316 3666 27328
rect 3789 27319 3847 27325
rect 3789 27316 3801 27319
rect 3660 27288 3801 27316
rect 3660 27276 3666 27288
rect 3789 27285 3801 27288
rect 3835 27285 3847 27319
rect 3988 27316 4016 27344
rect 4816 27316 4844 27415
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 5092 27461 5120 27560
rect 11698 27548 11704 27560
rect 11756 27548 11762 27600
rect 12912 27588 12940 27628
rect 13078 27616 13084 27628
rect 13136 27616 13142 27668
rect 16114 27656 16120 27668
rect 13188 27628 16120 27656
rect 13188 27588 13216 27628
rect 16114 27616 16120 27628
rect 16172 27616 16178 27668
rect 23106 27656 23112 27668
rect 22066 27628 23112 27656
rect 19334 27588 19340 27600
rect 12912 27560 13216 27588
rect 19247 27560 19340 27588
rect 19334 27548 19340 27560
rect 19392 27588 19398 27600
rect 22066 27588 22094 27628
rect 23106 27616 23112 27628
rect 23164 27616 23170 27668
rect 25222 27616 25228 27668
rect 25280 27656 25286 27668
rect 32398 27656 32404 27668
rect 25280 27628 32404 27656
rect 25280 27616 25286 27628
rect 32398 27616 32404 27628
rect 32456 27616 32462 27668
rect 37274 27656 37280 27668
rect 37235 27628 37280 27656
rect 37274 27616 37280 27628
rect 37332 27616 37338 27668
rect 19392 27560 22094 27588
rect 19392 27548 19398 27560
rect 28442 27548 28448 27600
rect 28500 27588 28506 27600
rect 28905 27591 28963 27597
rect 28905 27588 28917 27591
rect 28500 27560 28917 27588
rect 28500 27548 28506 27560
rect 28905 27557 28917 27560
rect 28951 27557 28963 27591
rect 28905 27551 28963 27557
rect 7466 27520 7472 27532
rect 7300 27492 7472 27520
rect 5077 27455 5135 27461
rect 5077 27421 5089 27455
rect 5123 27421 5135 27455
rect 5077 27415 5135 27421
rect 5215 27455 5273 27461
rect 5215 27421 5227 27455
rect 5261 27452 5273 27455
rect 5442 27452 5448 27464
rect 5261 27424 5448 27452
rect 5261 27421 5273 27424
rect 5215 27415 5273 27421
rect 5442 27412 5448 27424
rect 5500 27412 5506 27464
rect 5902 27412 5908 27464
rect 5960 27452 5966 27464
rect 6457 27455 6515 27461
rect 6457 27452 6469 27455
rect 5960 27424 6469 27452
rect 5960 27412 5966 27424
rect 6457 27421 6469 27424
rect 6503 27452 6515 27455
rect 7098 27452 7104 27464
rect 6503 27424 7104 27452
rect 6503 27421 6515 27424
rect 6457 27415 6515 27421
rect 7098 27412 7104 27424
rect 7156 27452 7162 27464
rect 7300 27461 7328 27492
rect 7466 27480 7472 27492
rect 7524 27480 7530 27532
rect 8938 27480 8944 27532
rect 8996 27520 9002 27532
rect 15013 27523 15071 27529
rect 8996 27492 9996 27520
rect 8996 27480 9002 27492
rect 9968 27464 9996 27492
rect 15013 27489 15025 27523
rect 15059 27520 15071 27523
rect 15286 27520 15292 27532
rect 15059 27492 15292 27520
rect 15059 27489 15071 27492
rect 15013 27483 15071 27489
rect 15286 27480 15292 27492
rect 15344 27480 15350 27532
rect 21266 27480 21272 27532
rect 21324 27520 21330 27532
rect 22002 27520 22008 27532
rect 21324 27492 21496 27520
rect 21324 27480 21330 27492
rect 7193 27455 7251 27461
rect 7193 27452 7205 27455
rect 7156 27424 7205 27452
rect 7156 27412 7162 27424
rect 7193 27421 7205 27424
rect 7239 27421 7251 27455
rect 7193 27415 7251 27421
rect 7285 27455 7343 27461
rect 7285 27421 7297 27455
rect 7331 27421 7343 27455
rect 7285 27415 7343 27421
rect 7374 27412 7380 27464
rect 7432 27452 7438 27464
rect 7432 27424 7477 27452
rect 7432 27412 7438 27424
rect 7558 27412 7564 27464
rect 7616 27452 7622 27464
rect 9766 27452 9772 27464
rect 7616 27424 8156 27452
rect 9679 27424 9772 27452
rect 7616 27412 7622 27424
rect 5000 27356 5488 27384
rect 3988 27288 4844 27316
rect 3789 27279 3847 27285
rect 4890 27276 4896 27328
rect 4948 27316 4954 27328
rect 5000 27316 5028 27356
rect 4948 27288 5028 27316
rect 4948 27276 4954 27288
rect 5074 27276 5080 27328
rect 5132 27316 5138 27328
rect 5353 27319 5411 27325
rect 5353 27316 5365 27319
rect 5132 27288 5365 27316
rect 5132 27276 5138 27288
rect 5353 27285 5365 27288
rect 5399 27285 5411 27319
rect 5460 27316 5488 27356
rect 7576 27316 7604 27412
rect 8128 27328 8156 27424
rect 9766 27412 9772 27424
rect 9824 27412 9830 27464
rect 9950 27452 9956 27464
rect 9911 27424 9956 27452
rect 9950 27412 9956 27424
rect 10008 27412 10014 27464
rect 11701 27455 11759 27461
rect 11701 27421 11713 27455
rect 11747 27452 11759 27455
rect 11747 27424 12204 27452
rect 11747 27421 11759 27424
rect 11701 27415 11759 27421
rect 9784 27384 9812 27412
rect 12176 27396 12204 27424
rect 13446 27412 13452 27464
rect 13504 27452 13510 27464
rect 14737 27455 14795 27461
rect 14737 27452 14749 27455
rect 13504 27424 14749 27452
rect 13504 27412 13510 27424
rect 14737 27421 14749 27424
rect 14783 27421 14795 27455
rect 14737 27415 14795 27421
rect 20806 27412 20812 27464
rect 20864 27452 20870 27464
rect 21468 27461 21496 27492
rect 21560 27492 22008 27520
rect 21560 27461 21588 27492
rect 22002 27480 22008 27492
rect 22060 27480 22066 27532
rect 26786 27520 26792 27532
rect 26747 27492 26792 27520
rect 26786 27480 26792 27492
rect 26844 27480 26850 27532
rect 21177 27455 21235 27461
rect 21177 27452 21189 27455
rect 20864 27424 21189 27452
rect 20864 27412 20870 27424
rect 21177 27421 21189 27424
rect 21223 27421 21235 27455
rect 21177 27415 21235 27421
rect 21361 27455 21419 27461
rect 21361 27421 21373 27455
rect 21407 27421 21419 27455
rect 21361 27415 21419 27421
rect 21453 27455 21511 27461
rect 21453 27421 21465 27455
rect 21499 27421 21511 27455
rect 21453 27415 21511 27421
rect 21545 27455 21603 27461
rect 21545 27421 21557 27455
rect 21591 27421 21603 27455
rect 21545 27415 21603 27421
rect 11974 27393 11980 27396
rect 11968 27384 11980 27393
rect 9784 27356 10456 27384
rect 11935 27356 11980 27384
rect 10428 27328 10456 27356
rect 11968 27347 11980 27356
rect 11974 27344 11980 27347
rect 12032 27344 12038 27396
rect 12158 27344 12164 27396
rect 12216 27384 12222 27396
rect 14826 27384 14832 27396
rect 12216 27356 14832 27384
rect 12216 27344 12222 27356
rect 14826 27344 14832 27356
rect 14884 27344 14890 27396
rect 16853 27387 16911 27393
rect 16853 27353 16865 27387
rect 16899 27353 16911 27387
rect 17034 27384 17040 27396
rect 16995 27356 17040 27384
rect 16853 27347 16911 27353
rect 8110 27316 8116 27328
rect 5460 27288 7604 27316
rect 8071 27288 8116 27316
rect 5353 27279 5411 27285
rect 8110 27276 8116 27288
rect 8168 27276 8174 27328
rect 10410 27316 10416 27328
rect 10371 27288 10416 27316
rect 10410 27276 10416 27288
rect 10468 27276 10474 27328
rect 15010 27276 15016 27328
rect 15068 27316 15074 27328
rect 16301 27319 16359 27325
rect 16301 27316 16313 27319
rect 15068 27288 16313 27316
rect 15068 27276 15074 27288
rect 16301 27285 16313 27288
rect 16347 27316 16359 27319
rect 16868 27316 16896 27347
rect 17034 27344 17040 27356
rect 17092 27344 17098 27396
rect 21376 27384 21404 27415
rect 21634 27412 21640 27464
rect 21692 27452 21698 27464
rect 22465 27455 22523 27461
rect 22465 27452 22477 27455
rect 21692 27424 22477 27452
rect 21692 27412 21698 27424
rect 22465 27421 22477 27424
rect 22511 27452 22523 27455
rect 24949 27455 25007 27461
rect 24949 27452 24961 27455
rect 22511 27424 24961 27452
rect 22511 27421 22523 27424
rect 22465 27415 22523 27421
rect 24949 27421 24961 27424
rect 24995 27421 25007 27455
rect 28920 27452 28948 27551
rect 31754 27548 31760 27600
rect 31812 27588 31818 27600
rect 31812 27560 35020 27588
rect 31812 27548 31818 27560
rect 30929 27523 30987 27529
rect 30929 27489 30941 27523
rect 30975 27520 30987 27523
rect 31570 27520 31576 27532
rect 30975 27492 31576 27520
rect 30975 27489 30987 27492
rect 30929 27483 30987 27489
rect 31570 27480 31576 27492
rect 31628 27480 31634 27532
rect 31665 27523 31723 27529
rect 31665 27489 31677 27523
rect 31711 27520 31723 27523
rect 32490 27520 32496 27532
rect 31711 27492 32496 27520
rect 31711 27489 31723 27492
rect 31665 27483 31723 27489
rect 32490 27480 32496 27492
rect 32548 27480 32554 27532
rect 32766 27480 32772 27532
rect 32824 27480 32830 27532
rect 31386 27452 31392 27464
rect 28920 27424 31248 27452
rect 31347 27424 31392 27452
rect 24949 27415 25007 27421
rect 21376 27356 22094 27384
rect 21542 27316 21548 27328
rect 16347 27288 21548 27316
rect 16347 27285 16359 27288
rect 16301 27279 16359 27285
rect 21542 27276 21548 27288
rect 21600 27276 21606 27328
rect 21818 27316 21824 27328
rect 21779 27288 21824 27316
rect 21818 27276 21824 27288
rect 21876 27276 21882 27328
rect 22066 27316 22094 27356
rect 22554 27344 22560 27396
rect 22612 27384 22618 27396
rect 22710 27387 22768 27393
rect 22710 27384 22722 27387
rect 22612 27356 22722 27384
rect 22612 27344 22618 27356
rect 22710 27353 22722 27356
rect 22756 27353 22768 27387
rect 22710 27347 22768 27353
rect 23198 27344 23204 27396
rect 23256 27384 23262 27396
rect 23750 27384 23756 27396
rect 23256 27356 23756 27384
rect 23256 27344 23262 27356
rect 23750 27344 23756 27356
rect 23808 27344 23814 27396
rect 24854 27344 24860 27396
rect 24912 27384 24918 27396
rect 25194 27387 25252 27393
rect 25194 27384 25206 27387
rect 24912 27356 25206 27384
rect 24912 27344 24918 27356
rect 25194 27353 25206 27356
rect 25240 27353 25252 27387
rect 25194 27347 25252 27353
rect 25958 27344 25964 27396
rect 26016 27384 26022 27396
rect 27034 27387 27092 27393
rect 27034 27384 27046 27387
rect 26016 27356 27046 27384
rect 26016 27344 26022 27356
rect 27034 27353 27046 27356
rect 27080 27353 27092 27387
rect 27034 27347 27092 27353
rect 28721 27387 28779 27393
rect 28721 27353 28733 27387
rect 28767 27384 28779 27387
rect 28994 27384 29000 27396
rect 28767 27356 29000 27384
rect 28767 27353 28779 27356
rect 28721 27347 28779 27353
rect 28994 27344 29000 27356
rect 29052 27344 29058 27396
rect 30374 27344 30380 27396
rect 30432 27384 30438 27396
rect 30662 27387 30720 27393
rect 30662 27384 30674 27387
rect 30432 27356 30674 27384
rect 30432 27344 30438 27356
rect 30662 27353 30674 27356
rect 30708 27353 30720 27387
rect 31220 27384 31248 27424
rect 31386 27412 31392 27424
rect 31444 27412 31450 27464
rect 32677 27455 32735 27461
rect 32677 27421 32689 27455
rect 32723 27421 32735 27455
rect 32677 27415 32735 27421
rect 32784 27446 32812 27480
rect 32968 27461 32996 27560
rect 33226 27480 33232 27532
rect 33284 27520 33290 27532
rect 33284 27492 34652 27520
rect 33284 27480 33290 27492
rect 33134 27461 33140 27464
rect 32861 27455 32919 27461
rect 32861 27446 32873 27455
rect 32784 27421 32873 27446
rect 32907 27421 32919 27455
rect 32968 27455 33030 27461
rect 32968 27424 32984 27455
rect 32784 27418 32919 27421
rect 32861 27415 32919 27418
rect 32972 27421 32984 27424
rect 33018 27421 33030 27455
rect 32972 27415 33030 27421
rect 33091 27455 33140 27461
rect 33091 27421 33103 27455
rect 33137 27421 33140 27455
rect 33091 27415 33140 27421
rect 32692 27384 32720 27415
rect 33134 27412 33140 27415
rect 33192 27412 33198 27464
rect 33410 27412 33416 27464
rect 33468 27452 33474 27464
rect 33962 27452 33968 27464
rect 33468 27424 33968 27452
rect 33468 27412 33474 27424
rect 33962 27412 33968 27424
rect 34020 27412 34026 27464
rect 34149 27455 34207 27461
rect 34149 27421 34161 27455
rect 34195 27452 34207 27455
rect 34514 27452 34520 27464
rect 34195 27424 34520 27452
rect 34195 27421 34207 27424
rect 34149 27415 34207 27421
rect 34514 27412 34520 27424
rect 34572 27412 34578 27464
rect 34624 27452 34652 27492
rect 34698 27452 34704 27464
rect 34611 27424 34704 27452
rect 34624 27421 34704 27424
rect 34698 27412 34704 27421
rect 34756 27412 34762 27464
rect 34790 27412 34796 27464
rect 34848 27452 34854 27464
rect 34992 27461 35020 27560
rect 34885 27455 34943 27461
rect 34885 27452 34897 27455
rect 34848 27424 34897 27452
rect 34848 27412 34854 27424
rect 34885 27421 34897 27424
rect 34931 27421 34943 27455
rect 34885 27415 34943 27421
rect 34977 27455 35035 27461
rect 34977 27421 34989 27455
rect 35023 27421 35035 27455
rect 34977 27415 35035 27421
rect 35066 27412 35072 27464
rect 35124 27452 35130 27464
rect 35434 27452 35440 27464
rect 35124 27424 35440 27452
rect 35124 27412 35130 27424
rect 35434 27412 35440 27424
rect 35492 27412 35498 27464
rect 38562 27412 38568 27464
rect 38620 27452 38626 27464
rect 38657 27455 38715 27461
rect 38657 27452 38669 27455
rect 38620 27424 38669 27452
rect 38620 27412 38626 27424
rect 38657 27421 38669 27424
rect 38703 27452 38715 27455
rect 40218 27452 40224 27464
rect 38703 27424 40224 27452
rect 38703 27421 38715 27424
rect 38657 27415 38715 27421
rect 40218 27412 40224 27424
rect 40276 27412 40282 27464
rect 33778 27384 33784 27396
rect 31220 27356 32720 27384
rect 33739 27356 33784 27384
rect 30662 27347 30720 27353
rect 23382 27316 23388 27328
rect 22066 27288 23388 27316
rect 23382 27276 23388 27288
rect 23440 27276 23446 27328
rect 23842 27316 23848 27328
rect 23803 27288 23848 27316
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 24118 27276 24124 27328
rect 24176 27316 24182 27328
rect 24397 27319 24455 27325
rect 24397 27316 24409 27319
rect 24176 27288 24409 27316
rect 24176 27276 24182 27288
rect 24397 27285 24409 27288
rect 24443 27285 24455 27319
rect 26326 27316 26332 27328
rect 26287 27288 26332 27316
rect 24397 27279 24455 27285
rect 26326 27276 26332 27288
rect 26384 27276 26390 27328
rect 28169 27319 28227 27325
rect 28169 27285 28181 27319
rect 28215 27316 28227 27319
rect 29362 27316 29368 27328
rect 28215 27288 29368 27316
rect 28215 27285 28227 27288
rect 28169 27279 28227 27285
rect 29362 27276 29368 27288
rect 29420 27276 29426 27328
rect 29546 27316 29552 27328
rect 29507 27288 29552 27316
rect 29546 27276 29552 27288
rect 29604 27276 29610 27328
rect 32692 27316 32720 27356
rect 33778 27344 33784 27356
rect 33836 27344 33842 27396
rect 35345 27387 35403 27393
rect 35345 27353 35357 27387
rect 35391 27384 35403 27387
rect 38390 27387 38448 27393
rect 38390 27384 38402 27387
rect 35391 27356 38402 27384
rect 35391 27353 35403 27356
rect 35345 27347 35403 27353
rect 38390 27353 38402 27356
rect 38436 27353 38448 27387
rect 38390 27347 38448 27353
rect 33226 27316 33232 27328
rect 32692 27288 33232 27316
rect 33226 27276 33232 27288
rect 33284 27276 33290 27328
rect 33321 27319 33379 27325
rect 33321 27285 33333 27319
rect 33367 27316 33379 27319
rect 33410 27316 33416 27328
rect 33367 27288 33416 27316
rect 33367 27285 33379 27288
rect 33321 27279 33379 27285
rect 33410 27276 33416 27288
rect 33468 27276 33474 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 3510 27072 3516 27124
rect 3568 27072 3574 27124
rect 4341 27115 4399 27121
rect 4341 27081 4353 27115
rect 4387 27112 4399 27115
rect 4890 27112 4896 27124
rect 4387 27084 4896 27112
rect 4387 27081 4399 27084
rect 4341 27075 4399 27081
rect 3528 26991 3556 27072
rect 2682 26936 2688 26988
rect 2740 26976 2746 26988
rect 3418 26976 3424 26988
rect 2740 26948 3424 26976
rect 2740 26936 2746 26948
rect 3418 26936 3424 26948
rect 3476 26936 3482 26988
rect 3510 26985 3568 26991
rect 3510 26951 3522 26985
rect 3556 26951 3568 26985
rect 3510 26945 3568 26951
rect 3602 26936 3608 26988
rect 3660 26979 3666 26988
rect 3789 26979 3847 26985
rect 3660 26951 3702 26979
rect 3660 26936 3666 26951
rect 3789 26945 3801 26979
rect 3835 26976 3847 26979
rect 4356 26976 4384 27075
rect 4890 27072 4896 27084
rect 4948 27072 4954 27124
rect 4982 27072 4988 27124
rect 5040 27112 5046 27124
rect 8938 27112 8944 27124
rect 5040 27084 8944 27112
rect 5040 27072 5046 27084
rect 4798 26976 4804 26988
rect 3835 26948 4384 26976
rect 4759 26948 4804 26976
rect 3835 26945 3847 26948
rect 3789 26939 3847 26945
rect 4798 26936 4804 26948
rect 4856 26936 4862 26988
rect 5092 26985 5120 27084
rect 7024 27053 7052 27084
rect 8938 27072 8944 27084
rect 8996 27072 9002 27124
rect 15473 27115 15531 27121
rect 15473 27081 15485 27115
rect 15519 27112 15531 27115
rect 16114 27112 16120 27124
rect 15519 27084 16120 27112
rect 15519 27081 15531 27084
rect 15473 27075 15531 27081
rect 16114 27072 16120 27084
rect 16172 27072 16178 27124
rect 17126 27072 17132 27124
rect 17184 27112 17190 27124
rect 17313 27115 17371 27121
rect 17313 27112 17325 27115
rect 17184 27084 17325 27112
rect 17184 27072 17190 27084
rect 17313 27081 17325 27084
rect 17359 27112 17371 27115
rect 24670 27112 24676 27124
rect 17359 27084 24676 27112
rect 17359 27081 17371 27084
rect 17313 27075 17371 27081
rect 24670 27072 24676 27084
rect 24728 27072 24734 27124
rect 24854 27112 24860 27124
rect 24815 27084 24860 27112
rect 24854 27072 24860 27084
rect 24912 27072 24918 27124
rect 25958 27112 25964 27124
rect 25919 27084 25964 27112
rect 25958 27072 25964 27084
rect 26016 27072 26022 27124
rect 30558 27072 30564 27124
rect 30616 27112 30622 27124
rect 30653 27115 30711 27121
rect 30653 27112 30665 27115
rect 30616 27084 30665 27112
rect 30616 27072 30622 27084
rect 30653 27081 30665 27084
rect 30699 27081 30711 27115
rect 30653 27075 30711 27081
rect 31478 27072 31484 27124
rect 31536 27112 31542 27124
rect 32493 27115 32551 27121
rect 32493 27112 32505 27115
rect 31536 27084 32505 27112
rect 31536 27072 31542 27084
rect 32493 27081 32505 27084
rect 32539 27112 32551 27115
rect 33134 27112 33140 27124
rect 32539 27084 33140 27112
rect 32539 27081 32551 27084
rect 32493 27075 32551 27081
rect 33134 27072 33140 27084
rect 33192 27072 33198 27124
rect 33962 27072 33968 27124
rect 34020 27112 34026 27124
rect 34517 27115 34575 27121
rect 34517 27112 34529 27115
rect 34020 27084 34529 27112
rect 34020 27072 34026 27084
rect 34517 27081 34529 27084
rect 34563 27081 34575 27115
rect 35066 27112 35072 27124
rect 35027 27084 35072 27112
rect 34517 27075 34575 27081
rect 35066 27072 35072 27084
rect 35124 27072 35130 27124
rect 5169 27047 5227 27053
rect 5169 27013 5181 27047
rect 5215 27013 5227 27047
rect 5169 27007 5227 27013
rect 7009 27047 7067 27053
rect 7009 27013 7021 27047
rect 7055 27013 7067 27047
rect 7009 27007 7067 27013
rect 7101 27047 7159 27053
rect 7101 27013 7113 27047
rect 7147 27044 7159 27047
rect 7742 27044 7748 27056
rect 7147 27016 7748 27044
rect 7147 27013 7159 27016
rect 7101 27007 7159 27013
rect 4894 26979 4952 26985
rect 4894 26945 4906 26979
rect 4940 26945 4952 26979
rect 4894 26939 4952 26945
rect 5077 26979 5135 26985
rect 5077 26945 5089 26979
rect 5123 26945 5135 26979
rect 5077 26939 5135 26945
rect 3694 26868 3700 26920
rect 3752 26908 3758 26920
rect 4909 26908 4937 26939
rect 3752 26880 4937 26908
rect 3752 26868 3758 26880
rect 5184 26840 5212 27007
rect 7742 27004 7748 27016
rect 7800 27004 7806 27056
rect 12342 27004 12348 27056
rect 12400 27044 12406 27056
rect 13081 27047 13139 27053
rect 13081 27044 13093 27047
rect 12400 27016 13093 27044
rect 12400 27004 12406 27016
rect 13081 27013 13093 27016
rect 13127 27013 13139 27047
rect 14826 27044 14832 27056
rect 14787 27016 14832 27044
rect 13081 27007 13139 27013
rect 14826 27004 14832 27016
rect 14884 27004 14890 27056
rect 21818 27004 21824 27056
rect 21876 27044 21882 27056
rect 22250 27047 22308 27053
rect 22250 27044 22262 27047
rect 21876 27016 22262 27044
rect 21876 27004 21882 27016
rect 22250 27013 22262 27016
rect 22296 27013 22308 27047
rect 22250 27007 22308 27013
rect 24118 27004 24124 27056
rect 24176 27044 24182 27056
rect 24176 27016 24624 27044
rect 24176 27004 24182 27016
rect 5266 26979 5324 26985
rect 5266 26945 5278 26979
rect 5312 26976 5396 26979
rect 6730 26976 6736 26988
rect 5312 26951 5488 26976
rect 5312 26945 5324 26951
rect 5368 26948 5488 26951
rect 6691 26948 6736 26976
rect 5266 26939 5324 26945
rect 5460 26920 5488 26948
rect 6730 26936 6736 26948
rect 6788 26936 6794 26988
rect 6822 26936 6828 26988
rect 6880 26976 6886 26988
rect 7239 26979 7297 26985
rect 7239 26976 7251 26979
rect 6880 26948 6925 26976
rect 7024 26948 7251 26976
rect 6880 26936 6886 26948
rect 5442 26868 5448 26920
rect 5500 26908 5506 26920
rect 7024 26908 7052 26948
rect 7239 26945 7251 26948
rect 7285 26976 7297 26979
rect 9122 26976 9128 26988
rect 7285 26948 9128 26976
rect 7285 26945 7297 26948
rect 7239 26939 7297 26945
rect 9122 26936 9128 26948
rect 9180 26936 9186 26988
rect 9950 26936 9956 26988
rect 10008 26976 10014 26988
rect 10689 26979 10747 26985
rect 10689 26976 10701 26979
rect 10008 26948 10701 26976
rect 10008 26936 10014 26948
rect 10689 26945 10701 26948
rect 10735 26945 10747 26979
rect 10689 26939 10747 26945
rect 12069 26979 12127 26985
rect 12069 26945 12081 26979
rect 12115 26976 12127 26979
rect 13722 26976 13728 26988
rect 12115 26948 13728 26976
rect 12115 26945 12127 26948
rect 12069 26939 12127 26945
rect 13722 26936 13728 26948
rect 13780 26936 13786 26988
rect 15930 26976 15936 26988
rect 15891 26948 15936 26976
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 16114 26976 16120 26988
rect 16075 26948 16120 26976
rect 16114 26936 16120 26948
rect 16172 26936 16178 26988
rect 17129 26979 17187 26985
rect 17129 26976 17141 26979
rect 16224 26948 17141 26976
rect 5500 26880 7052 26908
rect 5500 26868 5506 26880
rect 10870 26868 10876 26920
rect 10928 26908 10934 26920
rect 10965 26911 11023 26917
rect 10965 26908 10977 26911
rect 10928 26880 10977 26908
rect 10928 26868 10934 26880
rect 10965 26877 10977 26880
rect 11011 26908 11023 26911
rect 11793 26911 11851 26917
rect 11793 26908 11805 26911
rect 11011 26880 11805 26908
rect 11011 26877 11023 26880
rect 10965 26871 11023 26877
rect 11793 26877 11805 26880
rect 11839 26877 11851 26911
rect 15948 26908 15976 26936
rect 16224 26908 16252 26948
rect 17129 26945 17141 26948
rect 17175 26945 17187 26979
rect 18966 26976 18972 26988
rect 18927 26948 18972 26976
rect 17129 26939 17187 26945
rect 18966 26936 18972 26948
rect 19024 26936 19030 26988
rect 19150 26976 19156 26988
rect 19111 26948 19156 26976
rect 19150 26936 19156 26948
rect 19208 26936 19214 26988
rect 20073 26979 20131 26985
rect 20073 26945 20085 26979
rect 20119 26976 20131 26979
rect 20898 26976 20904 26988
rect 20119 26948 20904 26976
rect 20119 26945 20131 26948
rect 20073 26939 20131 26945
rect 20898 26936 20904 26948
rect 20956 26936 20962 26988
rect 24210 26976 24216 26988
rect 24171 26948 24216 26976
rect 24210 26936 24216 26948
rect 24268 26936 24274 26988
rect 24394 26976 24400 26988
rect 24355 26948 24400 26976
rect 24394 26936 24400 26948
rect 24452 26936 24458 26988
rect 24596 26985 24624 27016
rect 31570 27004 31576 27056
rect 31628 27044 31634 27056
rect 31628 27016 33180 27044
rect 31628 27004 31634 27016
rect 24492 26979 24550 26985
rect 24492 26945 24504 26979
rect 24538 26945 24550 26979
rect 24492 26939 24550 26945
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26945 24639 26979
rect 24581 26939 24639 26945
rect 15948 26880 16252 26908
rect 11793 26871 11851 26877
rect 16574 26868 16580 26920
rect 16632 26908 16638 26920
rect 16945 26911 17003 26917
rect 16945 26908 16957 26911
rect 16632 26880 16957 26908
rect 16632 26868 16638 26880
rect 16945 26877 16957 26880
rect 16991 26908 17003 26911
rect 17773 26911 17831 26917
rect 17773 26908 17785 26911
rect 16991 26880 17785 26908
rect 16991 26877 17003 26880
rect 16945 26871 17003 26877
rect 17773 26877 17785 26880
rect 17819 26877 17831 26911
rect 17773 26871 17831 26877
rect 18690 26868 18696 26920
rect 18748 26908 18754 26920
rect 19797 26911 19855 26917
rect 19797 26908 19809 26911
rect 18748 26880 19809 26908
rect 18748 26868 18754 26880
rect 19797 26877 19809 26880
rect 19843 26877 19855 26911
rect 19797 26871 19855 26877
rect 21634 26868 21640 26920
rect 21692 26908 21698 26920
rect 22005 26911 22063 26917
rect 22005 26908 22017 26911
rect 21692 26880 22017 26908
rect 21692 26868 21698 26880
rect 22005 26877 22017 26880
rect 22051 26877 22063 26911
rect 24504 26908 24532 26939
rect 24762 26936 24768 26988
rect 24820 26976 24826 26988
rect 25317 26979 25375 26985
rect 25317 26976 25329 26979
rect 24820 26948 25329 26976
rect 24820 26936 24826 26948
rect 25317 26945 25329 26948
rect 25363 26945 25375 26979
rect 25498 26976 25504 26988
rect 25459 26948 25504 26976
rect 25317 26939 25375 26945
rect 25498 26936 25504 26948
rect 25556 26936 25562 26988
rect 25593 26979 25651 26985
rect 25593 26945 25605 26979
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 25685 26979 25743 26985
rect 25685 26945 25697 26979
rect 25731 26976 25743 26979
rect 25774 26976 25780 26988
rect 25731 26948 25780 26976
rect 25731 26945 25743 26948
rect 25685 26939 25743 26945
rect 25038 26908 25044 26920
rect 24504 26880 25044 26908
rect 22005 26871 22063 26877
rect 25038 26868 25044 26880
rect 25096 26908 25102 26920
rect 25608 26908 25636 26939
rect 25774 26936 25780 26948
rect 25832 26976 25838 26988
rect 26973 26979 27031 26985
rect 26973 26976 26985 26979
rect 25832 26948 26985 26976
rect 25832 26936 25838 26948
rect 26973 26945 26985 26948
rect 27019 26945 27031 26979
rect 28994 26976 29000 26988
rect 26973 26939 27031 26945
rect 28276 26948 29000 26976
rect 25096 26880 25636 26908
rect 25096 26868 25102 26880
rect 5258 26840 5264 26852
rect 5184 26812 5264 26840
rect 5258 26800 5264 26812
rect 5316 26800 5322 26852
rect 21450 26840 21456 26852
rect 16408 26812 21456 26840
rect 16408 26784 16436 26812
rect 21450 26800 21456 26812
rect 21508 26800 21514 26852
rect 22940 26812 24440 26840
rect 22940 26784 22968 26812
rect 2682 26772 2688 26784
rect 2643 26744 2688 26772
rect 2682 26732 2688 26744
rect 2740 26732 2746 26784
rect 3142 26772 3148 26784
rect 3103 26744 3148 26772
rect 3142 26732 3148 26744
rect 3200 26732 3206 26784
rect 5442 26772 5448 26784
rect 5403 26744 5448 26772
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 7374 26772 7380 26784
rect 7335 26744 7380 26772
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 16025 26775 16083 26781
rect 16025 26741 16037 26775
rect 16071 26772 16083 26775
rect 16390 26772 16396 26784
rect 16071 26744 16396 26772
rect 16071 26741 16083 26744
rect 16025 26735 16083 26741
rect 16390 26732 16396 26744
rect 16448 26732 16454 26784
rect 19337 26775 19395 26781
rect 19337 26741 19349 26775
rect 19383 26772 19395 26775
rect 19702 26772 19708 26784
rect 19383 26744 19708 26772
rect 19383 26741 19395 26744
rect 19337 26735 19395 26741
rect 19702 26732 19708 26744
rect 19760 26732 19766 26784
rect 22922 26732 22928 26784
rect 22980 26732 22986 26784
rect 23385 26775 23443 26781
rect 23385 26741 23397 26775
rect 23431 26772 23443 26775
rect 23658 26772 23664 26784
rect 23431 26744 23664 26772
rect 23431 26741 23443 26744
rect 23385 26735 23443 26741
rect 23658 26732 23664 26744
rect 23716 26732 23722 26784
rect 24412 26772 24440 26812
rect 28276 26781 28304 26948
rect 28994 26936 29000 26948
rect 29052 26936 29058 26988
rect 29641 26979 29699 26985
rect 29641 26945 29653 26979
rect 29687 26976 29699 26979
rect 29822 26976 29828 26988
rect 29687 26948 29828 26976
rect 29687 26945 29699 26948
rect 29641 26939 29699 26945
rect 29822 26936 29828 26948
rect 29880 26936 29886 26988
rect 33152 26985 33180 27016
rect 33410 26985 33416 26988
rect 33137 26979 33195 26985
rect 33137 26945 33149 26979
rect 33183 26945 33195 26979
rect 33404 26976 33416 26985
rect 33371 26948 33416 26976
rect 33137 26939 33195 26945
rect 33404 26939 33416 26948
rect 33410 26936 33416 26939
rect 33468 26936 33474 26988
rect 29365 26911 29423 26917
rect 29365 26908 29377 26911
rect 28828 26880 29377 26908
rect 28261 26775 28319 26781
rect 28261 26772 28273 26775
rect 24412 26744 28273 26772
rect 28261 26741 28273 26744
rect 28307 26741 28319 26775
rect 28261 26735 28319 26741
rect 28718 26732 28724 26784
rect 28776 26772 28782 26784
rect 28828 26781 28856 26880
rect 29365 26877 29377 26880
rect 29411 26908 29423 26911
rect 31205 26911 31263 26917
rect 31205 26908 31217 26911
rect 29411 26880 31217 26908
rect 29411 26877 29423 26880
rect 29365 26871 29423 26877
rect 31205 26877 31217 26880
rect 31251 26908 31263 26911
rect 31386 26908 31392 26920
rect 31251 26880 31392 26908
rect 31251 26877 31263 26880
rect 31205 26871 31263 26877
rect 31386 26868 31392 26880
rect 31444 26868 31450 26920
rect 28813 26775 28871 26781
rect 28813 26772 28825 26775
rect 28776 26744 28825 26772
rect 28776 26732 28782 26744
rect 28813 26741 28825 26744
rect 28859 26741 28871 26775
rect 58158 26772 58164 26784
rect 58119 26744 58164 26772
rect 28813 26735 28871 26741
rect 58158 26732 58164 26744
rect 58216 26732 58222 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 3878 26528 3884 26580
rect 3936 26568 3942 26580
rect 6273 26571 6331 26577
rect 3936 26540 5488 26568
rect 3936 26528 3942 26540
rect 2869 26503 2927 26509
rect 2869 26469 2881 26503
rect 2915 26500 2927 26503
rect 2915 26472 4292 26500
rect 2915 26469 2927 26472
rect 2869 26463 2927 26469
rect 3694 26432 3700 26444
rect 3068 26404 3700 26432
rect 2590 26324 2596 26376
rect 2648 26364 2654 26376
rect 3068 26373 3096 26404
rect 3694 26392 3700 26404
rect 3752 26392 3758 26444
rect 3053 26367 3111 26373
rect 3053 26364 3065 26367
rect 2648 26336 3065 26364
rect 2648 26324 2654 26336
rect 3053 26333 3065 26336
rect 3099 26333 3111 26367
rect 3053 26327 3111 26333
rect 3237 26367 3295 26373
rect 3237 26333 3249 26367
rect 3283 26364 3295 26367
rect 3878 26364 3884 26376
rect 3283 26336 3884 26364
rect 3283 26333 3295 26336
rect 3237 26327 3295 26333
rect 3878 26324 3884 26336
rect 3936 26324 3942 26376
rect 4062 26364 4068 26376
rect 4023 26336 4068 26364
rect 4062 26324 4068 26336
rect 4120 26324 4126 26376
rect 4264 26373 4292 26472
rect 4154 26364 4212 26370
rect 4154 26330 4166 26364
rect 4200 26330 4212 26364
rect 4154 26324 4212 26330
rect 4254 26367 4312 26373
rect 4254 26333 4266 26367
rect 4300 26333 4312 26367
rect 4254 26327 4312 26333
rect 4433 26367 4491 26373
rect 4433 26333 4445 26367
rect 4479 26364 4491 26367
rect 4890 26364 4896 26376
rect 4479 26336 4896 26364
rect 4479 26333 4491 26336
rect 4433 26327 4491 26333
rect 4890 26324 4896 26336
rect 4948 26324 4954 26376
rect 5460 26364 5488 26540
rect 6273 26537 6285 26571
rect 6319 26568 6331 26571
rect 7558 26568 7564 26580
rect 6319 26540 7564 26568
rect 6319 26537 6331 26540
rect 6273 26531 6331 26537
rect 7558 26528 7564 26540
rect 7616 26528 7622 26580
rect 8110 26528 8116 26580
rect 8168 26568 8174 26580
rect 10873 26571 10931 26577
rect 10873 26568 10885 26571
rect 8168 26540 10885 26568
rect 8168 26528 8174 26540
rect 10873 26537 10885 26540
rect 10919 26537 10931 26571
rect 10873 26531 10931 26537
rect 11054 26528 11060 26580
rect 11112 26568 11118 26580
rect 12342 26568 12348 26580
rect 11112 26540 12348 26568
rect 11112 26528 11118 26540
rect 12342 26528 12348 26540
rect 12400 26568 12406 26580
rect 12897 26571 12955 26577
rect 12897 26568 12909 26571
rect 12400 26540 12909 26568
rect 12400 26528 12406 26540
rect 12897 26537 12909 26540
rect 12943 26537 12955 26571
rect 21818 26568 21824 26580
rect 12897 26531 12955 26537
rect 15856 26540 21824 26568
rect 7466 26500 7472 26512
rect 7116 26472 7472 26500
rect 6546 26392 6552 26444
rect 6604 26432 6610 26444
rect 6604 26404 7052 26432
rect 6604 26392 6610 26404
rect 5905 26367 5963 26373
rect 5905 26364 5917 26367
rect 5460 26336 5917 26364
rect 5905 26333 5917 26336
rect 5951 26364 5963 26367
rect 5994 26364 6000 26376
rect 5951 26336 6000 26364
rect 5951 26333 5963 26336
rect 5905 26327 5963 26333
rect 5994 26324 6000 26336
rect 6052 26324 6058 26376
rect 6089 26367 6147 26373
rect 6089 26333 6101 26367
rect 6135 26364 6147 26367
rect 6362 26364 6368 26376
rect 6135 26336 6368 26364
rect 6135 26333 6147 26336
rect 6089 26327 6147 26333
rect 6362 26324 6368 26336
rect 6420 26364 6426 26376
rect 6822 26364 6828 26376
rect 6420 26336 6828 26364
rect 6420 26324 6426 26336
rect 6822 26324 6828 26336
rect 6880 26324 6886 26376
rect 7024 26373 7052 26404
rect 7116 26373 7144 26472
rect 7466 26460 7472 26472
rect 7524 26460 7530 26512
rect 7929 26503 7987 26509
rect 7929 26469 7941 26503
rect 7975 26500 7987 26503
rect 11885 26503 11943 26509
rect 11885 26500 11897 26503
rect 7975 26472 11897 26500
rect 7975 26469 7987 26472
rect 7929 26463 7987 26469
rect 11885 26469 11897 26472
rect 11931 26500 11943 26503
rect 15856 26500 15884 26540
rect 21818 26528 21824 26540
rect 21876 26568 21882 26580
rect 23753 26571 23811 26577
rect 23753 26568 23765 26571
rect 21876 26540 23765 26568
rect 21876 26528 21882 26540
rect 23753 26537 23765 26540
rect 23799 26568 23811 26571
rect 24210 26568 24216 26580
rect 23799 26540 24216 26568
rect 23799 26537 23811 26540
rect 23753 26531 23811 26537
rect 24210 26528 24216 26540
rect 24268 26528 24274 26580
rect 25498 26528 25504 26580
rect 25556 26568 25562 26580
rect 25869 26571 25927 26577
rect 25869 26568 25881 26571
rect 25556 26540 25881 26568
rect 25556 26528 25562 26540
rect 25869 26537 25881 26540
rect 25915 26537 25927 26571
rect 25869 26531 25927 26537
rect 31570 26528 31576 26580
rect 31628 26568 31634 26580
rect 31665 26571 31723 26577
rect 31665 26568 31677 26571
rect 31628 26540 31677 26568
rect 31628 26528 31634 26540
rect 31665 26537 31677 26540
rect 31711 26537 31723 26571
rect 32582 26568 32588 26580
rect 32543 26540 32588 26568
rect 31665 26531 31723 26537
rect 32582 26528 32588 26540
rect 32640 26528 32646 26580
rect 11931 26472 15884 26500
rect 11931 26469 11943 26472
rect 11885 26463 11943 26469
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26333 7067 26367
rect 7009 26327 7067 26333
rect 7114 26367 7172 26373
rect 7377 26367 7435 26373
rect 7114 26333 7126 26367
rect 7160 26333 7172 26367
rect 7114 26327 7172 26333
rect 7214 26361 7272 26367
rect 7214 26327 7226 26361
rect 7260 26358 7272 26361
rect 7260 26327 7282 26358
rect 7377 26333 7389 26367
rect 7423 26364 7435 26367
rect 7944 26364 7972 26463
rect 15930 26460 15936 26512
rect 15988 26500 15994 26512
rect 20346 26500 20352 26512
rect 15988 26472 18276 26500
rect 20307 26472 20352 26500
rect 15988 26460 15994 26472
rect 14366 26432 14372 26444
rect 14327 26404 14372 26432
rect 14366 26392 14372 26404
rect 14424 26392 14430 26444
rect 16390 26432 16396 26444
rect 16351 26404 16396 26432
rect 16390 26392 16396 26404
rect 16448 26392 16454 26444
rect 18248 26441 18276 26472
rect 20346 26460 20352 26472
rect 20404 26460 20410 26512
rect 23198 26460 23204 26512
rect 23256 26500 23262 26512
rect 24765 26503 24823 26509
rect 24765 26500 24777 26503
rect 23256 26472 24777 26500
rect 23256 26460 23262 26472
rect 24765 26469 24777 26472
rect 24811 26469 24823 26503
rect 24765 26463 24823 26469
rect 18233 26435 18291 26441
rect 18233 26401 18245 26435
rect 18279 26401 18291 26435
rect 18233 26395 18291 26401
rect 19058 26392 19064 26444
rect 19116 26432 19122 26444
rect 21266 26432 21272 26444
rect 19116 26404 21272 26432
rect 19116 26392 19122 26404
rect 7423 26336 7972 26364
rect 7423 26333 7435 26336
rect 7377 26327 7435 26333
rect 3694 26256 3700 26308
rect 3752 26296 3758 26308
rect 3789 26299 3847 26305
rect 3789 26296 3801 26299
rect 3752 26268 3801 26296
rect 3752 26256 3758 26268
rect 3789 26265 3801 26268
rect 3835 26265 3847 26299
rect 3789 26259 3847 26265
rect 3510 26188 3516 26240
rect 3568 26228 3574 26240
rect 4172 26228 4200 26324
rect 7214 26321 7282 26327
rect 10594 26324 10600 26376
rect 10652 26364 10658 26376
rect 10781 26367 10839 26373
rect 10781 26364 10793 26367
rect 10652 26336 10793 26364
rect 10652 26324 10658 26336
rect 10781 26333 10793 26336
rect 10827 26364 10839 26367
rect 11698 26364 11704 26376
rect 10827 26336 11704 26364
rect 10827 26333 10839 26336
rect 10781 26327 10839 26333
rect 11698 26324 11704 26336
rect 11756 26324 11762 26376
rect 13446 26324 13452 26376
rect 13504 26364 13510 26376
rect 14093 26367 14151 26373
rect 14093 26364 14105 26367
rect 13504 26336 14105 26364
rect 13504 26324 13510 26336
rect 14093 26333 14105 26336
rect 14139 26333 14151 26367
rect 16114 26364 16120 26376
rect 16075 26336 16120 26364
rect 14093 26327 14151 26333
rect 16114 26324 16120 26336
rect 16172 26324 16178 26376
rect 17129 26367 17187 26373
rect 17129 26364 17141 26367
rect 16224 26336 17141 26364
rect 4614 26256 4620 26308
rect 4672 26296 4678 26308
rect 4982 26296 4988 26308
rect 4672 26268 4988 26296
rect 4672 26256 4678 26268
rect 4982 26256 4988 26268
rect 5040 26296 5046 26308
rect 5353 26299 5411 26305
rect 5353 26296 5365 26299
rect 5040 26268 5365 26296
rect 5040 26256 5046 26268
rect 5353 26265 5365 26268
rect 5399 26296 5411 26299
rect 6546 26296 6552 26308
rect 5399 26268 6552 26296
rect 5399 26265 5411 26268
rect 5353 26259 5411 26265
rect 6546 26256 6552 26268
rect 6604 26256 6610 26308
rect 6730 26296 6736 26308
rect 6691 26268 6736 26296
rect 6730 26256 6736 26268
rect 6788 26256 6794 26308
rect 7254 26296 7282 26321
rect 7558 26296 7564 26308
rect 7254 26268 7564 26296
rect 7558 26256 7564 26268
rect 7616 26256 7622 26308
rect 10410 26256 10416 26308
rect 10468 26296 10474 26308
rect 15102 26296 15108 26308
rect 10468 26268 15108 26296
rect 10468 26256 10474 26268
rect 15102 26256 15108 26268
rect 15160 26296 15166 26308
rect 16224 26296 16252 26336
rect 17129 26333 17141 26336
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 18509 26367 18567 26373
rect 18509 26333 18521 26367
rect 18555 26364 18567 26367
rect 18690 26364 18696 26376
rect 18555 26336 18696 26364
rect 18555 26333 18567 26336
rect 18509 26327 18567 26333
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 19628 26373 19656 26404
rect 21266 26392 21272 26404
rect 21324 26392 21330 26444
rect 22002 26392 22008 26444
rect 22060 26432 22066 26444
rect 25774 26432 25780 26444
rect 22060 26404 25780 26432
rect 22060 26392 22066 26404
rect 25774 26392 25780 26404
rect 25832 26392 25838 26444
rect 37829 26435 37887 26441
rect 37829 26401 37841 26435
rect 37875 26432 37887 26435
rect 38562 26432 38568 26444
rect 37875 26404 38568 26432
rect 37875 26401 37887 26404
rect 37829 26395 37887 26401
rect 38562 26392 38568 26404
rect 38620 26392 38626 26444
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 16942 26296 16948 26308
rect 15160 26268 16252 26296
rect 16903 26268 16948 26296
rect 15160 26256 15166 26268
rect 16942 26256 16948 26268
rect 17000 26256 17006 26308
rect 19536 26296 19564 26327
rect 19702 26324 19708 26376
rect 19760 26364 19766 26376
rect 19889 26367 19947 26373
rect 19760 26336 19805 26364
rect 19760 26324 19766 26336
rect 19889 26333 19901 26367
rect 19935 26364 19947 26367
rect 20806 26364 20812 26376
rect 19935 26336 20812 26364
rect 19935 26333 19947 26336
rect 19889 26327 19947 26333
rect 20806 26324 20812 26336
rect 20864 26324 20870 26376
rect 23201 26367 23259 26373
rect 23201 26333 23213 26367
rect 23247 26364 23259 26367
rect 25225 26367 25283 26373
rect 25225 26364 25237 26367
rect 23247 26336 25237 26364
rect 23247 26333 23259 26336
rect 23201 26327 23259 26333
rect 25225 26333 25237 26336
rect 25271 26364 25283 26367
rect 30377 26367 30435 26373
rect 30377 26364 30389 26367
rect 25271 26336 30389 26364
rect 25271 26333 25283 26336
rect 25225 26327 25283 26333
rect 30377 26333 30389 26336
rect 30423 26364 30435 26367
rect 32582 26364 32588 26376
rect 30423 26336 32588 26364
rect 30423 26333 30435 26336
rect 30377 26327 30435 26333
rect 32582 26324 32588 26336
rect 32640 26324 32646 26376
rect 38473 26367 38531 26373
rect 38473 26333 38485 26367
rect 38519 26364 38531 26367
rect 38930 26364 38936 26376
rect 38519 26336 38936 26364
rect 38519 26333 38531 26336
rect 38473 26327 38531 26333
rect 38930 26324 38936 26336
rect 38988 26324 38994 26376
rect 20346 26296 20352 26308
rect 19536 26268 20352 26296
rect 20346 26256 20352 26268
rect 20404 26256 20410 26308
rect 21634 26296 21640 26308
rect 21595 26268 21640 26296
rect 21634 26256 21640 26268
rect 21692 26256 21698 26308
rect 23658 26256 23664 26308
rect 23716 26296 23722 26308
rect 24210 26296 24216 26308
rect 23716 26268 24216 26296
rect 23716 26256 23722 26268
rect 24210 26256 24216 26268
rect 24268 26256 24274 26308
rect 24394 26296 24400 26308
rect 24355 26268 24400 26296
rect 24394 26256 24400 26268
rect 24452 26256 24458 26308
rect 24581 26299 24639 26305
rect 24581 26265 24593 26299
rect 24627 26265 24639 26299
rect 24581 26259 24639 26265
rect 26053 26299 26111 26305
rect 26053 26265 26065 26299
rect 26099 26265 26111 26299
rect 26053 26259 26111 26265
rect 7466 26228 7472 26240
rect 3568 26200 7472 26228
rect 3568 26188 3574 26200
rect 7466 26188 7472 26200
rect 7524 26188 7530 26240
rect 18414 26188 18420 26240
rect 18472 26228 18478 26240
rect 18598 26228 18604 26240
rect 18472 26200 18604 26228
rect 18472 26188 18478 26200
rect 18598 26188 18604 26200
rect 18656 26188 18662 26240
rect 19242 26228 19248 26240
rect 19203 26200 19248 26228
rect 19242 26188 19248 26200
rect 19300 26188 19306 26240
rect 23474 26188 23480 26240
rect 23532 26228 23538 26240
rect 23842 26228 23848 26240
rect 23532 26200 23848 26228
rect 23532 26188 23538 26200
rect 23842 26188 23848 26200
rect 23900 26228 23906 26240
rect 24596 26228 24624 26259
rect 23900 26200 24624 26228
rect 26068 26228 26096 26259
rect 26142 26256 26148 26308
rect 26200 26296 26206 26308
rect 26237 26299 26295 26305
rect 26237 26296 26249 26299
rect 26200 26268 26249 26296
rect 26200 26256 26206 26268
rect 26237 26265 26249 26268
rect 26283 26265 26295 26299
rect 29362 26296 29368 26308
rect 26237 26259 26295 26265
rect 26344 26268 29368 26296
rect 26344 26228 26372 26268
rect 29362 26256 29368 26268
rect 29420 26256 29426 26308
rect 37274 26256 37280 26308
rect 37332 26296 37338 26308
rect 37562 26299 37620 26305
rect 37562 26296 37574 26299
rect 37332 26268 37574 26296
rect 37332 26256 37338 26268
rect 37562 26265 37574 26268
rect 37608 26265 37620 26299
rect 37562 26259 37620 26265
rect 38657 26299 38715 26305
rect 38657 26265 38669 26299
rect 38703 26296 38715 26299
rect 39022 26296 39028 26308
rect 38703 26268 39028 26296
rect 38703 26265 38715 26268
rect 38657 26259 38715 26265
rect 39022 26256 39028 26268
rect 39080 26256 39086 26308
rect 29638 26228 29644 26240
rect 26068 26200 26372 26228
rect 29599 26200 29644 26228
rect 23900 26188 23906 26200
rect 29638 26188 29644 26200
rect 29696 26188 29702 26240
rect 36449 26231 36507 26237
rect 36449 26197 36461 26231
rect 36495 26228 36507 26231
rect 36630 26228 36636 26240
rect 36495 26200 36636 26228
rect 36495 26197 36507 26200
rect 36449 26191 36507 26197
rect 36630 26188 36636 26200
rect 36688 26188 36694 26240
rect 38010 26188 38016 26240
rect 38068 26228 38074 26240
rect 38289 26231 38347 26237
rect 38289 26228 38301 26231
rect 38068 26200 38301 26228
rect 38068 26188 38074 26200
rect 38289 26197 38301 26200
rect 38335 26197 38347 26231
rect 38289 26191 38347 26197
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 3970 26024 3976 26036
rect 3931 25996 3976 26024
rect 3970 25984 3976 25996
rect 4028 25984 4034 26036
rect 4062 25984 4068 26036
rect 4120 26024 4126 26036
rect 5261 26027 5319 26033
rect 5261 26024 5273 26027
rect 4120 25996 5273 26024
rect 4120 25984 4126 25996
rect 5261 25993 5273 25996
rect 5307 25993 5319 26027
rect 6362 26024 6368 26036
rect 6323 25996 6368 26024
rect 5261 25987 5319 25993
rect 6362 25984 6368 25996
rect 6420 25984 6426 26036
rect 14185 26027 14243 26033
rect 14185 25993 14197 26027
rect 14231 26024 14243 26027
rect 14366 26024 14372 26036
rect 14231 25996 14372 26024
rect 14231 25993 14243 25996
rect 14185 25987 14243 25993
rect 14366 25984 14372 25996
rect 14424 26024 14430 26036
rect 18141 26027 18199 26033
rect 14424 25996 15056 26024
rect 14424 25984 14430 25996
rect 15028 25968 15056 25996
rect 18141 25993 18153 26027
rect 18187 26024 18199 26027
rect 19150 26024 19156 26036
rect 18187 25996 19156 26024
rect 18187 25993 18199 25996
rect 18141 25987 18199 25993
rect 19150 25984 19156 25996
rect 19208 26024 19214 26036
rect 20714 26024 20720 26036
rect 19208 25996 20720 26024
rect 19208 25984 19214 25996
rect 20714 25984 20720 25996
rect 20772 25984 20778 26036
rect 21082 25984 21088 26036
rect 21140 26024 21146 26036
rect 21177 26027 21235 26033
rect 21177 26024 21189 26027
rect 21140 25996 21189 26024
rect 21140 25984 21146 25996
rect 21177 25993 21189 25996
rect 21223 25993 21235 26027
rect 21177 25987 21235 25993
rect 21266 25984 21272 26036
rect 21324 26024 21330 26036
rect 22465 26027 22523 26033
rect 21324 25996 22140 26024
rect 21324 25984 21330 25996
rect 2860 25959 2918 25965
rect 2860 25925 2872 25959
rect 2906 25956 2918 25959
rect 3142 25956 3148 25968
rect 2906 25928 3148 25956
rect 2906 25925 2918 25928
rect 2860 25919 2918 25925
rect 3142 25916 3148 25928
rect 3200 25916 3206 25968
rect 4801 25959 4859 25965
rect 4801 25925 4813 25959
rect 4847 25956 4859 25959
rect 4890 25956 4896 25968
rect 4847 25928 4896 25956
rect 4847 25925 4859 25928
rect 4801 25919 4859 25925
rect 4890 25916 4896 25928
rect 4948 25916 4954 25968
rect 6730 25916 6736 25968
rect 6788 25956 6794 25968
rect 7478 25959 7536 25965
rect 7478 25956 7490 25959
rect 6788 25928 7490 25956
rect 6788 25916 6794 25928
rect 7478 25925 7490 25928
rect 7524 25925 7536 25959
rect 7478 25919 7536 25925
rect 13449 25959 13507 25965
rect 13449 25925 13461 25959
rect 13495 25956 13507 25959
rect 13906 25956 13912 25968
rect 13495 25928 13912 25956
rect 13495 25925 13507 25928
rect 13449 25919 13507 25925
rect 13906 25916 13912 25928
rect 13964 25916 13970 25968
rect 14642 25956 14648 25968
rect 14603 25928 14648 25956
rect 14642 25916 14648 25928
rect 14700 25916 14706 25968
rect 15010 25916 15016 25968
rect 15068 25956 15074 25968
rect 15473 25959 15531 25965
rect 15473 25956 15485 25959
rect 15068 25928 15485 25956
rect 15068 25916 15074 25928
rect 15473 25925 15485 25928
rect 15519 25925 15531 25959
rect 15473 25919 15531 25925
rect 19242 25916 19248 25968
rect 19300 25965 19306 25968
rect 19300 25956 19312 25965
rect 19300 25928 19345 25956
rect 19300 25919 19312 25928
rect 19300 25916 19306 25919
rect 20806 25916 20812 25968
rect 20864 25956 20870 25968
rect 20864 25928 21864 25956
rect 20864 25916 20870 25928
rect 2314 25848 2320 25900
rect 2372 25888 2378 25900
rect 2593 25891 2651 25897
rect 2593 25888 2605 25891
rect 2372 25860 2605 25888
rect 2372 25848 2378 25860
rect 2593 25857 2605 25860
rect 2639 25857 2651 25891
rect 2593 25851 2651 25857
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25857 9551 25891
rect 9674 25888 9680 25900
rect 9635 25860 9680 25888
rect 9493 25851 9551 25857
rect 7745 25823 7803 25829
rect 7745 25789 7757 25823
rect 7791 25789 7803 25823
rect 9508 25820 9536 25851
rect 9674 25848 9680 25860
rect 9732 25848 9738 25900
rect 11698 25848 11704 25900
rect 11756 25888 11762 25900
rect 12529 25891 12587 25897
rect 12529 25888 12541 25891
rect 11756 25860 12541 25888
rect 11756 25848 11762 25860
rect 12529 25857 12541 25860
rect 12575 25857 12587 25891
rect 13633 25891 13691 25897
rect 13633 25888 13645 25891
rect 12529 25851 12587 25857
rect 12728 25860 13645 25888
rect 9766 25820 9772 25832
rect 9508 25792 9772 25820
rect 7745 25783 7803 25789
rect 6822 25644 6828 25696
rect 6880 25684 6886 25696
rect 7760 25684 7788 25783
rect 9766 25780 9772 25792
rect 9824 25820 9830 25832
rect 12728 25820 12756 25860
rect 13633 25857 13645 25860
rect 13679 25857 13691 25891
rect 13633 25851 13691 25857
rect 9824 25792 12756 25820
rect 12805 25823 12863 25829
rect 9824 25780 9830 25792
rect 12805 25789 12817 25823
rect 12851 25820 12863 25823
rect 12986 25820 12992 25832
rect 12851 25792 12992 25820
rect 12851 25789 12863 25792
rect 12805 25783 12863 25789
rect 10965 25755 11023 25761
rect 10965 25721 10977 25755
rect 11011 25752 11023 25755
rect 12820 25752 12848 25783
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 13648 25820 13676 25851
rect 14274 25848 14280 25900
rect 14332 25888 14338 25900
rect 14829 25891 14887 25897
rect 14829 25888 14841 25891
rect 14332 25860 14841 25888
rect 14332 25848 14338 25860
rect 14829 25857 14841 25860
rect 14875 25857 14887 25891
rect 17126 25888 17132 25900
rect 17087 25860 17132 25888
rect 14829 25851 14887 25857
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 17218 25848 17224 25900
rect 17276 25888 17282 25900
rect 21836 25897 21864 25928
rect 22112 25897 22140 25996
rect 22465 25993 22477 26027
rect 22511 26024 22523 26027
rect 22554 26024 22560 26036
rect 22511 25996 22560 26024
rect 22511 25993 22523 25996
rect 22465 25987 22523 25993
rect 22554 25984 22560 25996
rect 22612 25984 22618 26036
rect 23382 25984 23388 26036
rect 23440 26024 23446 26036
rect 24305 26027 24363 26033
rect 24305 26024 24317 26027
rect 23440 25996 24317 26024
rect 23440 25984 23446 25996
rect 24305 25993 24317 25996
rect 24351 25993 24363 26027
rect 24305 25987 24363 25993
rect 30285 26027 30343 26033
rect 30285 25993 30297 26027
rect 30331 26024 30343 26027
rect 30374 26024 30380 26036
rect 30331 25996 30380 26024
rect 30331 25993 30343 25996
rect 30285 25987 30343 25993
rect 30374 25984 30380 25996
rect 30432 25984 30438 26036
rect 37274 26024 37280 26036
rect 37235 25996 37280 26024
rect 37274 25984 37280 25996
rect 37332 25984 37338 26036
rect 23566 25956 23572 25968
rect 23527 25928 23572 25956
rect 23566 25916 23572 25928
rect 23624 25916 23630 25968
rect 24210 25956 24216 25968
rect 23768 25928 24216 25956
rect 21821 25891 21879 25897
rect 17276 25860 21772 25888
rect 17276 25848 17282 25860
rect 19521 25823 19579 25829
rect 13648 25792 15700 25820
rect 11011 25724 12848 25752
rect 11011 25721 11023 25724
rect 10965 25715 11023 25721
rect 15672 25696 15700 25792
rect 19521 25789 19533 25823
rect 19567 25820 19579 25823
rect 21634 25820 21640 25832
rect 19567 25792 21640 25820
rect 19567 25789 19579 25792
rect 19521 25783 19579 25789
rect 6880 25656 7788 25684
rect 9861 25687 9919 25693
rect 6880 25644 6886 25656
rect 9861 25653 9873 25687
rect 9907 25684 9919 25687
rect 10778 25684 10784 25696
rect 9907 25656 10784 25684
rect 9907 25653 9919 25656
rect 9861 25647 9919 25653
rect 10778 25644 10784 25656
rect 10836 25644 10842 25696
rect 13078 25644 13084 25696
rect 13136 25684 13142 25696
rect 13265 25687 13323 25693
rect 13265 25684 13277 25687
rect 13136 25656 13277 25684
rect 13136 25644 13142 25656
rect 13265 25653 13277 25656
rect 13311 25653 13323 25687
rect 15562 25684 15568 25696
rect 15523 25656 15568 25684
rect 13265 25647 13323 25653
rect 15562 25644 15568 25656
rect 15620 25644 15626 25696
rect 15654 25644 15660 25696
rect 15712 25684 15718 25696
rect 16945 25687 17003 25693
rect 16945 25684 16957 25687
rect 15712 25656 16957 25684
rect 15712 25644 15718 25656
rect 16945 25653 16957 25656
rect 16991 25653 17003 25687
rect 16945 25647 17003 25653
rect 19242 25644 19248 25696
rect 19300 25684 19306 25696
rect 19536 25684 19564 25783
rect 21634 25780 21640 25792
rect 21692 25780 21698 25832
rect 21744 25752 21772 25860
rect 21821 25857 21833 25891
rect 21867 25857 21879 25891
rect 21821 25851 21879 25857
rect 22005 25891 22063 25897
rect 22005 25857 22017 25891
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22097 25891 22155 25897
rect 22097 25857 22109 25891
rect 22143 25857 22155 25891
rect 22097 25851 22155 25857
rect 22020 25820 22048 25851
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22244 25860 22289 25888
rect 22244 25848 22250 25860
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 23768 25897 23796 25928
rect 24210 25916 24216 25928
rect 24268 25956 24274 25968
rect 24489 25959 24547 25965
rect 24489 25956 24501 25959
rect 24268 25928 24501 25956
rect 24268 25916 24274 25928
rect 24489 25925 24501 25928
rect 24535 25925 24547 25959
rect 24489 25919 24547 25925
rect 25777 25959 25835 25965
rect 25777 25925 25789 25959
rect 25823 25956 25835 25959
rect 26326 25956 26332 25968
rect 25823 25928 26332 25956
rect 25823 25925 25835 25928
rect 25777 25919 25835 25925
rect 26326 25916 26332 25928
rect 26384 25956 26390 25968
rect 27430 25956 27436 25968
rect 26384 25928 27436 25956
rect 26384 25916 26390 25928
rect 27430 25916 27436 25928
rect 27488 25916 27494 25968
rect 31570 25956 31576 25968
rect 28828 25928 31576 25956
rect 23339 25891 23397 25897
rect 23339 25888 23351 25891
rect 23164 25860 23351 25888
rect 23164 25848 23170 25860
rect 23339 25857 23351 25860
rect 23385 25857 23397 25891
rect 23339 25851 23397 25857
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 23752 25891 23810 25897
rect 23752 25857 23764 25891
rect 23798 25857 23810 25891
rect 23752 25851 23810 25857
rect 23198 25820 23204 25832
rect 22020 25792 23204 25820
rect 23198 25780 23204 25792
rect 23256 25780 23262 25832
rect 23382 25752 23388 25764
rect 21744 25724 23388 25752
rect 23382 25712 23388 25724
rect 23440 25712 23446 25764
rect 23492 25752 23520 25851
rect 23842 25848 23848 25900
rect 23900 25888 23906 25900
rect 23900 25860 23945 25888
rect 23900 25848 23906 25860
rect 24394 25848 24400 25900
rect 24452 25888 24458 25900
rect 24673 25891 24731 25897
rect 24673 25888 24685 25891
rect 24452 25860 24685 25888
rect 24452 25848 24458 25860
rect 24673 25857 24685 25860
rect 24719 25857 24731 25891
rect 24673 25851 24731 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25888 26019 25891
rect 26050 25888 26056 25900
rect 26007 25860 26056 25888
rect 26007 25857 26019 25860
rect 25961 25851 26019 25857
rect 26050 25848 26056 25860
rect 26108 25848 26114 25900
rect 27614 25848 27620 25900
rect 27672 25888 27678 25900
rect 28546 25891 28604 25897
rect 28546 25888 28558 25891
rect 27672 25860 28558 25888
rect 27672 25848 27678 25860
rect 28546 25857 28558 25860
rect 28592 25857 28604 25891
rect 28546 25851 28604 25857
rect 28828 25832 28856 25928
rect 31570 25916 31576 25928
rect 31628 25916 31634 25968
rect 38746 25916 38752 25968
rect 38804 25956 38810 25968
rect 40742 25959 40800 25965
rect 40742 25956 40754 25959
rect 38804 25928 40754 25956
rect 38804 25916 38810 25928
rect 40742 25925 40754 25928
rect 40788 25925 40800 25959
rect 40742 25919 40800 25925
rect 29638 25888 29644 25900
rect 29599 25860 29644 25888
rect 29638 25848 29644 25860
rect 29696 25848 29702 25900
rect 29822 25888 29828 25900
rect 29783 25860 29828 25888
rect 29822 25848 29828 25860
rect 29880 25848 29886 25900
rect 29920 25891 29978 25897
rect 29920 25857 29932 25891
rect 29966 25857 29978 25891
rect 29920 25851 29978 25857
rect 30009 25891 30067 25897
rect 30009 25857 30021 25891
rect 30055 25888 30067 25891
rect 30190 25888 30196 25900
rect 30055 25860 30196 25888
rect 30055 25857 30067 25860
rect 30009 25851 30067 25857
rect 24486 25780 24492 25832
rect 24544 25820 24550 25832
rect 25593 25823 25651 25829
rect 25593 25820 25605 25823
rect 24544 25792 25605 25820
rect 24544 25780 24550 25792
rect 25593 25789 25605 25792
rect 25639 25789 25651 25823
rect 25593 25783 25651 25789
rect 28810 25780 28816 25832
rect 28868 25820 28874 25832
rect 28868 25792 28961 25820
rect 28868 25780 28874 25792
rect 29932 25764 29960 25851
rect 30190 25848 30196 25860
rect 30248 25848 30254 25900
rect 36633 25891 36691 25897
rect 36633 25888 36645 25891
rect 31726 25860 36645 25888
rect 27798 25752 27804 25764
rect 23492 25724 27804 25752
rect 27798 25712 27804 25724
rect 27856 25712 27862 25764
rect 29914 25712 29920 25764
rect 29972 25712 29978 25764
rect 30374 25712 30380 25764
rect 30432 25752 30438 25764
rect 31297 25755 31355 25761
rect 31297 25752 31309 25755
rect 30432 25724 31309 25752
rect 30432 25712 30438 25724
rect 31297 25721 31309 25724
rect 31343 25752 31355 25755
rect 31726 25752 31754 25860
rect 36633 25857 36645 25860
rect 36679 25888 36691 25891
rect 37182 25888 37188 25900
rect 36679 25860 37188 25888
rect 36679 25857 36691 25860
rect 36633 25851 36691 25857
rect 37182 25848 37188 25860
rect 37240 25888 37246 25900
rect 37533 25891 37591 25897
rect 37533 25888 37545 25891
rect 37240 25860 37545 25888
rect 37240 25848 37246 25860
rect 37533 25857 37545 25860
rect 37579 25857 37591 25891
rect 37533 25851 37591 25857
rect 37642 25891 37700 25897
rect 37642 25857 37654 25891
rect 37688 25857 37700 25891
rect 37642 25851 37700 25857
rect 37737 25891 37795 25897
rect 37737 25857 37749 25891
rect 37783 25888 37795 25891
rect 37826 25888 37832 25900
rect 37783 25860 37832 25888
rect 37783 25857 37795 25860
rect 37737 25851 37795 25857
rect 31343 25724 31754 25752
rect 31343 25721 31355 25724
rect 31297 25715 31355 25721
rect 37550 25712 37556 25764
rect 37608 25752 37614 25764
rect 37660 25752 37688 25851
rect 37826 25848 37832 25860
rect 37884 25848 37890 25900
rect 37918 25848 37924 25900
rect 37976 25888 37982 25900
rect 37976 25860 38021 25888
rect 37976 25848 37982 25860
rect 38562 25848 38568 25900
rect 38620 25888 38626 25900
rect 39770 25891 39828 25897
rect 39770 25888 39782 25891
rect 38620 25860 39782 25888
rect 38620 25848 38626 25860
rect 39770 25857 39782 25860
rect 39816 25857 39828 25891
rect 39770 25851 39828 25857
rect 40037 25891 40095 25897
rect 40037 25857 40049 25891
rect 40083 25888 40095 25891
rect 40218 25888 40224 25900
rect 40083 25860 40224 25888
rect 40083 25857 40095 25860
rect 40037 25851 40095 25857
rect 40218 25848 40224 25860
rect 40276 25888 40282 25900
rect 40497 25891 40555 25897
rect 40497 25888 40509 25891
rect 40276 25860 40509 25888
rect 40276 25848 40282 25860
rect 40497 25857 40509 25860
rect 40543 25857 40555 25891
rect 40497 25851 40555 25857
rect 37608 25724 37688 25752
rect 37608 25712 37614 25724
rect 19300 25656 19564 25684
rect 19300 25644 19306 25656
rect 22186 25644 22192 25696
rect 22244 25684 22250 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 22244 25656 23213 25684
rect 22244 25644 22250 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 23290 25644 23296 25696
rect 23348 25684 23354 25696
rect 27433 25687 27491 25693
rect 27433 25684 27445 25687
rect 23348 25656 27445 25684
rect 23348 25644 23354 25656
rect 27433 25653 27445 25656
rect 27479 25684 27491 25687
rect 27890 25684 27896 25696
rect 27479 25656 27896 25684
rect 27479 25653 27491 25656
rect 27433 25647 27491 25653
rect 27890 25644 27896 25656
rect 27948 25644 27954 25696
rect 30190 25644 30196 25696
rect 30248 25684 30254 25696
rect 30745 25687 30803 25693
rect 30745 25684 30757 25687
rect 30248 25656 30757 25684
rect 30248 25644 30254 25656
rect 30745 25653 30757 25656
rect 30791 25684 30803 25687
rect 37458 25684 37464 25696
rect 30791 25656 37464 25684
rect 30791 25653 30803 25656
rect 30745 25647 30803 25653
rect 37458 25644 37464 25656
rect 37516 25644 37522 25696
rect 38657 25687 38715 25693
rect 38657 25653 38669 25687
rect 38703 25684 38715 25687
rect 38930 25684 38936 25696
rect 38703 25656 38936 25684
rect 38703 25653 38715 25656
rect 38657 25647 38715 25653
rect 38930 25644 38936 25656
rect 38988 25644 38994 25696
rect 39850 25644 39856 25696
rect 39908 25684 39914 25696
rect 41877 25687 41935 25693
rect 41877 25684 41889 25687
rect 39908 25656 41889 25684
rect 39908 25644 39914 25656
rect 41877 25653 41889 25656
rect 41923 25653 41935 25687
rect 41877 25647 41935 25653
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 9030 25480 9036 25492
rect 8991 25452 9036 25480
rect 9030 25440 9036 25452
rect 9088 25440 9094 25492
rect 17218 25480 17224 25492
rect 10704 25452 17224 25480
rect 3786 25372 3792 25424
rect 3844 25412 3850 25424
rect 10134 25412 10140 25424
rect 3844 25384 10140 25412
rect 3844 25372 3850 25384
rect 10134 25372 10140 25384
rect 10192 25412 10198 25424
rect 10704 25421 10732 25452
rect 17218 25440 17224 25452
rect 17276 25440 17282 25492
rect 18414 25440 18420 25492
rect 18472 25480 18478 25492
rect 18509 25483 18567 25489
rect 18509 25480 18521 25483
rect 18472 25452 18521 25480
rect 18472 25440 18478 25452
rect 18509 25449 18521 25452
rect 18555 25449 18567 25483
rect 22370 25480 22376 25492
rect 18509 25443 18567 25449
rect 18616 25452 22376 25480
rect 10689 25415 10747 25421
rect 10689 25412 10701 25415
rect 10192 25384 10701 25412
rect 10192 25372 10198 25384
rect 10689 25381 10701 25384
rect 10735 25381 10747 25415
rect 10689 25375 10747 25381
rect 16761 25415 16819 25421
rect 16761 25381 16773 25415
rect 16807 25412 16819 25415
rect 16942 25412 16948 25424
rect 16807 25384 16948 25412
rect 16807 25381 16819 25384
rect 16761 25375 16819 25381
rect 16942 25372 16948 25384
rect 17000 25372 17006 25424
rect 11054 25344 11060 25356
rect 7668 25316 11060 25344
rect 7668 25285 7696 25316
rect 11054 25304 11060 25316
rect 11112 25304 11118 25356
rect 12158 25344 12164 25356
rect 12119 25316 12164 25344
rect 12158 25304 12164 25316
rect 12216 25304 12222 25356
rect 18616 25353 18644 25452
rect 22370 25440 22376 25452
rect 22428 25440 22434 25492
rect 23382 25440 23388 25492
rect 23440 25480 23446 25492
rect 26970 25480 26976 25492
rect 23440 25452 26976 25480
rect 23440 25440 23446 25452
rect 26970 25440 26976 25452
rect 27028 25440 27034 25492
rect 28997 25483 29055 25489
rect 28997 25449 29009 25483
rect 29043 25480 29055 25483
rect 29822 25480 29828 25492
rect 29043 25452 29828 25480
rect 29043 25449 29055 25452
rect 28997 25443 29055 25449
rect 29822 25440 29828 25452
rect 29880 25440 29886 25492
rect 36817 25483 36875 25489
rect 36817 25449 36829 25483
rect 36863 25480 36875 25483
rect 37826 25480 37832 25492
rect 36863 25452 37832 25480
rect 36863 25449 36875 25452
rect 36817 25443 36875 25449
rect 37826 25440 37832 25452
rect 37884 25440 37890 25492
rect 38562 25480 38568 25492
rect 38523 25452 38568 25480
rect 38562 25440 38568 25452
rect 38620 25440 38626 25492
rect 37752 25384 38352 25412
rect 18601 25347 18659 25353
rect 18601 25313 18613 25347
rect 18647 25313 18659 25347
rect 19242 25344 19248 25356
rect 19203 25316 19248 25344
rect 18601 25307 18659 25313
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 22646 25304 22652 25356
rect 22704 25344 22710 25356
rect 27249 25347 27307 25353
rect 22704 25316 23612 25344
rect 22704 25304 22710 25316
rect 7193 25279 7251 25285
rect 7193 25245 7205 25279
rect 7239 25276 7251 25279
rect 7653 25279 7711 25285
rect 7653 25276 7665 25279
rect 7239 25248 7665 25276
rect 7239 25245 7251 25248
rect 7193 25239 7251 25245
rect 7653 25245 7665 25248
rect 7699 25245 7711 25279
rect 7653 25239 7711 25245
rect 9030 25236 9036 25288
rect 9088 25276 9094 25288
rect 9815 25279 9873 25285
rect 9815 25276 9827 25279
rect 9088 25248 9827 25276
rect 9088 25236 9094 25248
rect 9815 25245 9827 25248
rect 9861 25245 9873 25279
rect 9815 25239 9873 25245
rect 9950 25276 10008 25282
rect 9950 25242 9962 25276
rect 9996 25242 10008 25276
rect 9950 25236 10008 25242
rect 10042 25236 10048 25288
rect 10100 25285 10106 25288
rect 10100 25276 10108 25285
rect 10229 25279 10287 25285
rect 10100 25248 10145 25276
rect 10100 25239 10108 25248
rect 10229 25245 10241 25279
rect 10275 25276 10287 25279
rect 10962 25276 10968 25288
rect 10275 25248 10968 25276
rect 10275 25245 10287 25248
rect 10229 25239 10287 25245
rect 10100 25236 10106 25239
rect 10962 25236 10968 25248
rect 11020 25236 11026 25288
rect 13814 25236 13820 25288
rect 13872 25276 13878 25288
rect 23106 25285 23112 25288
rect 14829 25279 14887 25285
rect 14829 25276 14841 25279
rect 13872 25248 14841 25276
rect 13872 25236 13878 25248
rect 14829 25245 14841 25248
rect 14875 25245 14887 25279
rect 14829 25239 14887 25245
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25276 18751 25279
rect 23104 25276 23112 25285
rect 18739 25248 22094 25276
rect 23067 25248 23112 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 5534 25208 5540 25220
rect 5495 25180 5540 25208
rect 5534 25168 5540 25180
rect 5592 25168 5598 25220
rect 9582 25140 9588 25152
rect 9543 25112 9588 25140
rect 9582 25100 9588 25112
rect 9640 25100 9646 25152
rect 9965 25140 9993 25236
rect 12428 25211 12486 25217
rect 12428 25177 12440 25211
rect 12474 25208 12486 25211
rect 12618 25208 12624 25220
rect 12474 25180 12624 25208
rect 12474 25177 12486 25180
rect 12428 25171 12486 25177
rect 12618 25168 12624 25180
rect 12676 25168 12682 25220
rect 14734 25168 14740 25220
rect 14792 25208 14798 25220
rect 15074 25211 15132 25217
rect 15074 25208 15086 25211
rect 14792 25180 15086 25208
rect 14792 25168 14798 25180
rect 15074 25177 15086 25180
rect 15120 25177 15132 25211
rect 15074 25171 15132 25177
rect 19512 25211 19570 25217
rect 19512 25177 19524 25211
rect 19558 25177 19570 25211
rect 19512 25171 19570 25177
rect 11054 25140 11060 25152
rect 9965 25112 11060 25140
rect 11054 25100 11060 25112
rect 11112 25140 11118 25152
rect 12158 25140 12164 25152
rect 11112 25112 12164 25140
rect 11112 25100 11118 25112
rect 12158 25100 12164 25112
rect 12216 25140 12222 25152
rect 12710 25140 12716 25152
rect 12216 25112 12716 25140
rect 12216 25100 12222 25112
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 13541 25143 13599 25149
rect 13541 25109 13553 25143
rect 13587 25140 13599 25143
rect 13906 25140 13912 25152
rect 13587 25112 13912 25140
rect 13587 25109 13599 25112
rect 13541 25103 13599 25109
rect 13906 25100 13912 25112
rect 13964 25100 13970 25152
rect 14274 25140 14280 25152
rect 14235 25112 14280 25140
rect 14274 25100 14280 25112
rect 14332 25100 14338 25152
rect 16206 25140 16212 25152
rect 16167 25112 16212 25140
rect 16206 25100 16212 25112
rect 16264 25100 16270 25152
rect 18322 25140 18328 25152
rect 18283 25112 18328 25140
rect 18322 25100 18328 25112
rect 18380 25100 18386 25152
rect 19426 25100 19432 25152
rect 19484 25140 19490 25152
rect 19536 25140 19564 25171
rect 20622 25140 20628 25152
rect 19484 25112 19564 25140
rect 20583 25112 20628 25140
rect 19484 25100 19490 25112
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 22066 25140 22094 25248
rect 23104 25239 23112 25248
rect 23106 25236 23112 25239
rect 23164 25236 23170 25288
rect 23198 25236 23204 25288
rect 23256 25276 23262 25288
rect 23474 25276 23480 25288
rect 23256 25248 23301 25276
rect 23435 25248 23480 25276
rect 23256 25236 23262 25248
rect 23474 25236 23480 25248
rect 23532 25236 23538 25288
rect 23584 25285 23612 25316
rect 27249 25313 27261 25347
rect 27295 25344 27307 25347
rect 28810 25344 28816 25356
rect 27295 25316 28816 25344
rect 27295 25313 27307 25316
rect 27249 25307 27307 25313
rect 28810 25304 28816 25316
rect 28868 25304 28874 25356
rect 29914 25304 29920 25356
rect 29972 25344 29978 25356
rect 29972 25316 30144 25344
rect 29972 25304 29978 25316
rect 23569 25279 23627 25285
rect 23569 25245 23581 25279
rect 23615 25245 23627 25279
rect 24762 25276 24768 25288
rect 24723 25248 24768 25276
rect 23569 25239 23627 25245
rect 24762 25236 24768 25248
rect 24820 25236 24826 25288
rect 24946 25276 24952 25288
rect 24907 25248 24952 25276
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25038 25236 25044 25288
rect 25096 25276 25102 25288
rect 25179 25279 25237 25285
rect 25096 25248 25141 25276
rect 25096 25236 25102 25248
rect 25179 25245 25191 25279
rect 25225 25245 25237 25279
rect 25179 25239 25237 25245
rect 28629 25279 28687 25285
rect 28629 25245 28641 25279
rect 28675 25276 28687 25279
rect 28902 25276 28908 25288
rect 28675 25248 28908 25276
rect 28675 25245 28687 25248
rect 28629 25239 28687 25245
rect 23293 25211 23351 25217
rect 23293 25177 23305 25211
rect 23339 25177 23351 25211
rect 23293 25171 23351 25177
rect 22925 25143 22983 25149
rect 22925 25140 22937 25143
rect 22066 25112 22937 25140
rect 22925 25109 22937 25112
rect 22971 25109 22983 25143
rect 22925 25103 22983 25109
rect 23198 25100 23204 25152
rect 23256 25140 23262 25152
rect 23308 25140 23336 25171
rect 24026 25168 24032 25220
rect 24084 25208 24090 25220
rect 24578 25208 24584 25220
rect 24084 25180 24584 25208
rect 24084 25168 24090 25180
rect 24578 25168 24584 25180
rect 24636 25208 24642 25220
rect 25194 25208 25222 25239
rect 28902 25236 28908 25248
rect 28960 25236 28966 25288
rect 29730 25236 29736 25288
rect 29788 25276 29794 25288
rect 29825 25279 29883 25285
rect 29825 25276 29837 25279
rect 29788 25248 29837 25276
rect 29788 25236 29794 25248
rect 29825 25245 29837 25248
rect 29871 25245 29883 25279
rect 30006 25276 30012 25288
rect 29967 25248 30012 25276
rect 29825 25239 29883 25245
rect 30006 25236 30012 25248
rect 30064 25236 30070 25288
rect 30116 25285 30144 25316
rect 37752 25288 37780 25384
rect 38010 25304 38016 25356
rect 38068 25304 38074 25356
rect 30101 25279 30159 25285
rect 30101 25245 30113 25279
rect 30147 25245 30159 25279
rect 30101 25239 30159 25245
rect 30193 25279 30251 25285
rect 30193 25245 30205 25279
rect 30239 25276 30251 25279
rect 30374 25276 30380 25288
rect 30239 25248 30380 25276
rect 30239 25245 30251 25248
rect 30193 25239 30251 25245
rect 24636 25180 25222 25208
rect 25409 25211 25467 25217
rect 24636 25168 24642 25180
rect 25409 25177 25421 25211
rect 25455 25208 25467 25211
rect 26982 25211 27040 25217
rect 26982 25208 26994 25211
rect 25455 25180 26994 25208
rect 25455 25177 25467 25180
rect 25409 25171 25467 25177
rect 26982 25177 26994 25180
rect 27028 25177 27040 25211
rect 26982 25171 27040 25177
rect 27798 25168 27804 25220
rect 27856 25208 27862 25220
rect 28813 25211 28871 25217
rect 28813 25208 28825 25211
rect 27856 25180 28825 25208
rect 27856 25168 27862 25180
rect 28813 25177 28825 25180
rect 28859 25208 28871 25211
rect 29546 25208 29552 25220
rect 28859 25180 29552 25208
rect 28859 25177 28871 25180
rect 28813 25171 28871 25177
rect 29546 25168 29552 25180
rect 29604 25168 29610 25220
rect 23566 25140 23572 25152
rect 23256 25112 23572 25140
rect 23256 25100 23262 25112
rect 23566 25100 23572 25112
rect 23624 25100 23630 25152
rect 25774 25100 25780 25152
rect 25832 25140 25838 25152
rect 25869 25143 25927 25149
rect 25869 25140 25881 25143
rect 25832 25112 25881 25140
rect 25832 25100 25838 25112
rect 25869 25109 25881 25112
rect 25915 25109 25927 25143
rect 25869 25103 25927 25109
rect 28534 25100 28540 25152
rect 28592 25140 28598 25152
rect 30116 25140 30144 25239
rect 30374 25236 30380 25248
rect 30432 25236 30438 25288
rect 31570 25236 31576 25288
rect 31628 25276 31634 25288
rect 32309 25279 32367 25285
rect 32309 25276 32321 25279
rect 31628 25248 32321 25276
rect 31628 25236 31634 25248
rect 32309 25245 32321 25248
rect 32355 25245 32367 25279
rect 32309 25239 32367 25245
rect 36449 25279 36507 25285
rect 36449 25245 36461 25279
rect 36495 25276 36507 25279
rect 36722 25276 36728 25288
rect 36495 25248 36728 25276
rect 36495 25245 36507 25248
rect 36449 25239 36507 25245
rect 36722 25236 36728 25248
rect 36780 25236 36786 25288
rect 37458 25276 37464 25288
rect 37371 25248 37464 25276
rect 37458 25236 37464 25248
rect 37516 25276 37522 25288
rect 37734 25276 37740 25288
rect 37516 25248 37740 25276
rect 37516 25236 37522 25248
rect 37734 25236 37740 25248
rect 37792 25236 37798 25288
rect 37918 25276 37924 25288
rect 37879 25248 37924 25276
rect 37918 25236 37924 25248
rect 37976 25236 37982 25288
rect 38028 25276 38056 25304
rect 38324 25285 38352 25384
rect 38100 25276 38158 25282
rect 38028 25248 38112 25276
rect 38100 25242 38112 25248
rect 38146 25242 38158 25276
rect 38100 25236 38158 25242
rect 38197 25279 38255 25285
rect 38197 25245 38209 25279
rect 38243 25245 38255 25279
rect 38197 25239 38255 25245
rect 38309 25279 38367 25285
rect 38309 25245 38321 25279
rect 38355 25245 38367 25279
rect 58158 25276 58164 25288
rect 58119 25248 58164 25276
rect 38309 25239 38367 25245
rect 30469 25211 30527 25217
rect 30469 25177 30481 25211
rect 30515 25208 30527 25211
rect 32042 25211 32100 25217
rect 32042 25208 32054 25211
rect 30515 25180 32054 25208
rect 30515 25177 30527 25180
rect 30469 25171 30527 25177
rect 32042 25177 32054 25180
rect 32088 25177 32100 25211
rect 36630 25208 36636 25220
rect 36591 25180 36636 25208
rect 32042 25171 32100 25177
rect 36630 25168 36636 25180
rect 36688 25168 36694 25220
rect 28592 25112 30144 25140
rect 28592 25100 28598 25112
rect 30558 25100 30564 25152
rect 30616 25140 30622 25152
rect 30929 25143 30987 25149
rect 30929 25140 30941 25143
rect 30616 25112 30941 25140
rect 30616 25100 30622 25112
rect 30929 25109 30941 25112
rect 30975 25109 30987 25143
rect 30929 25103 30987 25109
rect 37550 25100 37556 25152
rect 37608 25140 37614 25152
rect 38212 25140 38240 25239
rect 58158 25236 58164 25248
rect 58216 25236 58222 25288
rect 37608 25112 38240 25140
rect 37608 25100 37614 25112
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 2590 24936 2596 24948
rect 2551 24908 2596 24936
rect 2590 24896 2596 24908
rect 2648 24896 2654 24948
rect 12618 24936 12624 24948
rect 12579 24908 12624 24936
rect 12618 24896 12624 24908
rect 12676 24896 12682 24948
rect 14734 24936 14740 24948
rect 14695 24908 14740 24936
rect 14734 24896 14740 24908
rect 14792 24896 14798 24948
rect 15562 24896 15568 24948
rect 15620 24936 15626 24948
rect 16022 24936 16028 24948
rect 15620 24908 16028 24936
rect 15620 24896 15626 24908
rect 16022 24896 16028 24908
rect 16080 24936 16086 24948
rect 16080 24908 19380 24936
rect 16080 24896 16086 24908
rect 2314 24828 2320 24880
rect 2372 24868 2378 24880
rect 8748 24871 8806 24877
rect 2372 24840 4016 24868
rect 2372 24828 2378 24840
rect 3694 24760 3700 24812
rect 3752 24809 3758 24812
rect 3988 24809 4016 24840
rect 8748 24837 8760 24871
rect 8794 24868 8806 24871
rect 9582 24868 9588 24880
rect 8794 24840 9588 24868
rect 8794 24837 8806 24840
rect 8748 24831 8806 24837
rect 9582 24828 9588 24840
rect 9640 24828 9646 24880
rect 10134 24828 10140 24880
rect 10192 24868 10198 24880
rect 11054 24868 11060 24880
rect 10192 24840 10548 24868
rect 10192 24828 10198 24840
rect 3752 24800 3764 24809
rect 3973 24803 4031 24809
rect 3752 24772 3797 24800
rect 3752 24763 3764 24772
rect 3973 24769 3985 24803
rect 4019 24800 4031 24803
rect 5534 24800 5540 24812
rect 4019 24772 5540 24800
rect 4019 24769 4031 24772
rect 3973 24763 4031 24769
rect 3752 24760 3758 24763
rect 5534 24760 5540 24772
rect 5592 24760 5598 24812
rect 6086 24760 6092 24812
rect 6144 24800 6150 24812
rect 10520 24806 10548 24840
rect 10704 24840 11060 24868
rect 10704 24812 10732 24840
rect 11054 24828 11060 24840
rect 11112 24828 11118 24880
rect 12710 24828 12716 24880
rect 12768 24868 12774 24880
rect 16114 24868 16120 24880
rect 12768 24840 16120 24868
rect 12768 24828 12774 24840
rect 10597 24806 10655 24809
rect 10520 24803 10655 24806
rect 6144 24772 9536 24800
rect 10520 24778 10609 24803
rect 6144 24760 6150 24772
rect 6822 24692 6828 24744
rect 6880 24732 6886 24744
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 6880 24704 8493 24732
rect 6880 24692 6886 24704
rect 8481 24701 8493 24704
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 9508 24664 9536 24772
rect 10597 24769 10609 24778
rect 10643 24769 10655 24803
rect 10597 24763 10655 24769
rect 10686 24806 10744 24812
rect 10686 24772 10698 24806
rect 10732 24772 10744 24806
rect 10686 24766 10744 24772
rect 10778 24760 10784 24812
rect 10836 24809 10842 24812
rect 10836 24800 10844 24809
rect 10836 24772 10881 24800
rect 10836 24763 10844 24772
rect 10836 24760 10842 24763
rect 10962 24760 10968 24812
rect 11020 24800 11026 24812
rect 12894 24800 12900 24812
rect 11020 24772 11065 24800
rect 12855 24772 12900 24800
rect 11020 24760 11026 24772
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13004 24809 13032 24840
rect 12989 24803 13047 24809
rect 12989 24769 13001 24803
rect 13035 24769 13047 24803
rect 12989 24763 13047 24769
rect 13078 24760 13084 24812
rect 13136 24800 13142 24812
rect 13136 24772 13181 24800
rect 13136 24760 13142 24772
rect 13262 24760 13268 24812
rect 13320 24800 13326 24812
rect 13320 24772 13365 24800
rect 13320 24760 13326 24772
rect 14182 24760 14188 24812
rect 14240 24800 14246 24812
rect 15120 24809 15148 24840
rect 16114 24828 16120 24840
rect 16172 24828 16178 24880
rect 19352 24868 19380 24908
rect 19426 24896 19432 24948
rect 19484 24936 19490 24948
rect 19521 24939 19579 24945
rect 19521 24936 19533 24939
rect 19484 24908 19533 24936
rect 19484 24896 19490 24908
rect 19521 24905 19533 24908
rect 19567 24905 19579 24939
rect 24762 24936 24768 24948
rect 19521 24899 19579 24905
rect 20088 24908 24768 24936
rect 20088 24868 20116 24908
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 24946 24896 24952 24948
rect 25004 24936 25010 24948
rect 25317 24939 25375 24945
rect 25317 24936 25329 24939
rect 25004 24908 25329 24936
rect 25004 24896 25010 24908
rect 25317 24905 25329 24908
rect 25363 24905 25375 24939
rect 27614 24936 27620 24948
rect 27575 24908 27620 24936
rect 25317 24899 25375 24905
rect 27614 24896 27620 24908
rect 27672 24896 27678 24948
rect 29733 24939 29791 24945
rect 27724 24908 28304 24936
rect 19352 24840 20116 24868
rect 20165 24871 20223 24877
rect 20165 24837 20177 24871
rect 20211 24868 20223 24871
rect 20622 24868 20628 24880
rect 20211 24840 20628 24868
rect 20211 24837 20223 24840
rect 20165 24831 20223 24837
rect 20622 24828 20628 24840
rect 20680 24828 20686 24880
rect 22922 24828 22928 24880
rect 22980 24868 22986 24880
rect 23198 24868 23204 24880
rect 22980 24840 23204 24868
rect 22980 24828 22986 24840
rect 23198 24828 23204 24840
rect 23256 24868 23262 24880
rect 23477 24871 23535 24877
rect 23477 24868 23489 24871
rect 23256 24840 23489 24868
rect 23256 24828 23262 24840
rect 23477 24837 23489 24840
rect 23523 24837 23535 24871
rect 23477 24831 23535 24837
rect 25501 24871 25559 24877
rect 25501 24837 25513 24871
rect 25547 24868 25559 24871
rect 25774 24868 25780 24880
rect 25547 24840 25780 24868
rect 25547 24837 25559 24840
rect 25501 24831 25559 24837
rect 25774 24828 25780 24840
rect 25832 24828 25838 24880
rect 26421 24871 26479 24877
rect 26421 24837 26433 24871
rect 26467 24868 26479 24871
rect 27724 24868 27752 24908
rect 26467 24840 27752 24868
rect 26467 24837 26479 24840
rect 26421 24831 26479 24837
rect 28276 24812 28304 24908
rect 29733 24905 29745 24939
rect 29779 24936 29791 24939
rect 30006 24936 30012 24948
rect 29779 24908 30012 24936
rect 29779 24905 29791 24908
rect 29733 24899 29791 24905
rect 30006 24896 30012 24908
rect 30064 24896 30070 24948
rect 39393 24939 39451 24945
rect 39393 24936 39405 24939
rect 38120 24908 39405 24936
rect 38120 24815 38148 24908
rect 39393 24905 39405 24908
rect 39439 24905 39451 24939
rect 39393 24899 39451 24905
rect 38838 24828 38844 24880
rect 38896 24868 38902 24880
rect 39850 24868 39856 24880
rect 38896 24840 39856 24868
rect 38896 24828 38902 24840
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 14240 24772 15025 24800
rect 14240 24760 14246 24772
rect 15013 24769 15025 24772
rect 15059 24769 15071 24803
rect 15013 24763 15071 24769
rect 15105 24803 15163 24809
rect 15105 24769 15117 24803
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15252 24772 15297 24800
rect 15252 24760 15258 24772
rect 15378 24760 15384 24812
rect 15436 24800 15442 24812
rect 16945 24803 17003 24809
rect 15436 24772 15481 24800
rect 15436 24760 15442 24772
rect 16945 24769 16957 24803
rect 16991 24769 17003 24803
rect 18874 24800 18880 24812
rect 18835 24772 18880 24800
rect 16945 24763 17003 24769
rect 12069 24667 12127 24673
rect 12069 24664 12081 24667
rect 9508 24636 12081 24664
rect 12069 24633 12081 24636
rect 12115 24664 12127 24667
rect 12894 24664 12900 24676
rect 12115 24636 12900 24664
rect 12115 24633 12127 24636
rect 12069 24627 12127 24633
rect 12894 24624 12900 24636
rect 12952 24624 12958 24676
rect 16960 24664 16988 24763
rect 18874 24760 18880 24772
rect 18932 24760 18938 24812
rect 19334 24809 19340 24812
rect 19040 24803 19098 24809
rect 19040 24769 19052 24803
rect 19086 24769 19098 24803
rect 19040 24763 19098 24769
rect 19156 24803 19214 24809
rect 19156 24769 19168 24803
rect 19202 24769 19214 24803
rect 19156 24763 19214 24769
rect 19291 24803 19340 24809
rect 19291 24769 19303 24803
rect 19337 24769 19340 24803
rect 19291 24763 19340 24769
rect 19055 24732 19083 24763
rect 19055 24704 19104 24732
rect 16132 24636 16988 24664
rect 16132 24608 16160 24636
rect 6454 24556 6460 24608
rect 6512 24596 6518 24608
rect 6641 24599 6699 24605
rect 6641 24596 6653 24599
rect 6512 24568 6653 24596
rect 6512 24556 6518 24568
rect 6641 24565 6653 24568
rect 6687 24596 6699 24599
rect 8018 24596 8024 24608
rect 6687 24568 8024 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 8018 24556 8024 24568
rect 8076 24556 8082 24608
rect 9858 24596 9864 24608
rect 9819 24568 9864 24596
rect 9858 24556 9864 24568
rect 9916 24556 9922 24608
rect 10318 24596 10324 24608
rect 10279 24568 10324 24596
rect 10318 24556 10324 24568
rect 10376 24556 10382 24608
rect 11054 24556 11060 24608
rect 11112 24596 11118 24608
rect 11517 24599 11575 24605
rect 11517 24596 11529 24599
rect 11112 24568 11529 24596
rect 11112 24556 11118 24568
rect 11517 24565 11529 24568
rect 11563 24565 11575 24599
rect 14182 24596 14188 24608
rect 14143 24568 14188 24596
rect 11517 24559 11575 24565
rect 14182 24556 14188 24568
rect 14240 24556 14246 24608
rect 16114 24596 16120 24608
rect 16075 24568 16120 24596
rect 16114 24556 16120 24568
rect 16172 24556 16178 24608
rect 16761 24599 16819 24605
rect 16761 24565 16773 24599
rect 16807 24596 16819 24599
rect 17402 24596 17408 24608
rect 16807 24568 17408 24596
rect 16807 24565 16819 24568
rect 16761 24559 16819 24565
rect 17402 24556 17408 24568
rect 17460 24556 17466 24608
rect 19076 24596 19104 24704
rect 19168 24676 19196 24763
rect 19334 24760 19340 24763
rect 19392 24760 19398 24812
rect 20254 24760 20260 24812
rect 20312 24800 20318 24812
rect 20349 24803 20407 24809
rect 20349 24800 20361 24803
rect 20312 24772 20361 24800
rect 20312 24760 20318 24772
rect 20349 24769 20361 24772
rect 20395 24769 20407 24803
rect 20349 24763 20407 24769
rect 22646 24760 22652 24812
rect 22704 24800 22710 24812
rect 23106 24800 23112 24812
rect 22704 24772 23112 24800
rect 22704 24760 22710 24772
rect 23106 24760 23112 24772
rect 23164 24800 23170 24812
rect 23288 24803 23346 24809
rect 23288 24800 23300 24803
rect 23164 24772 23300 24800
rect 23164 24760 23170 24772
rect 23288 24769 23300 24772
rect 23334 24769 23346 24803
rect 23288 24763 23346 24769
rect 23385 24803 23443 24809
rect 23385 24769 23397 24803
rect 23431 24769 23443 24803
rect 23385 24763 23443 24769
rect 23400 24732 23428 24763
rect 23566 24760 23572 24812
rect 23624 24809 23630 24812
rect 23624 24803 23663 24809
rect 23651 24769 23663 24803
rect 23624 24763 23663 24769
rect 23624 24760 23630 24763
rect 23750 24760 23756 24812
rect 23808 24800 23814 24812
rect 24578 24800 24584 24812
rect 23808 24772 23853 24800
rect 24539 24772 24584 24800
rect 23808 24760 23814 24772
rect 24578 24760 24584 24772
rect 24636 24760 24642 24812
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24800 25743 24803
rect 26050 24800 26056 24812
rect 25731 24772 26056 24800
rect 25731 24769 25743 24772
rect 25685 24763 25743 24769
rect 26050 24760 26056 24772
rect 26108 24760 26114 24812
rect 27798 24760 27804 24812
rect 27856 24809 27862 24812
rect 27856 24803 27905 24809
rect 27856 24769 27859 24803
rect 27893 24769 27905 24803
rect 27856 24763 27905 24769
rect 27982 24803 28040 24809
rect 27982 24769 27994 24803
rect 28028 24769 28040 24803
rect 27982 24763 28040 24769
rect 27856 24760 27862 24763
rect 23400 24704 27752 24732
rect 19150 24624 19156 24676
rect 19208 24624 19214 24676
rect 19981 24599 20039 24605
rect 19981 24596 19993 24599
rect 19076 24568 19993 24596
rect 19981 24565 19993 24568
rect 20027 24565 20039 24599
rect 23106 24596 23112 24608
rect 23067 24568 23112 24596
rect 19981 24559 20039 24565
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 27157 24599 27215 24605
rect 27157 24565 27169 24599
rect 27203 24596 27215 24599
rect 27246 24596 27252 24608
rect 27203 24568 27252 24596
rect 27203 24565 27215 24568
rect 27157 24559 27215 24565
rect 27246 24556 27252 24568
rect 27304 24556 27310 24608
rect 27724 24596 27752 24704
rect 27798 24624 27804 24676
rect 27856 24664 27862 24676
rect 28000 24664 28028 24763
rect 28074 24760 28080 24812
rect 28132 24809 28138 24812
rect 28132 24800 28140 24809
rect 28258 24800 28264 24812
rect 28132 24772 28177 24800
rect 28219 24772 28264 24800
rect 28132 24763 28140 24772
rect 28132 24760 28138 24763
rect 28258 24760 28264 24772
rect 28316 24760 28322 24812
rect 28902 24760 28908 24812
rect 28960 24800 28966 24812
rect 29365 24803 29423 24809
rect 29365 24800 29377 24803
rect 28960 24772 29377 24800
rect 28960 24760 28966 24772
rect 29365 24769 29377 24772
rect 29411 24769 29423 24803
rect 29365 24763 29423 24769
rect 29549 24803 29607 24809
rect 29549 24769 29561 24803
rect 29595 24800 29607 24803
rect 30558 24800 30564 24812
rect 29595 24772 30564 24800
rect 29595 24769 29607 24772
rect 29549 24763 29607 24769
rect 29564 24732 29592 24763
rect 30558 24760 30564 24772
rect 30616 24760 30622 24812
rect 30834 24760 30840 24812
rect 30892 24800 30898 24812
rect 31306 24803 31364 24809
rect 31306 24800 31318 24803
rect 30892 24772 31318 24800
rect 30892 24760 30898 24772
rect 31306 24769 31318 24772
rect 31352 24769 31364 24803
rect 31570 24800 31576 24812
rect 31531 24772 31576 24800
rect 31306 24763 31364 24769
rect 31570 24760 31576 24772
rect 31628 24760 31634 24812
rect 33594 24760 33600 24812
rect 33652 24800 33658 24812
rect 34986 24803 35044 24809
rect 34986 24800 34998 24803
rect 33652 24772 34998 24800
rect 33652 24760 33658 24772
rect 34986 24769 34998 24772
rect 35032 24769 35044 24803
rect 34986 24763 35044 24769
rect 37366 24760 37372 24812
rect 37424 24800 37430 24812
rect 37918 24800 37924 24812
rect 37424 24772 37924 24800
rect 37424 24760 37430 24772
rect 37918 24760 37924 24772
rect 37976 24760 37982 24812
rect 38084 24809 38148 24815
rect 38084 24775 38096 24809
rect 38130 24778 38148 24809
rect 38184 24809 38242 24815
rect 38130 24775 38142 24778
rect 38084 24769 38142 24775
rect 38184 24775 38196 24809
rect 38230 24775 38242 24809
rect 38335 24803 38393 24809
rect 38335 24800 38347 24803
rect 38184 24769 38242 24775
rect 38324 24769 38347 24800
rect 38381 24769 38393 24803
rect 39022 24800 39028 24812
rect 38983 24772 39028 24800
rect 27856 24636 28028 24664
rect 28276 24704 29592 24732
rect 35253 24735 35311 24741
rect 27856 24624 27862 24636
rect 28276 24596 28304 24704
rect 35253 24701 35265 24735
rect 35299 24732 35311 24735
rect 37458 24732 37464 24744
rect 35299 24704 37464 24732
rect 35299 24701 35311 24704
rect 35253 24695 35311 24701
rect 37458 24692 37464 24704
rect 37516 24692 37522 24744
rect 33042 24624 33048 24676
rect 33100 24664 33106 24676
rect 33100 24636 34008 24664
rect 33100 24624 33106 24636
rect 27724 24568 28304 24596
rect 28626 24556 28632 24608
rect 28684 24596 28690 24608
rect 28813 24599 28871 24605
rect 28813 24596 28825 24599
rect 28684 24568 28825 24596
rect 28684 24556 28690 24568
rect 28813 24565 28825 24568
rect 28859 24565 28871 24599
rect 28813 24559 28871 24565
rect 29822 24556 29828 24608
rect 29880 24596 29886 24608
rect 30193 24599 30251 24605
rect 30193 24596 30205 24599
rect 29880 24568 30205 24596
rect 29880 24556 29886 24568
rect 30193 24565 30205 24568
rect 30239 24565 30251 24599
rect 33870 24596 33876 24608
rect 33831 24568 33876 24596
rect 30193 24559 30251 24565
rect 33870 24556 33876 24568
rect 33928 24556 33934 24608
rect 33980 24596 34008 24636
rect 37550 24624 37556 24676
rect 37608 24664 37614 24676
rect 38212 24664 38240 24769
rect 37608 24636 38240 24664
rect 38324 24763 38393 24769
rect 37608 24624 37614 24636
rect 37461 24599 37519 24605
rect 37461 24596 37473 24599
rect 33980 24568 37473 24596
rect 37461 24565 37473 24568
rect 37507 24596 37519 24599
rect 38324 24596 38352 24763
rect 39022 24760 39028 24772
rect 39080 24760 39086 24812
rect 39224 24809 39252 24840
rect 39850 24828 39856 24840
rect 39908 24828 39914 24880
rect 39209 24803 39267 24809
rect 39209 24769 39221 24803
rect 39255 24769 39267 24803
rect 39209 24763 39267 24769
rect 38565 24667 38623 24673
rect 38565 24633 38577 24667
rect 38611 24664 38623 24667
rect 38746 24664 38752 24676
rect 38611 24636 38752 24664
rect 38611 24633 38623 24636
rect 38565 24627 38623 24633
rect 38746 24624 38752 24636
rect 38804 24624 38810 24676
rect 40126 24596 40132 24608
rect 37507 24568 40132 24596
rect 37507 24565 37519 24568
rect 37461 24559 37519 24565
rect 40126 24556 40132 24568
rect 40184 24556 40190 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 5810 24392 5816 24404
rect 5723 24364 5816 24392
rect 5810 24352 5816 24364
rect 5868 24392 5874 24404
rect 12526 24392 12532 24404
rect 5868 24364 12532 24392
rect 5868 24352 5874 24364
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 15010 24392 15016 24404
rect 12728 24364 15016 24392
rect 8018 24284 8024 24336
rect 8076 24324 8082 24336
rect 12728 24324 12756 24364
rect 15010 24352 15016 24364
rect 15068 24352 15074 24404
rect 15194 24392 15200 24404
rect 15155 24364 15200 24392
rect 15194 24352 15200 24364
rect 15252 24352 15258 24404
rect 15378 24352 15384 24404
rect 15436 24392 15442 24404
rect 16117 24395 16175 24401
rect 16117 24392 16129 24395
rect 15436 24364 16129 24392
rect 15436 24352 15442 24364
rect 16117 24361 16129 24364
rect 16163 24392 16175 24395
rect 16298 24392 16304 24404
rect 16163 24364 16304 24392
rect 16163 24361 16175 24364
rect 16117 24355 16175 24361
rect 16298 24352 16304 24364
rect 16356 24352 16362 24404
rect 17402 24352 17408 24404
rect 17460 24392 17466 24404
rect 19978 24392 19984 24404
rect 17460 24364 19984 24392
rect 17460 24352 17466 24364
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 21450 24392 21456 24404
rect 21363 24364 21456 24392
rect 21450 24352 21456 24364
rect 21508 24392 21514 24404
rect 21910 24392 21916 24404
rect 21508 24364 21916 24392
rect 21508 24352 21514 24364
rect 21910 24352 21916 24364
rect 21968 24352 21974 24404
rect 24578 24392 24584 24404
rect 22664 24364 24584 24392
rect 13262 24324 13268 24336
rect 8076 24296 12756 24324
rect 12820 24296 13268 24324
rect 8076 24284 8082 24296
rect 5534 24216 5540 24268
rect 5592 24256 5598 24268
rect 6822 24256 6828 24268
rect 5592 24228 6828 24256
rect 5592 24216 5598 24228
rect 6822 24216 6828 24228
rect 6880 24256 6886 24268
rect 7009 24259 7067 24265
rect 7009 24256 7021 24259
rect 6880 24228 7021 24256
rect 6880 24216 6886 24228
rect 7009 24225 7021 24228
rect 7055 24225 7067 24259
rect 10042 24256 10048 24268
rect 10003 24228 10048 24256
rect 7009 24219 7067 24225
rect 10042 24216 10048 24228
rect 10100 24216 10106 24268
rect 6454 24188 6460 24200
rect 6415 24160 6460 24188
rect 6454 24148 6460 24160
rect 6512 24148 6518 24200
rect 7276 24191 7334 24197
rect 7276 24157 7288 24191
rect 7322 24188 7334 24191
rect 10318 24188 10324 24200
rect 7322 24160 10324 24188
rect 7322 24157 7334 24160
rect 7276 24151 7334 24157
rect 10318 24148 10324 24160
rect 10376 24148 10382 24200
rect 11054 24148 11060 24200
rect 11112 24188 11118 24200
rect 12049 24191 12107 24197
rect 12253 24191 12311 24197
rect 12049 24188 12061 24191
rect 11112 24160 12061 24188
rect 11112 24148 11118 24160
rect 12049 24157 12061 24160
rect 12095 24157 12107 24191
rect 12049 24151 12107 24157
rect 12158 24185 12216 24191
rect 12158 24151 12170 24185
rect 12204 24151 12216 24185
rect 12253 24157 12265 24191
rect 12299 24188 12311 24191
rect 12342 24188 12348 24200
rect 12299 24160 12348 24188
rect 12299 24157 12311 24160
rect 12253 24151 12311 24157
rect 12158 24145 12216 24151
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24188 12495 24191
rect 12618 24188 12624 24200
rect 12483 24160 12624 24188
rect 12483 24157 12495 24160
rect 12437 24151 12495 24157
rect 12618 24148 12624 24160
rect 12676 24188 12682 24200
rect 12820 24188 12848 24296
rect 13262 24284 13268 24296
rect 13320 24324 13326 24336
rect 14185 24327 14243 24333
rect 14185 24324 14197 24327
rect 13320 24296 14197 24324
rect 13320 24284 13326 24296
rect 14185 24293 14197 24296
rect 14231 24324 14243 24327
rect 15396 24324 15424 24352
rect 14231 24296 15424 24324
rect 14231 24293 14243 24296
rect 14185 24287 14243 24293
rect 19334 24284 19340 24336
rect 19392 24324 19398 24336
rect 19705 24327 19763 24333
rect 19705 24324 19717 24327
rect 19392 24296 19717 24324
rect 19392 24284 19398 24296
rect 19705 24293 19717 24296
rect 19751 24324 19763 24327
rect 22664 24324 22692 24364
rect 24578 24352 24584 24364
rect 24636 24352 24642 24404
rect 28074 24392 28080 24404
rect 28035 24364 28080 24392
rect 28074 24352 28080 24364
rect 28132 24352 28138 24404
rect 28626 24352 28632 24404
rect 28684 24392 28690 24404
rect 29549 24395 29607 24401
rect 29549 24392 29561 24395
rect 28684 24364 29561 24392
rect 28684 24352 28690 24364
rect 29549 24361 29561 24364
rect 29595 24392 29607 24395
rect 29730 24392 29736 24404
rect 29595 24364 29736 24392
rect 29595 24361 29607 24364
rect 29549 24355 29607 24361
rect 29730 24352 29736 24364
rect 29788 24392 29794 24404
rect 30098 24392 30104 24404
rect 29788 24364 30104 24392
rect 29788 24352 29794 24364
rect 30098 24352 30104 24364
rect 30156 24352 30162 24404
rect 30745 24395 30803 24401
rect 30745 24361 30757 24395
rect 30791 24392 30803 24395
rect 30834 24392 30840 24404
rect 30791 24364 30840 24392
rect 30791 24361 30803 24364
rect 30745 24355 30803 24361
rect 30834 24352 30840 24364
rect 30892 24352 30898 24404
rect 31297 24395 31355 24401
rect 31297 24361 31309 24395
rect 31343 24392 31355 24395
rect 31754 24392 31760 24404
rect 31343 24364 31760 24392
rect 31343 24361 31355 24364
rect 31297 24355 31355 24361
rect 31754 24352 31760 24364
rect 31812 24352 31818 24404
rect 33594 24392 33600 24404
rect 33555 24364 33600 24392
rect 33594 24352 33600 24364
rect 33652 24352 33658 24404
rect 36541 24395 36599 24401
rect 36541 24361 36553 24395
rect 36587 24392 36599 24395
rect 38654 24392 38660 24404
rect 36587 24364 38660 24392
rect 36587 24361 36599 24364
rect 36541 24355 36599 24361
rect 38654 24352 38660 24364
rect 38712 24352 38718 24404
rect 19751 24296 22692 24324
rect 19751 24293 19763 24296
rect 19705 24287 19763 24293
rect 22738 24284 22744 24336
rect 22796 24324 22802 24336
rect 22796 24296 23244 24324
rect 22796 24284 22802 24296
rect 18322 24216 18328 24268
rect 18380 24256 18386 24268
rect 18966 24256 18972 24268
rect 18380 24228 18972 24256
rect 18380 24216 18386 24228
rect 18966 24216 18972 24228
rect 19024 24256 19030 24268
rect 20254 24256 20260 24268
rect 19024 24228 20260 24256
rect 19024 24216 19030 24228
rect 20254 24216 20260 24228
rect 20312 24216 20318 24268
rect 20622 24216 20628 24268
rect 20680 24256 20686 24268
rect 20680 24228 22876 24256
rect 20680 24216 20686 24228
rect 12676 24160 12848 24188
rect 13449 24191 13507 24197
rect 12676 24148 12682 24160
rect 13449 24157 13461 24191
rect 13495 24188 13507 24191
rect 14366 24188 14372 24200
rect 13495 24160 14372 24188
rect 13495 24157 13507 24160
rect 13449 24151 13507 24157
rect 6086 24080 6092 24132
rect 6144 24120 6150 24132
rect 6822 24120 6828 24132
rect 6144 24092 6828 24120
rect 6144 24080 6150 24092
rect 6822 24080 6828 24092
rect 6880 24080 6886 24132
rect 9677 24123 9735 24129
rect 9677 24089 9689 24123
rect 9723 24089 9735 24123
rect 9858 24120 9864 24132
rect 9819 24092 9864 24120
rect 9677 24083 9735 24089
rect 6270 24052 6276 24064
rect 6231 24024 6276 24052
rect 6270 24012 6276 24024
rect 6328 24012 6334 24064
rect 8389 24055 8447 24061
rect 8389 24021 8401 24055
rect 8435 24052 8447 24055
rect 9582 24052 9588 24064
rect 8435 24024 9588 24052
rect 8435 24021 8447 24024
rect 8389 24015 8447 24021
rect 9582 24012 9588 24024
rect 9640 24012 9646 24064
rect 9692 24052 9720 24083
rect 9858 24080 9864 24092
rect 9916 24080 9922 24132
rect 10965 24123 11023 24129
rect 10965 24089 10977 24123
rect 11011 24089 11023 24123
rect 11146 24120 11152 24132
rect 11107 24092 11152 24120
rect 10965 24083 11023 24089
rect 9766 24052 9772 24064
rect 9692 24024 9772 24052
rect 9766 24012 9772 24024
rect 9824 24052 9830 24064
rect 10980 24052 11008 24083
rect 11146 24080 11152 24092
rect 11204 24080 11210 24132
rect 11330 24120 11336 24132
rect 11291 24092 11336 24120
rect 11330 24080 11336 24092
rect 11388 24080 11394 24132
rect 12176 24064 12204 24145
rect 12986 24080 12992 24132
rect 13044 24120 13050 24132
rect 13265 24123 13323 24129
rect 13265 24120 13277 24123
rect 13044 24092 13277 24120
rect 13044 24080 13050 24092
rect 13265 24089 13277 24092
rect 13311 24089 13323 24123
rect 13265 24083 13323 24089
rect 11790 24052 11796 24064
rect 9824 24024 11008 24052
rect 11751 24024 11796 24052
rect 9824 24012 9830 24024
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 12158 24012 12164 24064
rect 12216 24012 12222 24064
rect 12526 24012 12532 24064
rect 12584 24052 12590 24064
rect 13464 24052 13492 24151
rect 14366 24148 14372 24160
rect 14424 24148 14430 24200
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 15470 24188 15476 24200
rect 15427 24160 15476 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 15470 24148 15476 24160
rect 15528 24188 15534 24200
rect 16206 24188 16212 24200
rect 15528 24160 16212 24188
rect 15528 24148 15534 24160
rect 16206 24148 16212 24160
rect 16264 24148 16270 24200
rect 17402 24188 17408 24200
rect 16868 24160 17408 24188
rect 14090 24080 14096 24132
rect 14148 24120 14154 24132
rect 15286 24120 15292 24132
rect 14148 24092 15292 24120
rect 14148 24080 14154 24092
rect 15286 24080 15292 24092
rect 15344 24080 15350 24132
rect 15565 24123 15623 24129
rect 15565 24089 15577 24123
rect 15611 24120 15623 24123
rect 15654 24120 15660 24132
rect 15611 24092 15660 24120
rect 15611 24089 15623 24092
rect 15565 24083 15623 24089
rect 15654 24080 15660 24092
rect 15712 24080 15718 24132
rect 12584 24024 13492 24052
rect 12584 24012 12590 24024
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 14366 24052 14372 24064
rect 13964 24024 14372 24052
rect 13964 24012 13970 24024
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 14734 24052 14740 24064
rect 14695 24024 14740 24052
rect 14734 24012 14740 24024
rect 14792 24012 14798 24064
rect 15010 24012 15016 24064
rect 15068 24052 15074 24064
rect 16868 24052 16896 24160
rect 17402 24148 17408 24160
rect 17460 24148 17466 24200
rect 17586 24188 17592 24200
rect 17547 24160 17592 24188
rect 17586 24148 17592 24160
rect 17644 24148 17650 24200
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24157 17739 24191
rect 17681 24151 17739 24157
rect 17696 24120 17724 24151
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 22646 24188 22652 24200
rect 20036 24160 22652 24188
rect 20036 24148 20042 24160
rect 22646 24148 22652 24160
rect 22704 24197 22710 24200
rect 22704 24191 22753 24197
rect 22704 24157 22707 24191
rect 22741 24157 22753 24191
rect 22848 24188 22876 24228
rect 23216 24197 23244 24296
rect 27246 24256 27252 24268
rect 27159 24228 27252 24256
rect 27246 24216 27252 24228
rect 27304 24256 27310 24268
rect 27706 24256 27712 24268
rect 27304 24228 27712 24256
rect 27304 24216 27310 24228
rect 27706 24216 27712 24228
rect 27764 24256 27770 24268
rect 32493 24259 32551 24265
rect 32493 24256 32505 24259
rect 27764 24228 32505 24256
rect 27764 24216 27770 24228
rect 32493 24225 32505 24228
rect 32539 24256 32551 24259
rect 32766 24256 32772 24268
rect 32539 24228 32772 24256
rect 32539 24225 32551 24228
rect 32493 24219 32551 24225
rect 32766 24216 32772 24228
rect 32824 24256 32830 24268
rect 32824 24228 33364 24256
rect 32824 24216 32830 24228
rect 23053 24191 23111 24197
rect 23053 24188 23065 24191
rect 22848 24160 23065 24188
rect 22704 24151 22753 24157
rect 23053 24157 23065 24160
rect 23099 24157 23111 24191
rect 23053 24151 23111 24157
rect 23201 24191 23259 24197
rect 23201 24157 23213 24191
rect 23247 24157 23259 24191
rect 27890 24188 27896 24200
rect 27851 24160 27896 24188
rect 23201 24151 23259 24157
rect 22704 24148 22710 24151
rect 27890 24148 27896 24160
rect 27948 24148 27954 24200
rect 30098 24188 30104 24200
rect 30059 24160 30104 24188
rect 30098 24148 30104 24160
rect 30156 24148 30162 24200
rect 30282 24188 30288 24200
rect 30243 24160 30288 24188
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 30377 24191 30435 24197
rect 30377 24157 30389 24191
rect 30423 24157 30435 24191
rect 30377 24151 30435 24157
rect 30469 24191 30527 24197
rect 30469 24157 30481 24191
rect 30515 24188 30527 24191
rect 31754 24188 31760 24200
rect 30515 24160 31760 24188
rect 30515 24157 30527 24160
rect 30469 24151 30527 24157
rect 22278 24120 22284 24132
rect 17144 24092 17724 24120
rect 17788 24092 22284 24120
rect 17144 24064 17172 24092
rect 15068 24024 16896 24052
rect 16945 24055 17003 24061
rect 15068 24012 15074 24024
rect 16945 24021 16957 24055
rect 16991 24052 17003 24055
rect 17126 24052 17132 24064
rect 16991 24024 17132 24052
rect 16991 24021 17003 24024
rect 16945 24015 17003 24021
rect 17126 24012 17132 24024
rect 17184 24012 17190 24064
rect 17494 24012 17500 24064
rect 17552 24052 17558 24064
rect 17788 24052 17816 24092
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 22833 24123 22891 24129
rect 22833 24089 22845 24123
rect 22879 24089 22891 24123
rect 22833 24083 22891 24089
rect 17552 24024 17816 24052
rect 17552 24012 17558 24024
rect 19426 24012 19432 24064
rect 19484 24052 19490 24064
rect 22557 24055 22615 24061
rect 22557 24052 22569 24055
rect 19484 24024 22569 24052
rect 19484 24012 19490 24024
rect 22557 24021 22569 24024
rect 22603 24021 22615 24055
rect 22848 24052 22876 24083
rect 22922 24080 22928 24132
rect 22980 24120 22986 24132
rect 26510 24120 26516 24132
rect 22980 24092 23025 24120
rect 26423 24092 26516 24120
rect 22980 24080 22986 24092
rect 26510 24080 26516 24092
rect 26568 24120 26574 24132
rect 27062 24120 27068 24132
rect 26568 24092 27068 24120
rect 26568 24080 26574 24092
rect 27062 24080 27068 24092
rect 27120 24080 27126 24132
rect 27614 24080 27620 24132
rect 27672 24120 27678 24132
rect 27709 24123 27767 24129
rect 27709 24120 27721 24123
rect 27672 24092 27721 24120
rect 27672 24080 27678 24092
rect 27709 24089 27721 24092
rect 27755 24089 27767 24123
rect 27709 24083 27767 24089
rect 27798 24080 27804 24132
rect 27856 24120 27862 24132
rect 28534 24120 28540 24132
rect 27856 24092 28540 24120
rect 27856 24080 27862 24092
rect 28534 24080 28540 24092
rect 28592 24120 28598 24132
rect 30392 24120 30420 24151
rect 28592 24092 30420 24120
rect 31726 24148 31760 24160
rect 31812 24148 31818 24200
rect 31938 24148 31944 24200
rect 31996 24188 32002 24200
rect 32953 24191 33011 24197
rect 32953 24188 32965 24191
rect 31996 24160 32965 24188
rect 31996 24148 32002 24160
rect 32953 24157 32965 24160
rect 32999 24157 33011 24191
rect 33134 24188 33140 24200
rect 33095 24160 33140 24188
rect 32953 24151 33011 24157
rect 33134 24148 33140 24160
rect 33192 24148 33198 24200
rect 33336 24197 33364 24228
rect 36722 24216 36728 24268
rect 36780 24256 36786 24268
rect 39022 24256 39028 24268
rect 36780 24228 39028 24256
rect 36780 24216 36786 24228
rect 39022 24216 39028 24228
rect 39080 24216 39086 24268
rect 33229 24191 33287 24197
rect 33229 24157 33241 24191
rect 33275 24157 33287 24191
rect 33229 24151 33287 24157
rect 33321 24191 33379 24197
rect 33321 24157 33333 24191
rect 33367 24157 33379 24191
rect 33321 24151 33379 24157
rect 31726 24120 31754 24148
rect 33042 24120 33048 24132
rect 31726 24092 33048 24120
rect 28592 24080 28598 24092
rect 33042 24080 33048 24092
rect 33100 24080 33106 24132
rect 33244 24120 33272 24151
rect 38654 24148 38660 24200
rect 38712 24188 38718 24200
rect 38749 24191 38807 24197
rect 38749 24188 38761 24191
rect 38712 24160 38761 24188
rect 38712 24148 38718 24160
rect 38749 24157 38761 24160
rect 38795 24157 38807 24191
rect 58158 24188 58164 24200
rect 58119 24160 58164 24188
rect 38749 24151 38807 24157
rect 58158 24148 58164 24160
rect 58216 24148 58222 24200
rect 33502 24120 33508 24132
rect 33244 24092 33508 24120
rect 33502 24080 33508 24092
rect 33560 24080 33566 24132
rect 29822 24052 29828 24064
rect 22848 24024 29828 24052
rect 22557 24015 22615 24021
rect 29822 24012 29828 24024
rect 29880 24012 29886 24064
rect 37458 24052 37464 24064
rect 37371 24024 37464 24052
rect 37458 24012 37464 24024
rect 37516 24052 37522 24064
rect 37918 24052 37924 24064
rect 37516 24024 37924 24052
rect 37516 24012 37522 24024
rect 37918 24012 37924 24024
rect 37976 24012 37982 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 11146 23808 11152 23860
rect 11204 23848 11210 23860
rect 11517 23851 11575 23857
rect 11517 23848 11529 23851
rect 11204 23820 11529 23848
rect 11204 23808 11210 23820
rect 11517 23817 11529 23820
rect 11563 23848 11575 23851
rect 11606 23848 11612 23860
rect 11563 23820 11612 23848
rect 11563 23817 11575 23820
rect 11517 23811 11575 23817
rect 11606 23808 11612 23820
rect 11664 23808 11670 23860
rect 14090 23848 14096 23860
rect 11716 23820 14096 23848
rect 2685 23783 2743 23789
rect 2685 23749 2697 23783
rect 2731 23780 2743 23783
rect 3513 23783 3571 23789
rect 3513 23780 3525 23783
rect 2731 23752 3525 23780
rect 2731 23749 2743 23752
rect 2685 23743 2743 23749
rect 3513 23749 3525 23752
rect 3559 23780 3571 23783
rect 3786 23780 3792 23792
rect 3559 23752 3792 23780
rect 3559 23749 3571 23752
rect 3513 23743 3571 23749
rect 3786 23740 3792 23752
rect 3844 23780 3850 23792
rect 6270 23780 6276 23792
rect 3844 23752 6276 23780
rect 3844 23740 3850 23752
rect 6270 23740 6276 23752
rect 6328 23740 6334 23792
rect 7745 23783 7803 23789
rect 7745 23780 7757 23783
rect 7208 23752 7757 23780
rect 1854 23672 1860 23724
rect 1912 23712 1918 23724
rect 2501 23715 2559 23721
rect 2501 23712 2513 23715
rect 1912 23684 2513 23712
rect 1912 23672 1918 23684
rect 2501 23681 2513 23684
rect 2547 23681 2559 23715
rect 2501 23675 2559 23681
rect 3329 23715 3387 23721
rect 3329 23681 3341 23715
rect 3375 23712 3387 23715
rect 3418 23712 3424 23724
rect 3375 23684 3424 23712
rect 3375 23681 3387 23684
rect 3329 23675 3387 23681
rect 3418 23672 3424 23684
rect 3476 23672 3482 23724
rect 5810 23712 5816 23724
rect 5771 23684 5816 23712
rect 5810 23672 5816 23684
rect 5868 23672 5874 23724
rect 7208 23721 7236 23752
rect 7745 23749 7757 23752
rect 7791 23780 7803 23783
rect 9953 23783 10011 23789
rect 9953 23780 9965 23783
rect 7791 23752 9965 23780
rect 7791 23749 7803 23752
rect 7745 23743 7803 23749
rect 9953 23749 9965 23752
rect 9999 23780 10011 23783
rect 11716 23780 11744 23820
rect 14090 23808 14096 23820
rect 14148 23808 14154 23860
rect 14734 23848 14740 23860
rect 14292 23820 14740 23848
rect 9999 23752 11744 23780
rect 9999 23749 10011 23752
rect 9953 23743 10011 23749
rect 11790 23740 11796 23792
rect 11848 23780 11854 23792
rect 12630 23783 12688 23789
rect 12630 23780 12642 23783
rect 11848 23752 12642 23780
rect 11848 23740 11854 23752
rect 12630 23749 12642 23752
rect 12676 23749 12688 23783
rect 12630 23743 12688 23749
rect 12986 23740 12992 23792
rect 13044 23780 13050 23792
rect 13357 23783 13415 23789
rect 13357 23780 13369 23783
rect 13044 23752 13369 23780
rect 13044 23740 13050 23752
rect 13357 23749 13369 23752
rect 13403 23749 13415 23783
rect 13357 23743 13415 23749
rect 7193 23715 7251 23721
rect 7193 23681 7205 23715
rect 7239 23681 7251 23715
rect 7193 23675 7251 23681
rect 10137 23715 10195 23721
rect 10137 23681 10149 23715
rect 10183 23681 10195 23715
rect 10137 23675 10195 23681
rect 5537 23647 5595 23653
rect 5537 23613 5549 23647
rect 5583 23644 5595 23647
rect 6362 23644 6368 23656
rect 5583 23616 6368 23644
rect 5583 23613 5595 23616
rect 5537 23607 5595 23613
rect 6362 23604 6368 23616
rect 6420 23604 6426 23656
rect 6914 23644 6920 23656
rect 6875 23616 6920 23644
rect 6914 23604 6920 23616
rect 6972 23604 6978 23656
rect 10152 23644 10180 23675
rect 10318 23672 10324 23724
rect 10376 23712 10382 23724
rect 11698 23712 11704 23724
rect 10376 23684 11704 23712
rect 10376 23672 10382 23684
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23712 12955 23715
rect 13814 23712 13820 23724
rect 12943 23684 13820 23712
rect 12943 23681 12955 23684
rect 12897 23675 12955 23681
rect 13814 23672 13820 23684
rect 13872 23672 13878 23724
rect 14292 23721 14320 23820
rect 14734 23808 14740 23820
rect 14792 23848 14798 23860
rect 17313 23851 17371 23857
rect 17313 23848 17325 23851
rect 14792 23820 17325 23848
rect 14792 23808 14798 23820
rect 14366 23740 14372 23792
rect 14424 23780 14430 23792
rect 15470 23780 15476 23792
rect 14424 23752 14469 23780
rect 14568 23752 15056 23780
rect 15431 23752 15476 23780
rect 14424 23740 14430 23752
rect 14277 23715 14335 23721
rect 14277 23681 14289 23715
rect 14323 23681 14335 23715
rect 14277 23675 14335 23681
rect 14461 23715 14519 23721
rect 14461 23681 14473 23715
rect 14507 23712 14519 23715
rect 14568 23712 14596 23752
rect 14507 23684 14596 23712
rect 14645 23715 14703 23721
rect 14507 23681 14519 23684
rect 14461 23675 14519 23681
rect 14645 23681 14657 23715
rect 14691 23681 14703 23715
rect 14645 23675 14703 23681
rect 10410 23644 10416 23656
rect 10152 23616 10416 23644
rect 10410 23604 10416 23616
rect 10468 23644 10474 23656
rect 10781 23647 10839 23653
rect 10781 23644 10793 23647
rect 10468 23616 10793 23644
rect 10468 23604 10474 23616
rect 10781 23613 10793 23616
rect 10827 23613 10839 23647
rect 14660 23644 14688 23675
rect 15028 23656 15056 23752
rect 15470 23740 15476 23752
rect 15528 23740 15534 23792
rect 15194 23712 15200 23724
rect 15155 23684 15200 23712
rect 15194 23672 15200 23684
rect 15252 23672 15258 23724
rect 15580 23721 15608 23820
rect 17313 23817 17325 23820
rect 17359 23848 17371 23851
rect 17494 23848 17500 23860
rect 17359 23820 17500 23848
rect 17359 23817 17371 23820
rect 17313 23811 17371 23817
rect 17494 23808 17500 23820
rect 17552 23808 17558 23860
rect 17586 23808 17592 23860
rect 17644 23848 17650 23860
rect 19797 23851 19855 23857
rect 19797 23848 19809 23851
rect 17644 23820 19809 23848
rect 17644 23808 17650 23820
rect 19797 23817 19809 23820
rect 19843 23817 19855 23851
rect 19797 23811 19855 23817
rect 20254 23808 20260 23860
rect 20312 23848 20318 23860
rect 21542 23848 21548 23860
rect 20312 23820 21548 23848
rect 20312 23808 20318 23820
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 21726 23808 21732 23860
rect 21784 23848 21790 23860
rect 25133 23851 25191 23857
rect 25133 23848 25145 23851
rect 21784 23820 25145 23848
rect 21784 23808 21790 23820
rect 25133 23817 25145 23820
rect 25179 23848 25191 23851
rect 30009 23851 30067 23857
rect 25179 23820 25820 23848
rect 25179 23817 25191 23820
rect 25133 23811 25191 23817
rect 15654 23740 15660 23792
rect 15712 23780 15718 23792
rect 16114 23780 16120 23792
rect 15712 23752 16120 23780
rect 15712 23740 15718 23752
rect 16114 23740 16120 23752
rect 16172 23780 16178 23792
rect 19058 23780 19064 23792
rect 16172 23752 19064 23780
rect 16172 23740 16178 23752
rect 19058 23740 19064 23752
rect 19116 23740 19122 23792
rect 19889 23783 19947 23789
rect 19889 23749 19901 23783
rect 19935 23780 19947 23783
rect 20162 23780 20168 23792
rect 19935 23752 20168 23780
rect 19935 23749 19947 23752
rect 19889 23743 19947 23749
rect 20162 23740 20168 23752
rect 20220 23780 20226 23792
rect 20438 23780 20444 23792
rect 20220 23752 20444 23780
rect 20220 23740 20226 23752
rect 20438 23740 20444 23752
rect 20496 23740 20502 23792
rect 21821 23783 21879 23789
rect 21821 23780 21833 23783
rect 20824 23752 21833 23780
rect 15381 23715 15439 23721
rect 15381 23681 15393 23715
rect 15427 23681 15439 23715
rect 15381 23675 15439 23681
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23681 15623 23715
rect 15565 23675 15623 23681
rect 18141 23715 18199 23721
rect 18141 23681 18153 23715
rect 18187 23712 18199 23715
rect 18966 23712 18972 23724
rect 18187 23684 18972 23712
rect 18187 23681 18199 23684
rect 18141 23675 18199 23681
rect 10781 23607 10839 23613
rect 13280 23616 14688 23644
rect 2317 23579 2375 23585
rect 2317 23545 2329 23579
rect 2363 23576 2375 23579
rect 3326 23576 3332 23588
rect 2363 23548 3332 23576
rect 2363 23545 2375 23548
rect 2317 23539 2375 23545
rect 3326 23536 3332 23548
rect 3384 23536 3390 23588
rect 7466 23536 7472 23588
rect 7524 23576 7530 23588
rect 7524 23548 10916 23576
rect 7524 23536 7530 23548
rect 3142 23508 3148 23520
rect 3103 23480 3148 23508
rect 3142 23468 3148 23480
rect 3200 23468 3206 23520
rect 10888 23508 10916 23548
rect 13280 23508 13308 23616
rect 15010 23604 15016 23656
rect 15068 23644 15074 23656
rect 15396 23644 15424 23675
rect 18966 23672 18972 23684
rect 19024 23672 19030 23724
rect 20824 23721 20852 23752
rect 21821 23749 21833 23752
rect 21867 23749 21879 23783
rect 21821 23743 21879 23749
rect 22005 23783 22063 23789
rect 22005 23749 22017 23783
rect 22051 23780 22063 23783
rect 23382 23780 23388 23792
rect 22051 23752 23388 23780
rect 22051 23749 22063 23752
rect 22005 23743 22063 23749
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 25792 23789 25820 23820
rect 30009 23817 30021 23851
rect 30055 23848 30067 23851
rect 30282 23848 30288 23860
rect 30055 23820 30288 23848
rect 30055 23817 30067 23820
rect 30009 23811 30067 23817
rect 30282 23808 30288 23820
rect 30340 23808 30346 23860
rect 39301 23851 39359 23857
rect 39301 23848 39313 23851
rect 36556 23820 39313 23848
rect 25777 23783 25835 23789
rect 25777 23749 25789 23783
rect 25823 23749 25835 23783
rect 25777 23743 25835 23749
rect 27338 23740 27344 23792
rect 27396 23780 27402 23792
rect 27709 23783 27767 23789
rect 27709 23780 27721 23783
rect 27396 23752 27721 23780
rect 27396 23740 27402 23752
rect 27709 23749 27721 23752
rect 27755 23749 27767 23783
rect 29822 23780 29828 23792
rect 29783 23752 29828 23780
rect 27709 23743 27767 23749
rect 29822 23740 29828 23752
rect 29880 23740 29886 23792
rect 35710 23740 35716 23792
rect 35768 23780 35774 23792
rect 36556 23789 36584 23820
rect 39301 23817 39313 23820
rect 39347 23817 39359 23851
rect 39301 23811 39359 23817
rect 36541 23783 36599 23789
rect 36541 23780 36553 23783
rect 35768 23752 36553 23780
rect 35768 23740 35774 23752
rect 36541 23749 36553 23752
rect 36587 23749 36599 23783
rect 36541 23743 36599 23749
rect 20625 23715 20683 23721
rect 20625 23712 20637 23715
rect 19306 23684 20637 23712
rect 15068 23616 16804 23644
rect 15068 23604 15074 23616
rect 16776 23585 16804 23616
rect 18874 23604 18880 23656
rect 18932 23644 18938 23656
rect 19306 23644 19334 23684
rect 20625 23681 20637 23684
rect 20671 23681 20683 23715
rect 20625 23675 20683 23681
rect 20809 23715 20867 23721
rect 20809 23681 20821 23715
rect 20855 23681 20867 23715
rect 20809 23675 20867 23681
rect 20901 23715 20959 23721
rect 20901 23681 20913 23715
rect 20947 23681 20959 23715
rect 20901 23675 20959 23681
rect 20993 23715 21051 23721
rect 20993 23681 21005 23715
rect 21039 23712 21051 23715
rect 21450 23712 21456 23724
rect 21039 23684 21456 23712
rect 21039 23681 21051 23684
rect 20993 23675 21051 23681
rect 18932 23616 19334 23644
rect 18932 23604 18938 23616
rect 16761 23579 16819 23585
rect 16761 23545 16773 23579
rect 16807 23576 16819 23579
rect 16807 23548 18460 23576
rect 16807 23545 16819 23548
rect 16761 23539 16819 23545
rect 14090 23508 14096 23520
rect 10888 23480 13308 23508
rect 14051 23480 14096 23508
rect 14090 23468 14096 23480
rect 14148 23468 14154 23520
rect 15470 23468 15476 23520
rect 15528 23508 15534 23520
rect 15749 23511 15807 23517
rect 15749 23508 15761 23511
rect 15528 23480 15761 23508
rect 15528 23468 15534 23480
rect 15749 23477 15761 23480
rect 15795 23477 15807 23511
rect 18322 23508 18328 23520
rect 18283 23480 18328 23508
rect 15749 23471 15807 23477
rect 18322 23468 18328 23480
rect 18380 23468 18386 23520
rect 18432 23508 18460 23548
rect 19150 23536 19156 23588
rect 19208 23576 19214 23588
rect 20916 23576 20944 23675
rect 21450 23672 21456 23684
rect 21508 23672 21514 23724
rect 21542 23672 21548 23724
rect 21600 23712 21606 23724
rect 22189 23715 22247 23721
rect 22189 23712 22201 23715
rect 21600 23684 22201 23712
rect 21600 23672 21606 23684
rect 22189 23681 22201 23684
rect 22235 23712 22247 23715
rect 24394 23712 24400 23724
rect 22235 23684 24400 23712
rect 22235 23681 22247 23684
rect 22189 23675 22247 23681
rect 24394 23672 24400 23684
rect 24452 23672 24458 23724
rect 27525 23715 27583 23721
rect 27525 23681 27537 23715
rect 27571 23712 27583 23715
rect 27614 23712 27620 23724
rect 27571 23684 27620 23712
rect 27571 23681 27583 23684
rect 27525 23675 27583 23681
rect 27614 23672 27620 23684
rect 27672 23712 27678 23724
rect 28902 23712 28908 23724
rect 27672 23684 28908 23712
rect 27672 23672 27678 23684
rect 28902 23672 28908 23684
rect 28960 23712 28966 23724
rect 29641 23715 29699 23721
rect 29641 23712 29653 23715
rect 28960 23684 29653 23712
rect 28960 23672 28966 23684
rect 29641 23681 29653 23684
rect 29687 23681 29699 23715
rect 29641 23675 29699 23681
rect 33226 23672 33232 23724
rect 33284 23712 33290 23724
rect 33974 23715 34032 23721
rect 33974 23712 33986 23715
rect 33284 23684 33986 23712
rect 33284 23672 33290 23684
rect 33974 23681 33986 23684
rect 34020 23681 34032 23715
rect 33974 23675 34032 23681
rect 36357 23715 36415 23721
rect 36357 23681 36369 23715
rect 36403 23712 36415 23715
rect 36722 23712 36728 23724
rect 36403 23684 36728 23712
rect 36403 23681 36415 23684
rect 36357 23675 36415 23681
rect 36722 23672 36728 23684
rect 36780 23672 36786 23724
rect 38194 23721 38200 23724
rect 38188 23675 38200 23721
rect 38252 23712 38258 23724
rect 38252 23684 38288 23712
rect 38194 23672 38200 23675
rect 38252 23672 38258 23684
rect 21468 23644 21496 23672
rect 24486 23644 24492 23656
rect 21468 23616 24492 23644
rect 24486 23604 24492 23616
rect 24544 23604 24550 23656
rect 34241 23647 34299 23653
rect 34241 23613 34253 23647
rect 34287 23644 34299 23647
rect 37918 23644 37924 23656
rect 34287 23616 37924 23644
rect 34287 23613 34299 23616
rect 34241 23607 34299 23613
rect 37918 23604 37924 23616
rect 37976 23604 37982 23656
rect 19208 23548 20944 23576
rect 21269 23579 21327 23585
rect 19208 23536 19214 23548
rect 21269 23545 21281 23579
rect 21315 23576 21327 23579
rect 22094 23576 22100 23588
rect 21315 23548 22100 23576
rect 21315 23545 21327 23548
rect 21269 23539 21327 23545
rect 22094 23536 22100 23548
rect 22152 23536 22158 23588
rect 25961 23579 26019 23585
rect 25961 23545 25973 23579
rect 26007 23576 26019 23579
rect 26510 23576 26516 23588
rect 26007 23548 26516 23576
rect 26007 23545 26019 23548
rect 25961 23539 26019 23545
rect 26510 23536 26516 23548
rect 26568 23576 26574 23588
rect 31938 23576 31944 23588
rect 26568 23548 31944 23576
rect 26568 23536 26574 23548
rect 31938 23536 31944 23548
rect 31996 23536 32002 23588
rect 22462 23508 22468 23520
rect 18432 23480 22468 23508
rect 22462 23468 22468 23480
rect 22520 23468 22526 23520
rect 27893 23511 27951 23517
rect 27893 23477 27905 23511
rect 27939 23508 27951 23511
rect 28166 23508 28172 23520
rect 27939 23480 28172 23508
rect 27939 23477 27951 23480
rect 27893 23471 27951 23477
rect 28166 23468 28172 23480
rect 28224 23468 28230 23520
rect 32306 23468 32312 23520
rect 32364 23508 32370 23520
rect 32861 23511 32919 23517
rect 32861 23508 32873 23511
rect 32364 23480 32873 23508
rect 32364 23468 32370 23480
rect 32861 23477 32873 23480
rect 32907 23477 32919 23511
rect 32861 23471 32919 23477
rect 36725 23511 36783 23517
rect 36725 23477 36737 23511
rect 36771 23508 36783 23511
rect 37642 23508 37648 23520
rect 36771 23480 37648 23508
rect 36771 23477 36783 23480
rect 36725 23471 36783 23477
rect 37642 23468 37648 23480
rect 37700 23468 37706 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 6914 23304 6920 23316
rect 4817 23276 6920 23304
rect 2682 23196 2688 23248
rect 2740 23236 2746 23248
rect 3881 23239 3939 23245
rect 3881 23236 3893 23239
rect 2740 23208 3893 23236
rect 2740 23196 2746 23208
rect 3881 23205 3893 23208
rect 3927 23236 3939 23239
rect 4706 23236 4712 23248
rect 3927 23208 4712 23236
rect 3927 23205 3939 23208
rect 3881 23199 3939 23205
rect 4706 23196 4712 23208
rect 4764 23196 4770 23248
rect 2700 23097 2728 23196
rect 3602 23168 3608 23180
rect 2976 23140 3608 23168
rect 2976 23109 3004 23140
rect 3602 23128 3608 23140
rect 3660 23168 3666 23180
rect 4817 23168 4845 23276
rect 6914 23264 6920 23276
rect 6972 23264 6978 23316
rect 12618 23304 12624 23316
rect 12579 23276 12624 23304
rect 12618 23264 12624 23276
rect 12676 23264 12682 23316
rect 15010 23304 15016 23316
rect 14971 23276 15016 23304
rect 15010 23264 15016 23276
rect 15068 23264 15074 23316
rect 22922 23304 22928 23316
rect 19306 23276 22928 23304
rect 7282 23196 7288 23248
rect 7340 23236 7346 23248
rect 12158 23236 12164 23248
rect 7340 23208 12164 23236
rect 7340 23196 7346 23208
rect 12158 23196 12164 23208
rect 12216 23196 12222 23248
rect 15194 23236 15200 23248
rect 12406 23208 15200 23236
rect 5442 23168 5448 23180
rect 3660 23140 4845 23168
rect 3660 23128 3666 23140
rect 2869 23103 2927 23109
rect 2700 23094 2774 23097
rect 2869 23094 2881 23103
rect 2700 23069 2881 23094
rect 2915 23069 2927 23103
rect 2746 23066 2927 23069
rect 2869 23063 2927 23066
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23069 3019 23103
rect 2961 23063 3019 23069
rect 3053 23100 3111 23106
rect 3053 23066 3065 23100
rect 3099 23066 3111 23100
rect 3053 23060 3111 23066
rect 3237 23103 3295 23109
rect 3237 23069 3249 23103
rect 3283 23100 3295 23103
rect 3510 23100 3516 23112
rect 3283 23072 3516 23100
rect 3283 23069 3295 23072
rect 3237 23063 3295 23069
rect 3510 23060 3516 23072
rect 3568 23100 3574 23112
rect 4817 23109 4845 23140
rect 4908 23140 5448 23168
rect 4908 23109 4936 23140
rect 5442 23128 5448 23140
rect 5500 23128 5506 23180
rect 5534 23128 5540 23180
rect 5592 23168 5598 23180
rect 5629 23171 5687 23177
rect 5629 23168 5641 23171
rect 5592 23140 5641 23168
rect 5592 23128 5598 23140
rect 5629 23137 5641 23140
rect 5675 23137 5687 23171
rect 12406 23168 12434 23208
rect 15194 23196 15200 23208
rect 15252 23196 15258 23248
rect 15930 23236 15936 23248
rect 15396 23208 15936 23236
rect 5629 23131 5687 23137
rect 9048 23140 12434 23168
rect 4525 23103 4583 23109
rect 4525 23100 4537 23103
rect 3568 23072 4537 23100
rect 3568 23060 3574 23072
rect 4525 23069 4537 23072
rect 4571 23100 4583 23103
rect 4709 23103 4767 23109
rect 4571 23072 4660 23100
rect 4571 23069 4583 23072
rect 4525 23063 4583 23069
rect 3068 23032 3096 23060
rect 3142 23032 3148 23044
rect 3068 23004 3148 23032
rect 3142 22992 3148 23004
rect 3200 22992 3206 23044
rect 2593 22967 2651 22973
rect 2593 22933 2605 22967
rect 2639 22964 2651 22967
rect 2682 22964 2688 22976
rect 2639 22936 2688 22964
rect 2639 22933 2651 22936
rect 2593 22927 2651 22933
rect 2682 22924 2688 22936
rect 2740 22924 2746 22976
rect 4632 22964 4660 23072
rect 4709 23069 4721 23103
rect 4755 23069 4767 23103
rect 4709 23063 4767 23069
rect 4801 23103 4859 23109
rect 4801 23069 4813 23103
rect 4847 23069 4859 23103
rect 4801 23063 4859 23069
rect 4893 23103 4951 23109
rect 4893 23069 4905 23103
rect 4939 23069 4951 23103
rect 7837 23103 7895 23109
rect 7837 23100 7849 23103
rect 4893 23063 4951 23069
rect 5000 23072 7849 23100
rect 4724 23032 4752 23063
rect 5000 23032 5028 23072
rect 7837 23069 7849 23072
rect 7883 23069 7895 23103
rect 7837 23063 7895 23069
rect 4724 23004 5028 23032
rect 5169 23035 5227 23041
rect 5169 23001 5181 23035
rect 5215 23032 5227 23035
rect 5874 23035 5932 23041
rect 5874 23032 5886 23035
rect 5215 23004 5886 23032
rect 5215 23001 5227 23004
rect 5169 22995 5227 23001
rect 5874 23001 5886 23004
rect 5920 23001 5932 23035
rect 5874 22995 5932 23001
rect 6270 22992 6276 23044
rect 6328 23032 6334 23044
rect 7469 23035 7527 23041
rect 7469 23032 7481 23035
rect 6328 23004 7481 23032
rect 6328 22992 6334 23004
rect 7469 23001 7481 23004
rect 7515 23001 7527 23035
rect 7469 22995 7527 23001
rect 7653 23035 7711 23041
rect 7653 23001 7665 23035
rect 7699 23032 7711 23035
rect 9048 23032 9076 23140
rect 9766 23060 9772 23112
rect 9824 23100 9830 23112
rect 11517 23103 11575 23109
rect 11517 23100 11529 23103
rect 9824 23072 11529 23100
rect 9824 23060 9830 23072
rect 11517 23069 11529 23072
rect 11563 23069 11575 23103
rect 11517 23063 11575 23069
rect 7699 23004 9076 23032
rect 7699 23001 7711 23004
rect 7653 22995 7711 23001
rect 6362 22964 6368 22976
rect 4632 22936 6368 22964
rect 6362 22924 6368 22936
rect 6420 22924 6426 22976
rect 7009 22967 7067 22973
rect 7009 22933 7021 22967
rect 7055 22964 7067 22967
rect 7668 22964 7696 22995
rect 7055 22936 7696 22964
rect 7055 22933 7067 22936
rect 7009 22927 7067 22933
rect 11238 22924 11244 22976
rect 11296 22964 11302 22976
rect 11333 22967 11391 22973
rect 11333 22964 11345 22967
rect 11296 22936 11345 22964
rect 11296 22924 11302 22936
rect 11333 22933 11345 22936
rect 11379 22933 11391 22967
rect 11532 22964 11560 23063
rect 11606 23060 11612 23112
rect 11664 23100 11670 23112
rect 11664 23072 11709 23100
rect 11664 23060 11670 23072
rect 11790 23060 11796 23112
rect 11848 23100 11854 23112
rect 11885 23103 11943 23109
rect 11885 23100 11897 23103
rect 11848 23072 11897 23100
rect 11848 23060 11854 23072
rect 11885 23069 11897 23072
rect 11931 23069 11943 23103
rect 15396 23100 15424 23208
rect 15930 23196 15936 23208
rect 15988 23196 15994 23248
rect 19306 23236 19334 23276
rect 22922 23264 22928 23276
rect 22980 23264 22986 23316
rect 24486 23304 24492 23316
rect 24447 23276 24492 23304
rect 24486 23264 24492 23276
rect 24544 23304 24550 23316
rect 25038 23304 25044 23316
rect 24544 23276 25044 23304
rect 24544 23264 24550 23276
rect 25038 23264 25044 23276
rect 25096 23264 25102 23316
rect 29546 23304 29552 23316
rect 27724 23276 29552 23304
rect 17144 23208 19334 23236
rect 17144 23177 17172 23208
rect 21266 23196 21272 23248
rect 21324 23236 21330 23248
rect 23106 23236 23112 23248
rect 21324 23208 23112 23236
rect 21324 23196 21330 23208
rect 23106 23196 23112 23208
rect 23164 23196 23170 23248
rect 17129 23171 17187 23177
rect 17129 23168 17141 23171
rect 15764 23140 17141 23168
rect 11885 23063 11943 23069
rect 11992 23072 15424 23100
rect 11698 23032 11704 23044
rect 11659 23004 11704 23032
rect 11698 22992 11704 23004
rect 11756 22992 11762 23044
rect 11992 22964 12020 23072
rect 15470 23060 15476 23112
rect 15528 23100 15534 23112
rect 15654 23109 15660 23112
rect 15621 23103 15660 23109
rect 15528 23072 15573 23100
rect 15528 23060 15534 23072
rect 15621 23069 15633 23103
rect 15621 23063 15660 23069
rect 15654 23060 15660 23063
rect 15712 23060 15718 23112
rect 15764 23109 15792 23140
rect 17129 23137 17141 23140
rect 17175 23137 17187 23171
rect 17129 23131 17187 23137
rect 18141 23171 18199 23177
rect 18141 23137 18153 23171
rect 18187 23168 18199 23171
rect 19150 23168 19156 23180
rect 18187 23140 19156 23168
rect 18187 23137 18199 23140
rect 18141 23131 18199 23137
rect 19150 23128 19156 23140
rect 19208 23128 19214 23180
rect 19797 23171 19855 23177
rect 19797 23137 19809 23171
rect 19843 23168 19855 23171
rect 20254 23168 20260 23180
rect 19843 23140 20260 23168
rect 19843 23137 19855 23140
rect 19797 23131 19855 23137
rect 20254 23128 20260 23140
rect 20312 23128 20318 23180
rect 27724 23168 27752 23276
rect 29546 23264 29552 23276
rect 29604 23264 29610 23316
rect 33134 23264 33140 23316
rect 33192 23304 33198 23316
rect 33505 23307 33563 23313
rect 33505 23304 33517 23307
rect 33192 23276 33517 23304
rect 33192 23264 33198 23276
rect 33505 23273 33517 23276
rect 33551 23273 33563 23307
rect 33505 23267 33563 23273
rect 38105 23307 38163 23313
rect 38105 23273 38117 23307
rect 38151 23304 38163 23307
rect 38194 23304 38200 23316
rect 38151 23276 38200 23304
rect 38151 23273 38163 23276
rect 38105 23267 38163 23273
rect 38194 23264 38200 23276
rect 38252 23264 38258 23316
rect 32677 23239 32735 23245
rect 32677 23205 32689 23239
rect 32723 23236 32735 23239
rect 33226 23236 33232 23248
rect 32723 23208 33232 23236
rect 32723 23205 32735 23208
rect 32677 23199 32735 23205
rect 33226 23196 33232 23208
rect 33284 23196 33290 23248
rect 22756 23140 27752 23168
rect 28721 23171 28779 23177
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 15979 23103 16037 23109
rect 15979 23069 15991 23103
rect 16025 23100 16037 23103
rect 17402 23100 17408 23112
rect 16025 23072 17264 23100
rect 17363 23072 17408 23100
rect 16025 23069 16037 23072
rect 15979 23063 16037 23069
rect 12158 22992 12164 23044
rect 12216 23032 12222 23044
rect 14182 23032 14188 23044
rect 12216 23004 14188 23032
rect 12216 22992 12222 23004
rect 14182 22992 14188 23004
rect 14240 22992 14246 23044
rect 15838 22992 15844 23044
rect 15896 23032 15902 23044
rect 17236 23032 17264 23072
rect 17402 23060 17408 23072
rect 17460 23060 17466 23112
rect 17770 23060 17776 23112
rect 17828 23100 17834 23112
rect 17865 23103 17923 23109
rect 17865 23100 17877 23103
rect 17828 23072 17877 23100
rect 17828 23060 17834 23072
rect 17865 23069 17877 23072
rect 17911 23069 17923 23103
rect 17865 23063 17923 23069
rect 20073 23103 20131 23109
rect 20073 23069 20085 23103
rect 20119 23069 20131 23103
rect 22756 23100 22784 23140
rect 28721 23137 28733 23171
rect 28767 23168 28779 23171
rect 28810 23168 28816 23180
rect 28767 23140 28816 23168
rect 28767 23137 28779 23140
rect 28721 23131 28779 23137
rect 28810 23128 28816 23140
rect 28868 23128 28874 23180
rect 32766 23128 32772 23180
rect 32824 23168 32830 23180
rect 36081 23171 36139 23177
rect 32824 23140 34008 23168
rect 32824 23128 32830 23140
rect 20073 23063 20131 23069
rect 20824 23072 22784 23100
rect 22833 23103 22891 23109
rect 19978 23032 19984 23044
rect 15896 23004 15941 23032
rect 17236 23004 19984 23032
rect 15896 22992 15902 23004
rect 19978 22992 19984 23004
rect 20036 23032 20042 23044
rect 20088 23032 20116 23063
rect 20036 23004 20116 23032
rect 20036 22992 20042 23004
rect 20254 22992 20260 23044
rect 20312 23032 20318 23044
rect 20438 23032 20444 23044
rect 20312 23004 20444 23032
rect 20312 22992 20318 23004
rect 20438 22992 20444 23004
rect 20496 22992 20502 23044
rect 20530 22992 20536 23044
rect 20588 23032 20594 23044
rect 20824 23032 20852 23072
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 30742 23100 30748 23112
rect 22879 23072 30748 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 20588 23004 20852 23032
rect 20588 22992 20594 23004
rect 20898 22992 20904 23044
rect 20956 23032 20962 23044
rect 21085 23035 21143 23041
rect 21085 23032 21097 23035
rect 20956 23004 21097 23032
rect 20956 22992 20962 23004
rect 21085 23001 21097 23004
rect 21131 23001 21143 23035
rect 21085 22995 21143 23001
rect 16114 22964 16120 22976
rect 11532 22936 12020 22964
rect 16075 22936 16120 22964
rect 11333 22927 11391 22933
rect 16114 22924 16120 22936
rect 16172 22924 16178 22976
rect 17218 22924 17224 22976
rect 17276 22964 17282 22976
rect 22370 22964 22376 22976
rect 17276 22936 22376 22964
rect 17276 22924 17282 22936
rect 22370 22924 22376 22936
rect 22428 22964 22434 22976
rect 22848 22964 22876 23063
rect 30742 23060 30748 23072
rect 30800 23060 30806 23112
rect 31938 23060 31944 23112
rect 31996 23100 32002 23112
rect 32033 23103 32091 23109
rect 32033 23100 32045 23103
rect 31996 23072 32045 23100
rect 31996 23060 32002 23072
rect 32033 23069 32045 23072
rect 32079 23069 32091 23103
rect 32033 23063 32091 23069
rect 32122 23060 32128 23112
rect 32180 23100 32186 23112
rect 32217 23103 32275 23109
rect 32217 23100 32229 23103
rect 32180 23072 32229 23100
rect 32180 23060 32186 23072
rect 32217 23069 32229 23072
rect 32263 23069 32275 23103
rect 32217 23063 32275 23069
rect 32309 23103 32367 23109
rect 32309 23069 32321 23103
rect 32355 23069 32367 23103
rect 32309 23063 32367 23069
rect 32401 23103 32459 23109
rect 32401 23069 32413 23103
rect 32447 23069 32459 23103
rect 33318 23100 33324 23112
rect 33231 23072 33324 23100
rect 32401 23063 32459 23069
rect 27706 22992 27712 23044
rect 27764 23032 27770 23044
rect 28454 23035 28512 23041
rect 28454 23032 28466 23035
rect 27764 23004 28466 23032
rect 27764 22992 27770 23004
rect 28454 23001 28466 23004
rect 28500 23001 28512 23035
rect 28454 22995 28512 23001
rect 31662 22992 31668 23044
rect 31720 23032 31726 23044
rect 32324 23032 32352 23063
rect 31720 23004 32352 23032
rect 31720 22992 31726 23004
rect 27338 22964 27344 22976
rect 22428 22936 22876 22964
rect 27299 22936 27344 22964
rect 22428 22924 22434 22936
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 30282 22924 30288 22976
rect 30340 22964 30346 22976
rect 31481 22967 31539 22973
rect 31481 22964 31493 22967
rect 30340 22936 31493 22964
rect 30340 22924 30346 22936
rect 31481 22933 31493 22936
rect 31527 22964 31539 22967
rect 32416 22964 32444 23063
rect 33318 23060 33324 23072
rect 33376 23100 33382 23112
rect 33870 23100 33876 23112
rect 33376 23072 33876 23100
rect 33376 23060 33382 23072
rect 33870 23060 33876 23072
rect 33928 23060 33934 23112
rect 33980 23100 34008 23140
rect 36081 23137 36093 23171
rect 36127 23168 36139 23171
rect 37918 23168 37924 23180
rect 36127 23140 37924 23168
rect 36127 23137 36139 23140
rect 36081 23131 36139 23137
rect 37918 23128 37924 23140
rect 37976 23128 37982 23180
rect 33980 23072 37044 23100
rect 32490 22992 32496 23044
rect 32548 23032 32554 23044
rect 33137 23035 33195 23041
rect 33137 23032 33149 23035
rect 32548 23004 33149 23032
rect 32548 22992 32554 23004
rect 33137 23001 33149 23004
rect 33183 23001 33195 23035
rect 33137 22995 33195 23001
rect 33686 22992 33692 23044
rect 33744 23032 33750 23044
rect 35814 23035 35872 23041
rect 35814 23032 35826 23035
rect 33744 23004 35826 23032
rect 33744 22992 33750 23004
rect 35814 23001 35826 23004
rect 35860 23001 35872 23035
rect 35814 22995 35872 23001
rect 34698 22964 34704 22976
rect 31527 22936 32444 22964
rect 34659 22936 34704 22964
rect 31527 22933 31539 22936
rect 31481 22927 31539 22933
rect 34698 22924 34704 22936
rect 34756 22924 34762 22976
rect 37016 22973 37044 23072
rect 37366 23060 37372 23112
rect 37424 23100 37430 23112
rect 37461 23103 37519 23109
rect 37461 23100 37473 23103
rect 37424 23072 37473 23100
rect 37424 23060 37430 23072
rect 37461 23069 37473 23072
rect 37507 23069 37519 23103
rect 37642 23100 37648 23112
rect 37603 23072 37648 23100
rect 37461 23063 37519 23069
rect 37642 23060 37648 23072
rect 37700 23060 37706 23112
rect 37737 23103 37795 23109
rect 37737 23069 37749 23103
rect 37783 23069 37795 23103
rect 37737 23063 37795 23069
rect 37829 23103 37887 23109
rect 37829 23069 37841 23103
rect 37875 23100 37887 23103
rect 39666 23100 39672 23112
rect 37875 23072 39672 23100
rect 37875 23069 37887 23072
rect 37829 23063 37887 23069
rect 37550 22992 37556 23044
rect 37608 23032 37614 23044
rect 37752 23032 37780 23063
rect 37608 23004 37780 23032
rect 37608 22992 37614 23004
rect 37001 22967 37059 22973
rect 37001 22933 37013 22967
rect 37047 22964 37059 22967
rect 37844 22964 37872 23063
rect 39666 23060 39672 23072
rect 39724 23060 39730 23112
rect 37047 22936 37872 22964
rect 37047 22933 37059 22936
rect 37001 22927 37059 22933
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 6270 22760 6276 22772
rect 3620 22732 4384 22760
rect 3620 22704 3648 22732
rect 3602 22692 3608 22704
rect 3252 22664 3608 22692
rect 3252 22633 3280 22664
rect 3602 22652 3608 22664
rect 3660 22652 3666 22704
rect 4356 22692 4384 22732
rect 4264 22664 4384 22692
rect 5460 22732 6276 22760
rect 4264 22636 4292 22664
rect 3145 22627 3203 22633
rect 3145 22593 3157 22627
rect 3191 22593 3203 22627
rect 3145 22587 3203 22593
rect 3234 22627 3292 22633
rect 3234 22593 3246 22627
rect 3280 22593 3292 22627
rect 3234 22587 3292 22593
rect 3160 22556 3188 22587
rect 3326 22584 3332 22636
rect 3384 22624 3390 22636
rect 3384 22596 3429 22624
rect 3384 22584 3390 22596
rect 3510 22584 3516 22636
rect 3568 22624 3574 22636
rect 3973 22627 4031 22633
rect 3973 22624 3985 22627
rect 3568 22596 3985 22624
rect 3568 22584 3574 22596
rect 3973 22593 3985 22596
rect 4019 22593 4031 22627
rect 4136 22627 4194 22633
rect 4136 22624 4148 22627
rect 3973 22587 4031 22593
rect 4080 22596 4148 22624
rect 3694 22556 3700 22568
rect 2746 22528 3700 22556
rect 2409 22491 2467 22497
rect 2409 22457 2421 22491
rect 2455 22488 2467 22491
rect 2746 22488 2774 22528
rect 3694 22516 3700 22528
rect 3752 22556 3758 22568
rect 3878 22556 3884 22568
rect 3752 22528 3884 22556
rect 3752 22516 3758 22528
rect 3878 22516 3884 22528
rect 3936 22516 3942 22568
rect 4080 22500 4108 22596
rect 4136 22593 4148 22596
rect 4182 22593 4194 22627
rect 4136 22587 4194 22593
rect 4252 22630 4310 22636
rect 4252 22596 4264 22630
rect 4298 22596 4310 22630
rect 4252 22590 4310 22596
rect 4341 22627 4399 22633
rect 4341 22593 4353 22627
rect 4387 22624 4399 22627
rect 4706 22624 4712 22636
rect 4387 22596 4712 22624
rect 4387 22593 4399 22596
rect 4341 22587 4399 22593
rect 4706 22584 4712 22596
rect 4764 22624 4770 22636
rect 4982 22624 4988 22636
rect 4764 22596 4988 22624
rect 4764 22584 4770 22596
rect 4982 22584 4988 22596
rect 5040 22584 5046 22636
rect 5460 22633 5488 22732
rect 6270 22720 6276 22732
rect 6328 22720 6334 22772
rect 10318 22760 10324 22772
rect 9600 22732 10324 22760
rect 9306 22652 9312 22704
rect 9364 22692 9370 22704
rect 9600 22701 9628 22732
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 17402 22760 17408 22772
rect 15252 22732 17408 22760
rect 15252 22720 15258 22732
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 20257 22763 20315 22769
rect 20257 22729 20269 22763
rect 20303 22729 20315 22763
rect 27338 22760 27344 22772
rect 20257 22723 20315 22729
rect 20548 22732 27344 22760
rect 9585 22695 9643 22701
rect 9585 22692 9597 22695
rect 9364 22664 9597 22692
rect 9364 22652 9370 22664
rect 9585 22661 9597 22664
rect 9631 22661 9643 22695
rect 9585 22655 9643 22661
rect 9677 22695 9735 22701
rect 9677 22661 9689 22695
rect 9723 22692 9735 22695
rect 9858 22692 9864 22704
rect 9723 22664 9864 22692
rect 9723 22661 9735 22664
rect 9677 22655 9735 22661
rect 9858 22652 9864 22664
rect 9916 22652 9922 22704
rect 5445 22627 5503 22633
rect 5445 22593 5457 22627
rect 5491 22593 5503 22627
rect 5445 22587 5503 22593
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22593 5687 22627
rect 6362 22624 6368 22636
rect 6323 22596 6368 22624
rect 5629 22587 5687 22593
rect 2455 22460 2774 22488
rect 2455 22457 2467 22460
rect 2409 22451 2467 22457
rect 4062 22448 4068 22500
rect 4120 22448 4126 22500
rect 5644 22488 5672 22587
rect 6362 22584 6368 22596
rect 6420 22584 6426 22636
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 6644 22627 6702 22633
rect 6644 22593 6656 22627
rect 6690 22593 6702 22627
rect 6644 22587 6702 22593
rect 6779 22627 6837 22633
rect 6779 22593 6791 22627
rect 6825 22624 6837 22627
rect 7098 22624 7104 22636
rect 6825 22596 7104 22624
rect 6825 22593 6837 22596
rect 6779 22587 6837 22593
rect 5813 22559 5871 22565
rect 5813 22525 5825 22559
rect 5859 22556 5871 22559
rect 6564 22556 6592 22587
rect 5859 22528 6592 22556
rect 6656 22556 6684 22587
rect 7098 22584 7104 22596
rect 7156 22584 7162 22636
rect 9398 22624 9404 22636
rect 9359 22596 9404 22624
rect 9398 22584 9404 22596
rect 9456 22584 9462 22636
rect 9766 22624 9772 22636
rect 9727 22596 9772 22624
rect 9766 22584 9772 22596
rect 9824 22584 9830 22636
rect 11514 22584 11520 22636
rect 11572 22624 11578 22636
rect 16114 22624 16120 22636
rect 11572 22596 16120 22624
rect 11572 22584 11578 22596
rect 16114 22584 16120 22596
rect 16172 22584 16178 22636
rect 6914 22556 6920 22568
rect 6656 22528 6920 22556
rect 5859 22525 5871 22528
rect 5813 22519 5871 22525
rect 6914 22516 6920 22528
rect 6972 22516 6978 22568
rect 7466 22516 7472 22568
rect 7524 22516 7530 22568
rect 12250 22516 12256 22568
rect 12308 22556 12314 22568
rect 17218 22556 17224 22568
rect 12308 22528 17224 22556
rect 12308 22516 12314 22528
rect 17218 22516 17224 22528
rect 17276 22516 17282 22568
rect 7484 22488 7512 22516
rect 5644 22460 7512 22488
rect 13906 22448 13912 22500
rect 13964 22488 13970 22500
rect 17420 22488 17448 22720
rect 19613 22627 19671 22633
rect 19613 22593 19625 22627
rect 19659 22624 19671 22627
rect 20272 22624 20300 22723
rect 20548 22701 20576 22732
rect 27338 22720 27344 22732
rect 27396 22720 27402 22772
rect 27706 22760 27712 22772
rect 27667 22732 27712 22760
rect 27706 22720 27712 22732
rect 27764 22720 27770 22772
rect 29270 22720 29276 22772
rect 29328 22760 29334 22772
rect 29457 22763 29515 22769
rect 29457 22760 29469 22763
rect 29328 22732 29469 22760
rect 29328 22720 29334 22732
rect 29457 22729 29469 22732
rect 29503 22760 29515 22763
rect 32122 22760 32128 22772
rect 29503 22732 30144 22760
rect 32083 22732 32128 22760
rect 29503 22729 29515 22732
rect 29457 22723 29515 22729
rect 22094 22701 22100 22704
rect 20533 22695 20591 22701
rect 20533 22661 20545 22695
rect 20579 22661 20591 22695
rect 20533 22655 20591 22661
rect 22088 22655 22100 22701
rect 22152 22692 22158 22704
rect 24762 22692 24768 22704
rect 22152 22664 22188 22692
rect 24688 22664 24768 22692
rect 22094 22652 22100 22655
rect 22152 22652 22158 22664
rect 20438 22633 20444 22636
rect 20436 22624 20444 22633
rect 19659 22596 20300 22624
rect 20399 22596 20444 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 20436 22587 20444 22596
rect 20438 22584 20444 22587
rect 20496 22584 20502 22636
rect 20625 22627 20683 22633
rect 20625 22593 20637 22627
rect 20671 22593 20683 22627
rect 20625 22587 20683 22593
rect 19521 22559 19579 22565
rect 19521 22525 19533 22559
rect 19567 22556 19579 22559
rect 20530 22556 20536 22568
rect 19567 22528 20536 22556
rect 19567 22525 19579 22528
rect 19521 22519 19579 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 20640 22488 20668 22587
rect 20714 22584 20720 22636
rect 20772 22633 20778 22636
rect 20772 22627 20811 22633
rect 20799 22593 20811 22627
rect 20772 22587 20811 22593
rect 20901 22627 20959 22633
rect 20901 22593 20913 22627
rect 20947 22624 20959 22627
rect 20990 22624 20996 22636
rect 20947 22596 20996 22624
rect 20947 22593 20959 22596
rect 20901 22587 20959 22593
rect 20772 22584 20778 22587
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 21634 22584 21640 22636
rect 21692 22624 21698 22636
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21692 22596 21833 22624
rect 21692 22584 21698 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 23842 22624 23848 22636
rect 23803 22596 23848 22624
rect 21821 22587 21879 22593
rect 23842 22584 23848 22596
rect 23900 22584 23906 22636
rect 24688 22633 24716 22664
rect 24762 22652 24768 22664
rect 24820 22652 24826 22704
rect 25961 22695 26019 22701
rect 25961 22661 25973 22695
rect 26007 22692 26019 22695
rect 26326 22692 26332 22704
rect 26007 22664 26332 22692
rect 26007 22661 26019 22664
rect 25961 22655 26019 22661
rect 26326 22652 26332 22664
rect 26384 22652 26390 22704
rect 30116 22701 30144 22732
rect 32122 22720 32128 22732
rect 32180 22720 32186 22772
rect 33686 22760 33692 22772
rect 33647 22732 33692 22760
rect 33686 22720 33692 22732
rect 33744 22720 33750 22772
rect 30101 22695 30159 22701
rect 30101 22661 30113 22695
rect 30147 22661 30159 22695
rect 30101 22655 30159 22661
rect 31726 22664 31892 22692
rect 24673 22627 24731 22633
rect 24673 22593 24685 22627
rect 24719 22593 24731 22627
rect 24854 22624 24860 22636
rect 24815 22596 24860 22624
rect 24673 22587 24731 22593
rect 24854 22584 24860 22596
rect 24912 22584 24918 22636
rect 24952 22627 25010 22633
rect 24952 22593 24964 22627
rect 24998 22593 25010 22627
rect 24952 22587 25010 22593
rect 24964 22500 24992 22587
rect 25038 22584 25044 22636
rect 25096 22624 25102 22636
rect 25096 22596 25141 22624
rect 25096 22584 25102 22596
rect 26050 22584 26056 22636
rect 26108 22624 26114 22636
rect 26145 22627 26203 22633
rect 27985 22627 28043 22633
rect 26145 22624 26157 22627
rect 26108 22596 26157 22624
rect 26108 22584 26114 22596
rect 26145 22593 26157 22596
rect 26191 22593 26203 22627
rect 27908 22624 27997 22627
rect 26145 22587 26203 22593
rect 27724 22599 27997 22624
rect 27724 22596 27936 22599
rect 13964 22460 16252 22488
rect 17420 22460 20668 22488
rect 23124 22460 23796 22488
rect 13964 22448 13970 22460
rect 2869 22423 2927 22429
rect 2869 22389 2881 22423
rect 2915 22420 2927 22423
rect 2958 22420 2964 22432
rect 2915 22392 2964 22420
rect 2915 22389 2927 22392
rect 2869 22383 2927 22389
rect 2958 22380 2964 22392
rect 3016 22380 3022 22432
rect 4614 22420 4620 22432
rect 4575 22392 4620 22420
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 7006 22420 7012 22432
rect 6967 22392 7012 22420
rect 7006 22380 7012 22392
rect 7064 22380 7070 22432
rect 7098 22380 7104 22432
rect 7156 22420 7162 22432
rect 7558 22420 7564 22432
rect 7156 22392 7564 22420
rect 7156 22380 7162 22392
rect 7558 22380 7564 22392
rect 7616 22380 7622 22432
rect 9950 22420 9956 22432
rect 9911 22392 9956 22420
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 16025 22423 16083 22429
rect 16025 22389 16037 22423
rect 16071 22420 16083 22423
rect 16114 22420 16120 22432
rect 16071 22392 16120 22420
rect 16071 22389 16083 22392
rect 16025 22383 16083 22389
rect 16114 22380 16120 22392
rect 16172 22380 16178 22432
rect 16224 22420 16252 22460
rect 18874 22420 18880 22432
rect 16224 22392 18880 22420
rect 18874 22380 18880 22392
rect 18932 22380 18938 22432
rect 19242 22420 19248 22432
rect 19203 22392 19248 22420
rect 19242 22380 19248 22392
rect 19300 22380 19306 22432
rect 19613 22423 19671 22429
rect 19613 22389 19625 22423
rect 19659 22420 19671 22423
rect 20070 22420 20076 22432
rect 19659 22392 20076 22420
rect 19659 22389 19671 22392
rect 19613 22383 19671 22389
rect 20070 22380 20076 22392
rect 20128 22380 20134 22432
rect 20346 22380 20352 22432
rect 20404 22420 20410 22432
rect 23124 22420 23152 22460
rect 20404 22392 23152 22420
rect 23201 22423 23259 22429
rect 20404 22380 20410 22392
rect 23201 22389 23213 22423
rect 23247 22420 23259 22423
rect 23382 22420 23388 22432
rect 23247 22392 23388 22420
rect 23247 22389 23259 22392
rect 23201 22383 23259 22389
rect 23382 22380 23388 22392
rect 23440 22380 23446 22432
rect 23768 22429 23796 22460
rect 24946 22448 24952 22500
rect 25004 22448 25010 22500
rect 25038 22448 25044 22500
rect 25096 22488 25102 22500
rect 25777 22491 25835 22497
rect 25777 22488 25789 22491
rect 25096 22460 25789 22488
rect 25096 22448 25102 22460
rect 25777 22457 25789 22460
rect 25823 22457 25835 22491
rect 25777 22451 25835 22457
rect 27062 22448 27068 22500
rect 27120 22488 27126 22500
rect 27522 22488 27528 22500
rect 27120 22460 27528 22488
rect 27120 22448 27126 22460
rect 27522 22448 27528 22460
rect 27580 22448 27586 22500
rect 23753 22423 23811 22429
rect 23753 22389 23765 22423
rect 23799 22420 23811 22423
rect 25130 22420 25136 22432
rect 23799 22392 25136 22420
rect 23799 22389 23811 22392
rect 23753 22383 23811 22389
rect 25130 22380 25136 22392
rect 25188 22380 25194 22432
rect 25314 22420 25320 22432
rect 25275 22392 25320 22420
rect 25314 22380 25320 22392
rect 25372 22380 25378 22432
rect 27249 22423 27307 22429
rect 27249 22389 27261 22423
rect 27295 22420 27307 22423
rect 27338 22420 27344 22432
rect 27295 22392 27344 22420
rect 27295 22389 27307 22392
rect 27249 22383 27307 22389
rect 27338 22380 27344 22392
rect 27396 22420 27402 22432
rect 27724 22420 27752 22596
rect 27985 22593 27997 22599
rect 28031 22593 28043 22627
rect 27985 22587 28043 22593
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 27798 22516 27804 22568
rect 27856 22556 27862 22568
rect 28092 22556 28120 22587
rect 28166 22584 28172 22636
rect 28224 22624 28230 22636
rect 28224 22596 28269 22624
rect 28224 22584 28230 22596
rect 28350 22584 28356 22636
rect 28408 22624 28414 22636
rect 28408 22596 28453 22624
rect 28408 22584 28414 22596
rect 31726 22556 31754 22664
rect 27856 22528 28120 22556
rect 28184 22528 31754 22556
rect 31864 22556 31892 22664
rect 32030 22652 32036 22704
rect 32088 22692 32094 22704
rect 32306 22692 32312 22704
rect 32088 22664 32312 22692
rect 32088 22652 32094 22664
rect 32306 22652 32312 22664
rect 32364 22652 32370 22704
rect 32490 22692 32496 22704
rect 32451 22664 32496 22692
rect 32490 22652 32496 22664
rect 32548 22652 32554 22704
rect 33134 22652 33140 22704
rect 33192 22692 33198 22704
rect 33502 22692 33508 22704
rect 33192 22664 33508 22692
rect 33192 22652 33198 22664
rect 31938 22584 31944 22636
rect 31996 22624 32002 22636
rect 33045 22627 33103 22633
rect 33045 22624 33057 22627
rect 31996 22596 33057 22624
rect 31996 22584 32002 22596
rect 33045 22593 33057 22596
rect 33091 22593 33103 22627
rect 33226 22624 33232 22636
rect 33187 22596 33232 22624
rect 33045 22587 33103 22593
rect 33226 22584 33232 22596
rect 33284 22584 33290 22636
rect 33336 22633 33364 22664
rect 33502 22652 33508 22664
rect 33560 22652 33566 22704
rect 33321 22627 33379 22633
rect 33321 22593 33333 22627
rect 33367 22593 33379 22627
rect 33321 22587 33379 22593
rect 33413 22627 33471 22633
rect 33413 22593 33425 22627
rect 33459 22593 33471 22627
rect 33413 22587 33471 22593
rect 31864 22528 33272 22556
rect 27856 22516 27862 22528
rect 28184 22420 28212 22528
rect 29270 22448 29276 22500
rect 29328 22488 29334 22500
rect 30282 22488 30288 22500
rect 29328 22460 30288 22488
rect 29328 22448 29334 22460
rect 30282 22448 30288 22460
rect 30340 22448 30346 22500
rect 31662 22448 31668 22500
rect 31720 22488 31726 22500
rect 33134 22488 33140 22500
rect 31720 22460 33140 22488
rect 31720 22448 31726 22460
rect 33134 22448 33140 22460
rect 33192 22448 33198 22500
rect 33244 22488 33272 22528
rect 33428 22488 33456 22587
rect 37918 22584 37924 22636
rect 37976 22624 37982 22636
rect 38657 22627 38715 22633
rect 38657 22624 38669 22627
rect 37976 22596 38669 22624
rect 37976 22584 37982 22596
rect 38657 22593 38669 22596
rect 38703 22593 38715 22627
rect 38657 22587 38715 22593
rect 38924 22627 38982 22633
rect 38924 22593 38936 22627
rect 38970 22624 38982 22627
rect 39850 22624 39856 22636
rect 38970 22596 39856 22624
rect 38970 22593 38982 22596
rect 38924 22587 38982 22593
rect 39850 22584 39856 22596
rect 39908 22584 39914 22636
rect 33502 22488 33508 22500
rect 33244 22460 33508 22488
rect 33502 22448 33508 22460
rect 33560 22448 33566 22500
rect 40126 22448 40132 22500
rect 40184 22488 40190 22500
rect 40497 22491 40555 22497
rect 40497 22488 40509 22491
rect 40184 22460 40509 22488
rect 40184 22448 40190 22460
rect 40497 22457 40509 22460
rect 40543 22457 40555 22491
rect 58158 22488 58164 22500
rect 58119 22460 58164 22488
rect 40497 22451 40555 22457
rect 58158 22448 58164 22460
rect 58216 22448 58222 22500
rect 27396 22392 28212 22420
rect 27396 22380 27402 22392
rect 38654 22380 38660 22432
rect 38712 22420 38718 22432
rect 40037 22423 40095 22429
rect 40037 22420 40049 22423
rect 38712 22392 40049 22420
rect 38712 22380 38718 22392
rect 40037 22389 40049 22392
rect 40083 22420 40095 22423
rect 40218 22420 40224 22432
rect 40083 22392 40224 22420
rect 40083 22389 40095 22392
rect 40037 22383 40095 22389
rect 40218 22380 40224 22392
rect 40276 22380 40282 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 4062 22176 4068 22228
rect 4120 22216 4126 22228
rect 4157 22219 4215 22225
rect 4157 22216 4169 22219
rect 4120 22188 4169 22216
rect 4120 22176 4126 22188
rect 4157 22185 4169 22188
rect 4203 22185 4215 22219
rect 4157 22179 4215 22185
rect 5353 22219 5411 22225
rect 5353 22185 5365 22219
rect 5399 22216 5411 22219
rect 5534 22216 5540 22228
rect 5399 22188 5540 22216
rect 5399 22185 5411 22188
rect 5353 22179 5411 22185
rect 5534 22176 5540 22188
rect 5592 22176 5598 22228
rect 6730 22176 6736 22228
rect 6788 22216 6794 22228
rect 7282 22216 7288 22228
rect 6788 22188 7288 22216
rect 6788 22176 6794 22188
rect 7282 22176 7288 22188
rect 7340 22176 7346 22228
rect 7466 22216 7472 22228
rect 7427 22188 7472 22216
rect 7466 22176 7472 22188
rect 7524 22176 7530 22228
rect 14642 22176 14648 22228
rect 14700 22216 14706 22228
rect 15654 22216 15660 22228
rect 14700 22188 15240 22216
rect 15615 22188 15660 22216
rect 14700 22176 14706 22188
rect 15212 22148 15240 22188
rect 15654 22176 15660 22188
rect 15712 22176 15718 22228
rect 16942 22176 16948 22228
rect 17000 22216 17006 22228
rect 17126 22216 17132 22228
rect 17000 22188 17132 22216
rect 17000 22176 17006 22188
rect 17126 22176 17132 22188
rect 17184 22176 17190 22228
rect 18506 22216 18512 22228
rect 18467 22188 18512 22216
rect 18506 22176 18512 22188
rect 18564 22176 18570 22228
rect 18782 22176 18788 22228
rect 18840 22216 18846 22228
rect 19429 22219 19487 22225
rect 19429 22216 19441 22219
rect 18840 22188 19441 22216
rect 18840 22176 18846 22188
rect 19429 22185 19441 22188
rect 19475 22185 19487 22219
rect 19429 22179 19487 22185
rect 22462 22176 22468 22228
rect 22520 22216 22526 22228
rect 22520 22188 27200 22216
rect 22520 22176 22526 22188
rect 21266 22148 21272 22160
rect 15212 22120 21272 22148
rect 21266 22108 21272 22120
rect 21324 22108 21330 22160
rect 26326 22148 26332 22160
rect 26239 22120 26332 22148
rect 26326 22108 26332 22120
rect 26384 22148 26390 22160
rect 27062 22148 27068 22160
rect 26384 22120 27068 22148
rect 26384 22108 26390 22120
rect 27062 22108 27068 22120
rect 27120 22108 27126 22160
rect 27172 22148 27200 22188
rect 28350 22176 28356 22228
rect 28408 22216 28414 22228
rect 29733 22219 29791 22225
rect 29733 22216 29745 22219
rect 28408 22188 29745 22216
rect 28408 22176 28414 22188
rect 29733 22185 29745 22188
rect 29779 22185 29791 22219
rect 39850 22216 39856 22228
rect 39811 22188 39856 22216
rect 29733 22179 29791 22185
rect 39850 22176 39856 22188
rect 39908 22176 39914 22228
rect 41325 22219 41383 22225
rect 41325 22216 41337 22219
rect 39960 22188 41337 22216
rect 29362 22148 29368 22160
rect 27172 22120 29368 22148
rect 29362 22108 29368 22120
rect 29420 22108 29426 22160
rect 29546 22148 29552 22160
rect 29507 22120 29552 22148
rect 29546 22108 29552 22120
rect 29604 22108 29610 22160
rect 33594 22148 33600 22160
rect 30024 22120 33600 22148
rect 13814 22040 13820 22092
rect 13872 22080 13878 22092
rect 14277 22083 14335 22089
rect 14277 22080 14289 22083
rect 13872 22052 14289 22080
rect 13872 22040 13878 22052
rect 14277 22049 14289 22052
rect 14323 22049 14335 22083
rect 14277 22043 14335 22049
rect 19521 22083 19579 22089
rect 19521 22049 19533 22083
rect 19567 22080 19579 22083
rect 20530 22080 20536 22092
rect 19567 22052 20536 22080
rect 19567 22049 19579 22052
rect 19521 22043 19579 22049
rect 2958 22012 2964 22024
rect 3016 22021 3022 22024
rect 2928 21984 2964 22012
rect 2958 21972 2964 21984
rect 3016 21975 3028 22021
rect 3237 22015 3295 22021
rect 3237 21981 3249 22015
rect 3283 22012 3295 22015
rect 4246 22012 4252 22024
rect 3283 21984 4252 22012
rect 3283 21981 3295 21984
rect 3237 21975 3295 21981
rect 3016 21972 3022 21975
rect 4246 21972 4252 21984
rect 4304 22012 4310 22024
rect 6089 22015 6147 22021
rect 6089 22012 6101 22015
rect 4304 21984 6101 22012
rect 4304 21972 4310 21984
rect 6089 21981 6101 21984
rect 6135 22012 6147 22015
rect 7742 22012 7748 22024
rect 6135 21984 7748 22012
rect 6135 21981 6147 21984
rect 6089 21975 6147 21981
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 9217 22015 9275 22021
rect 9217 21981 9229 22015
rect 9263 21981 9275 22015
rect 9217 21975 9275 21981
rect 3786 21944 3792 21956
rect 3747 21916 3792 21944
rect 3786 21904 3792 21916
rect 3844 21904 3850 21956
rect 3970 21944 3976 21956
rect 3931 21916 3976 21944
rect 3970 21904 3976 21916
rect 4028 21904 4034 21956
rect 6356 21947 6414 21953
rect 4080 21916 5028 21944
rect 1854 21876 1860 21888
rect 1815 21848 1860 21876
rect 1854 21836 1860 21848
rect 1912 21836 1918 21888
rect 3418 21836 3424 21888
rect 3476 21876 3482 21888
rect 3878 21876 3884 21888
rect 3476 21848 3884 21876
rect 3476 21836 3482 21848
rect 3878 21836 3884 21848
rect 3936 21876 3942 21888
rect 4080 21876 4108 21916
rect 4706 21876 4712 21888
rect 3936 21848 4108 21876
rect 4667 21848 4712 21876
rect 3936 21836 3942 21848
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 5000 21876 5028 21916
rect 6356 21913 6368 21947
rect 6402 21944 6414 21947
rect 7006 21944 7012 21956
rect 6402 21916 7012 21944
rect 6402 21913 6414 21916
rect 6356 21907 6414 21913
rect 7006 21904 7012 21916
rect 7064 21904 7070 21956
rect 9232 21876 9260 21975
rect 9306 21972 9312 22024
rect 9364 22012 9370 22024
rect 9401 22015 9459 22021
rect 9401 22012 9413 22015
rect 9364 21984 9413 22012
rect 9364 21972 9370 21984
rect 9401 21981 9413 21984
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 9585 22015 9643 22021
rect 9585 21981 9597 22015
rect 9631 22012 9643 22015
rect 9766 22012 9772 22024
rect 9631 21984 9772 22012
rect 9631 21981 9643 21984
rect 9585 21975 9643 21981
rect 9766 21972 9772 21984
rect 9824 21972 9830 22024
rect 14292 22012 14320 22043
rect 20530 22040 20536 22052
rect 20588 22040 20594 22092
rect 22002 22040 22008 22092
rect 22060 22080 22066 22092
rect 24397 22083 24455 22089
rect 24397 22080 24409 22083
rect 22060 22052 24409 22080
rect 22060 22040 22066 22052
rect 24397 22049 24409 22052
rect 24443 22049 24455 22083
rect 29914 22080 29920 22092
rect 24397 22043 24455 22049
rect 29748 22052 29920 22080
rect 17681 22015 17739 22021
rect 17681 22012 17693 22015
rect 14292 21984 17693 22012
rect 17681 21981 17693 21984
rect 17727 22012 17739 22015
rect 18138 22012 18144 22024
rect 17727 21984 18144 22012
rect 17727 21981 17739 21984
rect 17681 21975 17739 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 18598 22012 18604 22024
rect 18559 21984 18604 22012
rect 18598 21972 18604 21984
rect 18656 21972 18662 22024
rect 18693 22015 18751 22021
rect 18693 21981 18705 22015
rect 18739 21981 18751 22015
rect 18693 21975 18751 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 22012 19671 22015
rect 22186 22012 22192 22024
rect 19659 21984 22192 22012
rect 19659 21981 19671 21984
rect 19613 21975 19671 21981
rect 9493 21947 9551 21953
rect 9493 21913 9505 21947
rect 9539 21944 9551 21947
rect 9674 21944 9680 21956
rect 9539 21916 9680 21944
rect 9539 21913 9551 21916
rect 9493 21907 9551 21913
rect 9674 21904 9680 21916
rect 9732 21904 9738 21956
rect 14550 21953 14556 21956
rect 14544 21907 14556 21953
rect 14608 21944 14614 21956
rect 16114 21944 16120 21956
rect 14608 21916 14644 21944
rect 16075 21916 16120 21944
rect 14550 21904 14556 21907
rect 14608 21904 14614 21916
rect 16114 21904 16120 21916
rect 16172 21904 16178 21956
rect 18708 21944 18736 21975
rect 22186 21972 22192 21984
rect 22244 21972 22250 22024
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 22012 25007 22015
rect 26234 22012 26240 22024
rect 24995 21984 26240 22012
rect 24995 21981 25007 21984
rect 24949 21975 25007 21981
rect 26234 21972 26240 21984
rect 26292 21972 26298 22024
rect 29748 22021 29776 22052
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 30024 22021 30052 22120
rect 33594 22108 33600 22120
rect 33652 22108 33658 22160
rect 39114 22148 39120 22160
rect 39037 22120 39120 22148
rect 30374 22040 30380 22092
rect 30432 22080 30438 22092
rect 30745 22083 30803 22089
rect 30745 22080 30757 22083
rect 30432 22052 30757 22080
rect 30432 22040 30438 22052
rect 30745 22049 30757 22052
rect 30791 22080 30803 22083
rect 31018 22080 31024 22092
rect 30791 22052 31024 22080
rect 30791 22049 30803 22052
rect 30745 22043 30803 22049
rect 31018 22040 31024 22052
rect 31076 22040 31082 22092
rect 32953 22083 33011 22089
rect 32953 22049 32965 22083
rect 32999 22080 33011 22083
rect 33226 22080 33232 22092
rect 32999 22052 33232 22080
rect 32999 22049 33011 22052
rect 32953 22043 33011 22049
rect 33226 22040 33232 22052
rect 33284 22040 33290 22092
rect 35894 22080 35900 22092
rect 35820 22052 35900 22080
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 29825 22015 29883 22021
rect 29825 21981 29837 22015
rect 29871 21981 29883 22015
rect 29825 21975 29883 21981
rect 30009 22015 30067 22021
rect 30009 21981 30021 22015
rect 30055 21981 30067 22015
rect 30009 21975 30067 21981
rect 30561 22015 30619 22021
rect 30561 21981 30573 22015
rect 30607 22012 30619 22015
rect 30650 22012 30656 22024
rect 30607 21984 30656 22012
rect 30607 21981 30619 21984
rect 30561 21975 30619 21981
rect 19426 21944 19432 21956
rect 18708 21916 19432 21944
rect 19426 21904 19432 21916
rect 19484 21904 19490 21956
rect 21821 21947 21879 21953
rect 21821 21913 21833 21947
rect 21867 21944 21879 21947
rect 22649 21947 22707 21953
rect 22649 21944 22661 21947
rect 21867 21916 22661 21944
rect 21867 21913 21879 21916
rect 21821 21907 21879 21913
rect 22649 21913 22661 21916
rect 22695 21944 22707 21947
rect 25216 21947 25274 21953
rect 22695 21916 23612 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 9766 21876 9772 21888
rect 5000 21848 9260 21876
rect 9727 21848 9772 21876
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 18322 21876 18328 21888
rect 18283 21848 18328 21876
rect 18322 21836 18328 21848
rect 18380 21836 18386 21888
rect 18782 21836 18788 21888
rect 18840 21876 18846 21888
rect 19245 21879 19303 21885
rect 19245 21876 19257 21879
rect 18840 21848 19257 21876
rect 18840 21836 18846 21848
rect 19245 21845 19257 21848
rect 19291 21845 19303 21879
rect 19245 21839 19303 21845
rect 19978 21836 19984 21888
rect 20036 21876 20042 21888
rect 20073 21879 20131 21885
rect 20073 21876 20085 21879
rect 20036 21848 20085 21876
rect 20036 21836 20042 21848
rect 20073 21845 20085 21848
rect 20119 21845 20131 21879
rect 20898 21876 20904 21888
rect 20859 21848 20904 21876
rect 20073 21839 20131 21845
rect 20898 21836 20904 21848
rect 20956 21836 20962 21888
rect 22557 21879 22615 21885
rect 22557 21845 22569 21879
rect 22603 21876 22615 21879
rect 23382 21876 23388 21888
rect 22603 21848 23388 21876
rect 22603 21845 22615 21848
rect 22557 21839 22615 21845
rect 23382 21836 23388 21848
rect 23440 21836 23446 21888
rect 23584 21885 23612 21916
rect 25216 21913 25228 21947
rect 25262 21944 25274 21947
rect 25498 21944 25504 21956
rect 25262 21916 25504 21944
rect 25262 21913 25274 21916
rect 25216 21907 25274 21913
rect 25498 21904 25504 21916
rect 25556 21904 25562 21956
rect 26694 21904 26700 21956
rect 26752 21944 26758 21956
rect 27341 21947 27399 21953
rect 27341 21944 27353 21947
rect 26752 21916 27353 21944
rect 26752 21904 26758 21916
rect 27341 21913 27353 21916
rect 27387 21944 27399 21947
rect 28258 21944 28264 21956
rect 27387 21916 28264 21944
rect 27387 21913 27399 21916
rect 27341 21907 27399 21913
rect 28258 21904 28264 21916
rect 28316 21904 28322 21956
rect 29178 21904 29184 21956
rect 29236 21944 29242 21956
rect 29840 21944 29868 21975
rect 30650 21972 30656 21984
rect 30708 22012 30714 22024
rect 31110 22012 31116 22024
rect 30708 21984 31116 22012
rect 30708 21972 30714 21984
rect 31110 21972 31116 21984
rect 31168 22012 31174 22024
rect 31205 22015 31263 22021
rect 31205 22012 31217 22015
rect 31168 21984 31217 22012
rect 31168 21972 31174 21984
rect 31205 21981 31217 21984
rect 31251 21981 31263 22015
rect 32769 22015 32827 22021
rect 32769 22012 32781 22015
rect 31205 21975 31263 21981
rect 31726 21984 32781 22012
rect 31726 21944 31754 21984
rect 32769 21981 32781 21984
rect 32815 22012 32827 22015
rect 34698 22012 34704 22024
rect 32815 21984 34704 22012
rect 32815 21981 32827 21984
rect 32769 21975 32827 21981
rect 34698 21972 34704 21984
rect 34756 21972 34762 22024
rect 35820 22021 35848 22052
rect 35894 22040 35900 22052
rect 35952 22040 35958 22092
rect 37734 22040 37740 22092
rect 37792 22080 37798 22092
rect 38197 22083 38255 22089
rect 38197 22080 38209 22083
rect 37792 22052 38209 22080
rect 37792 22040 37798 22052
rect 38197 22049 38209 22052
rect 38243 22080 38255 22083
rect 38243 22052 38976 22080
rect 38243 22049 38255 22052
rect 38197 22043 38255 22049
rect 35805 22015 35863 22021
rect 35805 21981 35817 22015
rect 35851 21981 35863 22015
rect 35805 21975 35863 21981
rect 36173 22015 36231 22021
rect 36173 21981 36185 22015
rect 36219 22012 36231 22015
rect 38838 22012 38844 22024
rect 36219 21984 38844 22012
rect 36219 21981 36231 21984
rect 36173 21975 36231 21981
rect 38838 21972 38844 21984
rect 38896 21972 38902 22024
rect 38948 22021 38976 22052
rect 39037 22021 39065 22120
rect 39114 22108 39120 22120
rect 39172 22108 39178 22160
rect 39960 22080 39988 22188
rect 41325 22185 41337 22188
rect 41371 22185 41383 22219
rect 41325 22179 41383 22185
rect 39224 22052 39988 22080
rect 38933 22015 38991 22021
rect 38933 21981 38945 22015
rect 38979 21981 38991 22015
rect 38933 21975 38991 21981
rect 39022 22015 39080 22021
rect 39022 21981 39034 22015
rect 39068 21981 39080 22015
rect 39022 21975 39080 21981
rect 39138 22015 39196 22021
rect 39138 21981 39150 22015
rect 39184 22012 39196 22015
rect 39224 22012 39252 22052
rect 39184 21984 39252 22012
rect 39301 22015 39359 22021
rect 39184 21981 39196 21984
rect 39138 21975 39196 21981
rect 39301 21981 39313 22015
rect 39347 22012 39359 22015
rect 39850 22012 39856 22024
rect 39347 21984 39856 22012
rect 39347 21981 39359 21984
rect 39301 21975 39359 21981
rect 39850 21972 39856 21984
rect 39908 21972 39914 22024
rect 40126 22012 40132 22024
rect 40087 21984 40132 22012
rect 40126 21972 40132 21984
rect 40184 21972 40190 22024
rect 40221 22015 40279 22021
rect 40221 21981 40233 22015
rect 40267 21981 40279 22015
rect 40221 21975 40279 21981
rect 32582 21944 32588 21956
rect 29236 21916 29868 21944
rect 30576 21916 31754 21944
rect 32543 21916 32588 21944
rect 29236 21904 29242 21916
rect 23569 21879 23627 21885
rect 23569 21845 23581 21879
rect 23615 21876 23627 21879
rect 23842 21876 23848 21888
rect 23615 21848 23848 21876
rect 23615 21845 23627 21848
rect 23569 21839 23627 21845
rect 23842 21836 23848 21848
rect 23900 21876 23906 21888
rect 26602 21876 26608 21888
rect 23900 21848 26608 21876
rect 23900 21836 23906 21848
rect 26602 21836 26608 21848
rect 26660 21876 26666 21888
rect 26789 21879 26847 21885
rect 26789 21876 26801 21879
rect 26660 21848 26801 21876
rect 26660 21836 26666 21848
rect 26789 21845 26801 21848
rect 26835 21845 26847 21879
rect 26789 21839 26847 21845
rect 28074 21836 28080 21888
rect 28132 21876 28138 21888
rect 30576 21876 30604 21916
rect 32582 21904 32588 21916
rect 32640 21904 32646 21956
rect 35897 21947 35955 21953
rect 35897 21913 35909 21947
rect 35943 21913 35955 21947
rect 35897 21907 35955 21913
rect 28132 21848 30604 21876
rect 28132 21836 28138 21848
rect 31938 21836 31944 21888
rect 31996 21876 32002 21888
rect 33318 21876 33324 21888
rect 31996 21848 33324 21876
rect 31996 21836 32002 21848
rect 33318 21836 33324 21848
rect 33376 21836 33382 21888
rect 33502 21876 33508 21888
rect 33463 21848 33508 21876
rect 33502 21836 33508 21848
rect 33560 21836 33566 21888
rect 35618 21876 35624 21888
rect 35579 21848 35624 21876
rect 35618 21836 35624 21848
rect 35676 21836 35682 21888
rect 35912 21876 35940 21907
rect 35986 21904 35992 21956
rect 36044 21944 36050 21956
rect 38746 21944 38752 21956
rect 36044 21916 36089 21944
rect 37016 21916 38752 21944
rect 36044 21904 36050 21916
rect 37016 21876 37044 21916
rect 38746 21904 38752 21916
rect 38804 21904 38810 21956
rect 40236 21944 40264 21975
rect 40310 21972 40316 22024
rect 40368 22012 40374 22024
rect 40368 21984 40413 22012
rect 40368 21972 40374 21984
rect 40494 21972 40500 22024
rect 40552 22012 40558 22024
rect 40552 21984 40597 22012
rect 40552 21972 40558 21984
rect 40678 21944 40684 21956
rect 40236 21916 40684 21944
rect 40678 21904 40684 21916
rect 40736 21904 40742 21956
rect 40954 21944 40960 21956
rect 40915 21916 40960 21944
rect 40954 21904 40960 21916
rect 41012 21904 41018 21956
rect 41138 21944 41144 21956
rect 41099 21916 41144 21944
rect 41138 21904 41144 21916
rect 41196 21904 41202 21956
rect 37182 21876 37188 21888
rect 35912 21848 37044 21876
rect 37143 21848 37188 21876
rect 37182 21836 37188 21848
rect 37240 21836 37246 21888
rect 38654 21876 38660 21888
rect 38615 21848 38660 21876
rect 38654 21836 38660 21848
rect 38712 21836 38718 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 3789 21675 3847 21681
rect 3789 21641 3801 21675
rect 3835 21672 3847 21675
rect 3878 21672 3884 21684
rect 3835 21644 3884 21672
rect 3835 21641 3847 21644
rect 3789 21635 3847 21641
rect 3878 21632 3884 21644
rect 3936 21632 3942 21684
rect 3970 21632 3976 21684
rect 4028 21672 4034 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 4028 21644 5641 21672
rect 4028 21632 4034 21644
rect 5629 21641 5641 21644
rect 5675 21672 5687 21675
rect 9398 21672 9404 21684
rect 5675 21644 9404 21672
rect 5675 21641 5687 21644
rect 5629 21635 5687 21641
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 14274 21672 14280 21684
rect 12728 21644 14280 21672
rect 4516 21607 4574 21613
rect 2424 21576 4292 21604
rect 2424 21545 2452 21576
rect 4264 21548 4292 21576
rect 4516 21573 4528 21607
rect 4562 21604 4574 21607
rect 4614 21604 4620 21616
rect 4562 21576 4620 21604
rect 4562 21573 4574 21576
rect 4516 21567 4574 21573
rect 4614 21564 4620 21576
rect 4672 21564 4678 21616
rect 6730 21604 6736 21616
rect 6691 21576 6736 21604
rect 6730 21564 6736 21576
rect 6788 21564 6794 21616
rect 7101 21607 7159 21613
rect 7101 21573 7113 21607
rect 7147 21604 7159 21607
rect 7926 21604 7932 21616
rect 7147 21576 7932 21604
rect 7147 21573 7159 21576
rect 7101 21567 7159 21573
rect 7926 21564 7932 21576
rect 7984 21564 7990 21616
rect 12158 21564 12164 21616
rect 12216 21604 12222 21616
rect 12728 21613 12756 21644
rect 14274 21632 14280 21644
rect 14332 21632 14338 21684
rect 14550 21672 14556 21684
rect 14511 21644 14556 21672
rect 14550 21632 14556 21644
rect 14608 21632 14614 21684
rect 18230 21672 18236 21684
rect 17328 21644 18236 21672
rect 12713 21607 12771 21613
rect 12713 21604 12725 21607
rect 12216 21576 12725 21604
rect 12216 21564 12222 21576
rect 12713 21573 12725 21576
rect 12759 21573 12771 21607
rect 12713 21567 12771 21573
rect 12802 21564 12808 21616
rect 12860 21604 12866 21616
rect 17328 21613 17356 21644
rect 18230 21632 18236 21644
rect 18288 21672 18294 21684
rect 21177 21675 21235 21681
rect 21177 21672 21189 21675
rect 18288 21644 21189 21672
rect 18288 21632 18294 21644
rect 21177 21641 21189 21644
rect 21223 21641 21235 21675
rect 21177 21635 21235 21641
rect 22066 21644 22876 21672
rect 12897 21607 12955 21613
rect 12897 21604 12909 21607
rect 12860 21576 12909 21604
rect 12860 21564 12866 21576
rect 12897 21573 12909 21576
rect 12943 21604 12955 21607
rect 17313 21607 17371 21613
rect 17313 21604 17325 21607
rect 12943 21576 17325 21604
rect 12943 21573 12955 21576
rect 12897 21567 12955 21573
rect 17313 21573 17325 21576
rect 17359 21573 17371 21607
rect 17313 21567 17371 21573
rect 17880 21576 20668 21604
rect 17880 21548 17908 21576
rect 2682 21545 2688 21548
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21505 2467 21539
rect 2676 21536 2688 21545
rect 2643 21508 2688 21536
rect 2409 21499 2467 21505
rect 2676 21499 2688 21508
rect 2682 21496 2688 21499
rect 2740 21496 2746 21548
rect 4246 21536 4252 21548
rect 4207 21508 4252 21536
rect 4246 21496 4252 21508
rect 4304 21496 4310 21548
rect 8196 21539 8254 21545
rect 8196 21505 8208 21539
rect 8242 21536 8254 21539
rect 10134 21536 10140 21548
rect 8242 21508 10140 21536
rect 8242 21505 8254 21508
rect 8196 21499 8254 21505
rect 10134 21496 10140 21508
rect 10192 21496 10198 21548
rect 13906 21536 13912 21548
rect 13867 21508 13912 21536
rect 13906 21496 13912 21508
rect 13964 21496 13970 21548
rect 14090 21536 14096 21548
rect 14051 21508 14096 21536
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14323 21539 14381 21545
rect 14240 21508 14285 21536
rect 14240 21496 14246 21508
rect 14323 21505 14335 21539
rect 14369 21536 14381 21539
rect 15194 21536 15200 21548
rect 14369 21505 14403 21536
rect 15155 21508 15200 21536
rect 14323 21499 14403 21505
rect 7742 21428 7748 21480
rect 7800 21468 7806 21480
rect 7929 21471 7987 21477
rect 7929 21468 7941 21471
rect 7800 21440 7941 21468
rect 7800 21428 7806 21440
rect 7929 21437 7941 21440
rect 7975 21437 7987 21471
rect 14375 21468 14403 21499
rect 15194 21496 15200 21508
rect 15252 21496 15258 21548
rect 15381 21539 15439 21545
rect 15381 21505 15393 21539
rect 15427 21536 15439 21539
rect 16025 21539 16083 21545
rect 16025 21536 16037 21539
rect 15427 21508 16037 21536
rect 15427 21505 15439 21508
rect 15381 21499 15439 21505
rect 16025 21505 16037 21508
rect 16071 21536 16083 21539
rect 16942 21536 16948 21548
rect 16071 21508 16948 21536
rect 16071 21505 16083 21508
rect 16025 21499 16083 21505
rect 16942 21496 16948 21508
rect 17000 21496 17006 21548
rect 17862 21536 17868 21548
rect 17775 21508 17868 21536
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 18026 21536 18032 21548
rect 17987 21508 18032 21536
rect 18026 21496 18032 21508
rect 18084 21496 18090 21548
rect 18141 21539 18199 21545
rect 18141 21505 18153 21539
rect 18187 21505 18199 21539
rect 18141 21499 18199 21505
rect 7929 21431 7987 21437
rect 13372 21440 14403 21468
rect 11606 21400 11612 21412
rect 11519 21372 11612 21400
rect 11606 21360 11612 21372
rect 11664 21400 11670 21412
rect 12802 21400 12808 21412
rect 11664 21372 12808 21400
rect 11664 21360 11670 21372
rect 12802 21360 12808 21372
rect 12860 21360 12866 21412
rect 13372 21344 13400 21440
rect 14918 21428 14924 21480
rect 14976 21468 14982 21480
rect 15013 21471 15071 21477
rect 15013 21468 15025 21471
rect 14976 21440 15025 21468
rect 14976 21428 14982 21440
rect 15013 21437 15025 21440
rect 15059 21468 15071 21471
rect 15059 21440 16804 21468
rect 15059 21437 15071 21440
rect 15013 21431 15071 21437
rect 9309 21335 9367 21341
rect 9309 21301 9321 21335
rect 9355 21332 9367 21335
rect 11330 21332 11336 21344
rect 9355 21304 11336 21332
rect 9355 21301 9367 21304
rect 9309 21295 9367 21301
rect 11330 21292 11336 21304
rect 11388 21292 11394 21344
rect 12158 21332 12164 21344
rect 12119 21304 12164 21332
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 13354 21332 13360 21344
rect 13315 21304 13360 21332
rect 13354 21292 13360 21304
rect 13412 21292 13418 21344
rect 15746 21292 15752 21344
rect 15804 21332 15810 21344
rect 16776 21341 16804 21440
rect 17770 21428 17776 21480
rect 17828 21468 17834 21480
rect 18156 21468 18184 21499
rect 18230 21496 18236 21548
rect 18288 21536 18294 21548
rect 18966 21536 18972 21548
rect 18288 21508 18333 21536
rect 18927 21508 18972 21536
rect 18288 21496 18294 21508
rect 18966 21496 18972 21508
rect 19024 21496 19030 21548
rect 19153 21539 19211 21545
rect 19153 21505 19165 21539
rect 19199 21536 19211 21539
rect 20530 21536 20536 21548
rect 19199 21508 20536 21536
rect 19199 21505 19211 21508
rect 19153 21499 19211 21505
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 17828 21440 18184 21468
rect 17828 21428 17834 21440
rect 18598 21428 18604 21480
rect 18656 21468 18662 21480
rect 19797 21471 19855 21477
rect 19797 21468 19809 21471
rect 18656 21440 19809 21468
rect 18656 21428 18662 21440
rect 19797 21437 19809 21440
rect 19843 21468 19855 21471
rect 19978 21468 19984 21480
rect 19843 21440 19984 21468
rect 19843 21437 19855 21440
rect 19797 21431 19855 21437
rect 19978 21428 19984 21440
rect 20036 21428 20042 21480
rect 20073 21471 20131 21477
rect 20073 21437 20085 21471
rect 20119 21468 20131 21471
rect 20640 21468 20668 21576
rect 21192 21536 21220 21635
rect 22066 21616 22094 21644
rect 21266 21564 21272 21616
rect 21324 21604 21330 21616
rect 22002 21604 22008 21616
rect 21324 21576 22008 21604
rect 21324 21564 21330 21576
rect 22002 21564 22008 21576
rect 22060 21576 22094 21616
rect 22060 21564 22066 21576
rect 22848 21545 22876 21644
rect 24854 21632 24860 21684
rect 24912 21632 24918 21684
rect 25498 21672 25504 21684
rect 25459 21644 25504 21672
rect 25498 21632 25504 21644
rect 25556 21632 25562 21684
rect 27338 21672 27344 21684
rect 27299 21644 27344 21672
rect 27338 21632 27344 21644
rect 27396 21632 27402 21684
rect 28994 21672 29000 21684
rect 28092 21644 29000 21672
rect 24872 21604 24900 21632
rect 25961 21607 26019 21613
rect 25961 21604 25973 21607
rect 24872 21576 25973 21604
rect 25961 21573 25973 21576
rect 26007 21573 26019 21607
rect 25961 21567 26019 21573
rect 26050 21564 26056 21616
rect 26108 21604 26114 21616
rect 28092 21613 28120 21644
rect 28994 21632 29000 21644
rect 29052 21632 29058 21684
rect 29362 21672 29368 21684
rect 29323 21644 29368 21672
rect 29362 21632 29368 21644
rect 29420 21632 29426 21684
rect 31938 21672 31944 21684
rect 29748 21644 31944 21672
rect 26329 21607 26387 21613
rect 26329 21604 26341 21607
rect 26108 21576 26341 21604
rect 26108 21564 26114 21576
rect 26329 21573 26341 21576
rect 26375 21573 26387 21607
rect 26329 21567 26387 21573
rect 28077 21607 28135 21613
rect 28077 21573 28089 21607
rect 28123 21573 28135 21607
rect 28077 21567 28135 21573
rect 28169 21607 28227 21613
rect 28169 21573 28181 21607
rect 28215 21604 28227 21607
rect 29748 21604 29776 21644
rect 31938 21632 31944 21644
rect 31996 21632 32002 21684
rect 32122 21672 32128 21684
rect 32083 21644 32128 21672
rect 32122 21632 32128 21644
rect 32180 21632 32186 21684
rect 33502 21632 33508 21684
rect 33560 21672 33566 21684
rect 36446 21672 36452 21684
rect 33560 21644 36452 21672
rect 33560 21632 33566 21644
rect 36446 21632 36452 21644
rect 36504 21632 36510 21684
rect 39114 21672 39120 21684
rect 37660 21644 39120 21672
rect 28215 21576 29776 21604
rect 29825 21607 29883 21613
rect 28215 21573 28227 21576
rect 28169 21567 28227 21573
rect 29825 21573 29837 21607
rect 29871 21604 29883 21607
rect 30190 21604 30196 21616
rect 29871 21576 30196 21604
rect 29871 21573 29883 21576
rect 29825 21567 29883 21573
rect 30190 21564 30196 21576
rect 30248 21564 30254 21616
rect 30282 21564 30288 21616
rect 30340 21604 30346 21616
rect 30837 21607 30895 21613
rect 30837 21604 30849 21607
rect 30340 21576 30849 21604
rect 30340 21564 30346 21576
rect 30837 21573 30849 21576
rect 30883 21573 30895 21607
rect 30837 21567 30895 21573
rect 30929 21607 30987 21613
rect 30929 21573 30941 21607
rect 30975 21604 30987 21607
rect 32030 21604 32036 21616
rect 30975 21576 32036 21604
rect 30975 21573 30987 21576
rect 30929 21567 30987 21573
rect 32030 21564 32036 21576
rect 32088 21564 32094 21616
rect 32214 21564 32220 21616
rect 32272 21604 32278 21616
rect 32585 21607 32643 21613
rect 32585 21604 32597 21607
rect 32272 21576 32597 21604
rect 32272 21564 32278 21576
rect 32585 21573 32597 21576
rect 32631 21573 32643 21607
rect 32585 21567 32643 21573
rect 35612 21607 35670 21613
rect 35612 21573 35624 21607
rect 35658 21604 35670 21607
rect 37277 21607 37335 21613
rect 37277 21604 37289 21607
rect 35658 21576 37289 21604
rect 35658 21573 35670 21576
rect 35612 21567 35670 21573
rect 37277 21573 37289 21576
rect 37323 21573 37335 21607
rect 37277 21567 37335 21573
rect 22465 21539 22523 21545
rect 22465 21536 22477 21539
rect 21192 21508 22477 21536
rect 22465 21505 22477 21508
rect 22511 21505 22523 21539
rect 22465 21499 22523 21505
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 22649 21539 22707 21545
rect 22649 21505 22661 21539
rect 22695 21505 22707 21539
rect 22649 21499 22707 21505
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21536 22891 21539
rect 24857 21539 24915 21545
rect 24857 21536 24869 21539
rect 22879 21508 24869 21536
rect 22879 21505 22891 21508
rect 22833 21499 22891 21505
rect 24857 21505 24869 21508
rect 24903 21505 24915 21539
rect 25038 21536 25044 21548
rect 24999 21508 25044 21536
rect 24857 21499 24915 21505
rect 20806 21468 20812 21480
rect 20119 21440 20812 21468
rect 20119 21437 20131 21440
rect 20073 21431 20131 21437
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 21726 21428 21732 21480
rect 21784 21468 21790 21480
rect 22572 21468 22600 21499
rect 21784 21440 22600 21468
rect 22664 21468 22692 21499
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 25133 21539 25191 21545
rect 25133 21505 25145 21539
rect 25179 21505 25191 21539
rect 25133 21499 25191 21505
rect 23474 21468 23480 21480
rect 22664 21440 23480 21468
rect 21784 21428 21790 21440
rect 18230 21360 18236 21412
rect 18288 21400 18294 21412
rect 19337 21403 19395 21409
rect 19337 21400 19349 21403
rect 18288 21372 19349 21400
rect 18288 21360 18294 21372
rect 19337 21369 19349 21372
rect 19383 21369 19395 21403
rect 22572 21400 22600 21440
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21437 23627 21471
rect 23569 21431 23627 21437
rect 23845 21471 23903 21477
rect 23845 21437 23857 21471
rect 23891 21468 23903 21471
rect 24946 21468 24952 21480
rect 23891 21440 24952 21468
rect 23891 21437 23903 21440
rect 23845 21431 23903 21437
rect 23584 21400 23612 21431
rect 24946 21428 24952 21440
rect 25004 21468 25010 21480
rect 25148 21468 25176 21499
rect 25222 21496 25228 21548
rect 25280 21536 25286 21548
rect 25280 21508 25325 21536
rect 25280 21496 25286 21508
rect 25590 21496 25596 21548
rect 25648 21536 25654 21548
rect 26068 21536 26096 21564
rect 25648 21508 26096 21536
rect 26145 21539 26203 21545
rect 25648 21496 25654 21508
rect 26145 21505 26157 21539
rect 26191 21505 26203 21539
rect 26145 21499 26203 21505
rect 25004 21440 25176 21468
rect 26160 21468 26188 21499
rect 26602 21496 26608 21548
rect 26660 21536 26666 21548
rect 27249 21539 27307 21545
rect 27249 21536 27261 21539
rect 26660 21508 27261 21536
rect 26660 21496 26666 21508
rect 27249 21505 27261 21508
rect 27295 21505 27307 21539
rect 27249 21499 27307 21505
rect 27430 21496 27436 21548
rect 27488 21536 27494 21548
rect 27893 21539 27951 21545
rect 27893 21536 27905 21539
rect 27488 21508 27905 21536
rect 27488 21496 27494 21508
rect 27893 21505 27905 21508
rect 27939 21505 27951 21539
rect 27893 21499 27951 21505
rect 28261 21539 28319 21545
rect 28261 21505 28273 21539
rect 28307 21505 28319 21539
rect 28261 21499 28319 21505
rect 29549 21539 29607 21545
rect 29549 21505 29561 21539
rect 29595 21505 29607 21539
rect 29549 21499 29607 21505
rect 26970 21468 26976 21480
rect 26160 21440 26976 21468
rect 25004 21428 25010 21440
rect 26970 21428 26976 21440
rect 27028 21428 27034 21480
rect 28166 21428 28172 21480
rect 28224 21468 28230 21480
rect 28276 21468 28304 21499
rect 28224 21440 28304 21468
rect 28224 21428 28230 21440
rect 22572 21372 23612 21400
rect 19337 21363 19395 21369
rect 25774 21360 25780 21412
rect 25832 21400 25838 21412
rect 28534 21400 28540 21412
rect 25832 21372 28540 21400
rect 25832 21360 25838 21372
rect 28534 21360 28540 21372
rect 28592 21360 28598 21412
rect 29564 21400 29592 21499
rect 29730 21496 29736 21548
rect 29788 21536 29794 21548
rect 30653 21539 30711 21545
rect 30653 21536 30665 21539
rect 29788 21508 30665 21536
rect 29788 21496 29794 21508
rect 30653 21505 30665 21508
rect 30699 21505 30711 21539
rect 30653 21499 30711 21505
rect 31021 21539 31079 21545
rect 31021 21505 31033 21539
rect 31067 21536 31079 21539
rect 31110 21536 31116 21548
rect 31067 21508 31116 21536
rect 31067 21505 31079 21508
rect 31021 21499 31079 21505
rect 31110 21496 31116 21508
rect 31168 21496 31174 21548
rect 32306 21536 32312 21548
rect 32267 21508 32312 21536
rect 32306 21496 32312 21508
rect 32364 21496 32370 21548
rect 37182 21496 37188 21548
rect 37240 21536 37246 21548
rect 37660 21545 37688 21644
rect 39114 21632 39120 21644
rect 39172 21672 39178 21684
rect 40678 21672 40684 21684
rect 39172 21644 40684 21672
rect 39172 21632 39178 21644
rect 40678 21632 40684 21644
rect 40736 21632 40742 21684
rect 38654 21564 38660 21616
rect 38712 21604 38718 21616
rect 38994 21607 39052 21613
rect 38994 21604 39006 21607
rect 38712 21576 39006 21604
rect 38712 21564 38718 21576
rect 38994 21573 39006 21576
rect 39040 21573 39052 21607
rect 38994 21567 39052 21573
rect 39758 21564 39764 21616
rect 39816 21604 39822 21616
rect 40954 21604 40960 21616
rect 39816 21576 40960 21604
rect 39816 21564 39822 21576
rect 40954 21564 40960 21576
rect 41012 21564 41018 21616
rect 37553 21539 37611 21545
rect 37553 21536 37565 21539
rect 37240 21508 37565 21536
rect 37240 21496 37246 21508
rect 37553 21505 37565 21508
rect 37599 21505 37611 21539
rect 37553 21499 37611 21505
rect 37645 21539 37703 21545
rect 37645 21505 37657 21539
rect 37691 21505 37703 21539
rect 37645 21499 37703 21505
rect 37734 21496 37740 21548
rect 37792 21536 37798 21548
rect 37921 21539 37979 21545
rect 37792 21508 37837 21536
rect 37792 21496 37798 21508
rect 37921 21505 37933 21539
rect 37967 21505 37979 21539
rect 37921 21499 37979 21505
rect 29641 21471 29699 21477
rect 29641 21437 29653 21471
rect 29687 21468 29699 21471
rect 30006 21468 30012 21480
rect 29687 21440 30012 21468
rect 29687 21437 29699 21440
rect 29641 21431 29699 21437
rect 30006 21428 30012 21440
rect 30064 21428 30070 21480
rect 32030 21428 32036 21480
rect 32088 21468 32094 21480
rect 32401 21471 32459 21477
rect 32401 21468 32413 21471
rect 32088 21440 32413 21468
rect 32088 21428 32094 21440
rect 32401 21437 32413 21440
rect 32447 21437 32459 21471
rect 35342 21468 35348 21480
rect 35303 21440 35348 21468
rect 32401 21431 32459 21437
rect 35342 21428 35348 21440
rect 35400 21428 35406 21480
rect 36538 21428 36544 21480
rect 36596 21468 36602 21480
rect 37936 21468 37964 21499
rect 40034 21496 40040 21548
rect 40092 21536 40098 21548
rect 40402 21536 40408 21548
rect 40092 21508 40408 21536
rect 40092 21496 40098 21508
rect 40402 21496 40408 21508
rect 40460 21536 40466 21548
rect 40586 21536 40592 21548
rect 40460 21508 40592 21536
rect 40460 21496 40466 21508
rect 40586 21496 40592 21508
rect 40644 21496 40650 21548
rect 36596 21440 37964 21468
rect 38749 21471 38807 21477
rect 36596 21428 36602 21440
rect 38749 21437 38761 21471
rect 38795 21437 38807 21471
rect 38749 21431 38807 21437
rect 31205 21403 31263 21409
rect 29564 21372 30696 21400
rect 15841 21335 15899 21341
rect 15841 21332 15853 21335
rect 15804 21304 15853 21332
rect 15804 21292 15810 21304
rect 15841 21301 15853 21304
rect 15887 21301 15899 21335
rect 15841 21295 15899 21301
rect 16761 21335 16819 21341
rect 16761 21301 16773 21335
rect 16807 21332 16819 21335
rect 17954 21332 17960 21344
rect 16807 21304 17960 21332
rect 16807 21301 16819 21304
rect 16761 21295 16819 21301
rect 17954 21292 17960 21304
rect 18012 21292 18018 21344
rect 18506 21332 18512 21344
rect 18467 21304 18512 21332
rect 18506 21292 18512 21304
rect 18564 21292 18570 21344
rect 22189 21335 22247 21341
rect 22189 21301 22201 21335
rect 22235 21332 22247 21335
rect 22462 21332 22468 21344
rect 22235 21304 22468 21332
rect 22235 21301 22247 21304
rect 22189 21295 22247 21301
rect 22462 21292 22468 21304
rect 22520 21292 22526 21344
rect 28445 21335 28503 21341
rect 28445 21301 28457 21335
rect 28491 21332 28503 21335
rect 29549 21335 29607 21341
rect 29549 21332 29561 21335
rect 28491 21304 29561 21332
rect 28491 21301 28503 21304
rect 28445 21295 28503 21301
rect 29549 21301 29561 21304
rect 29595 21301 29607 21335
rect 30668 21332 30696 21372
rect 31205 21369 31217 21403
rect 31251 21400 31263 21403
rect 31251 21372 32444 21400
rect 31251 21369 31263 21372
rect 31205 21363 31263 21369
rect 32214 21332 32220 21344
rect 30668 21304 32220 21332
rect 29549 21295 29607 21301
rect 32214 21292 32220 21304
rect 32272 21292 32278 21344
rect 32416 21341 32444 21372
rect 32401 21335 32459 21341
rect 32401 21301 32413 21335
rect 32447 21301 32459 21335
rect 32401 21295 32459 21301
rect 36725 21335 36783 21341
rect 36725 21301 36737 21335
rect 36771 21332 36783 21335
rect 36906 21332 36912 21344
rect 36771 21304 36912 21332
rect 36771 21301 36783 21304
rect 36725 21295 36783 21301
rect 36906 21292 36912 21304
rect 36964 21292 36970 21344
rect 38764 21332 38792 21431
rect 40034 21332 40040 21344
rect 38764 21304 40040 21332
rect 40034 21292 40040 21304
rect 40092 21292 40098 21344
rect 40126 21292 40132 21344
rect 40184 21332 40190 21344
rect 41138 21332 41144 21344
rect 40184 21304 41144 21332
rect 40184 21292 40190 21304
rect 41138 21292 41144 21304
rect 41196 21292 41202 21344
rect 58158 21332 58164 21344
rect 58119 21304 58164 21332
rect 58158 21292 58164 21304
rect 58216 21292 58222 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 10134 21128 10140 21140
rect 10095 21100 10140 21128
rect 10134 21088 10140 21100
rect 10192 21088 10198 21140
rect 11790 21128 11796 21140
rect 10244 21100 11796 21128
rect 1854 21020 1860 21072
rect 1912 21060 1918 21072
rect 10244 21060 10272 21100
rect 11790 21088 11796 21100
rect 11848 21088 11854 21140
rect 14090 21088 14096 21140
rect 14148 21128 14154 21140
rect 15381 21131 15439 21137
rect 15381 21128 15393 21131
rect 14148 21100 15393 21128
rect 14148 21088 14154 21100
rect 15381 21097 15393 21100
rect 15427 21097 15439 21131
rect 15381 21091 15439 21097
rect 17589 21131 17647 21137
rect 17589 21097 17601 21131
rect 17635 21128 17647 21131
rect 18046 21128 18052 21140
rect 17635 21100 18052 21128
rect 17635 21097 17647 21100
rect 17589 21091 17647 21097
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 18138 21088 18144 21140
rect 18196 21128 18202 21140
rect 25130 21128 25136 21140
rect 18196 21100 19288 21128
rect 25091 21100 25136 21128
rect 18196 21088 18202 21100
rect 1912 21032 10272 21060
rect 1912 21020 1918 21032
rect 10502 21020 10508 21072
rect 10560 21060 10566 21072
rect 10560 21032 13216 21060
rect 10560 21020 10566 21032
rect 13188 21004 13216 21032
rect 16942 21020 16948 21072
rect 17000 21060 17006 21072
rect 18966 21060 18972 21072
rect 17000 21032 18972 21060
rect 17000 21020 17006 21032
rect 18966 21020 18972 21032
rect 19024 21020 19030 21072
rect 10226 20952 10232 21004
rect 10284 20992 10290 21004
rect 11241 20995 11299 21001
rect 11241 20992 11253 20995
rect 10284 20964 11253 20992
rect 10284 20952 10290 20964
rect 10796 20936 10824 20964
rect 11241 20961 11253 20964
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 13170 20952 13176 21004
rect 13228 20992 13234 21004
rect 14182 20992 14188 21004
rect 13228 20964 14188 20992
rect 13228 20952 13234 20964
rect 14182 20952 14188 20964
rect 14240 20992 14246 21004
rect 14369 20995 14427 21001
rect 14369 20992 14381 20995
rect 14240 20964 14381 20992
rect 14240 20952 14246 20964
rect 14369 20961 14381 20964
rect 14415 20961 14427 20995
rect 17770 20992 17776 21004
rect 14369 20955 14427 20961
rect 15495 20964 16436 20992
rect 9674 20924 9680 20936
rect 9635 20896 9680 20924
rect 9674 20884 9680 20896
rect 9732 20924 9738 20936
rect 10367 20927 10425 20933
rect 10367 20924 10379 20927
rect 9732 20896 10379 20924
rect 9732 20884 9738 20896
rect 10367 20893 10379 20896
rect 10413 20893 10425 20927
rect 10502 20924 10508 20936
rect 10463 20896 10508 20924
rect 10367 20887 10425 20893
rect 10502 20884 10508 20896
rect 10560 20884 10566 20936
rect 10597 20927 10655 20933
rect 10597 20893 10609 20927
rect 10643 20893 10655 20927
rect 10597 20887 10655 20893
rect 5721 20859 5779 20865
rect 5721 20825 5733 20859
rect 5767 20856 5779 20859
rect 6914 20856 6920 20868
rect 5767 20828 6920 20856
rect 5767 20825 5779 20828
rect 5721 20819 5779 20825
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 7469 20859 7527 20865
rect 7469 20825 7481 20859
rect 7515 20856 7527 20859
rect 7742 20856 7748 20868
rect 7515 20828 7748 20856
rect 7515 20825 7527 20828
rect 7469 20819 7527 20825
rect 7742 20816 7748 20828
rect 7800 20816 7806 20868
rect 10612 20856 10640 20887
rect 10778 20884 10784 20936
rect 10836 20924 10842 20936
rect 11425 20927 11483 20933
rect 10836 20896 10929 20924
rect 10836 20884 10842 20896
rect 11425 20893 11437 20927
rect 11471 20924 11483 20927
rect 11606 20924 11612 20936
rect 11471 20896 11612 20924
rect 11471 20893 11483 20896
rect 11425 20887 11483 20893
rect 11606 20884 11612 20896
rect 11664 20884 11670 20936
rect 14090 20924 14096 20936
rect 14051 20896 14096 20924
rect 14090 20884 14096 20896
rect 14148 20924 14154 20936
rect 15495 20924 15523 20964
rect 14148 20896 15523 20924
rect 15565 20927 15623 20933
rect 14148 20884 14154 20896
rect 15565 20893 15577 20927
rect 15611 20924 15623 20927
rect 15654 20924 15660 20936
rect 15611 20896 15660 20924
rect 15611 20893 15623 20896
rect 15565 20887 15623 20893
rect 15654 20884 15660 20896
rect 15712 20884 15718 20936
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 16408 20924 16436 20964
rect 17236 20964 17776 20992
rect 15804 20896 15849 20924
rect 16408 20921 17172 20924
rect 17236 20921 17264 20964
rect 17770 20952 17776 20964
rect 17828 20992 17834 21004
rect 19260 21001 19288 21100
rect 25130 21088 25136 21100
rect 25188 21088 25194 21140
rect 28350 21128 28356 21140
rect 28311 21100 28356 21128
rect 28350 21088 28356 21100
rect 28408 21088 28414 21140
rect 28534 21088 28540 21140
rect 28592 21128 28598 21140
rect 30190 21128 30196 21140
rect 28592 21100 30196 21128
rect 28592 21088 28598 21100
rect 30190 21088 30196 21100
rect 30248 21088 30254 21140
rect 31297 21131 31355 21137
rect 31297 21097 31309 21131
rect 31343 21128 31355 21131
rect 32125 21131 32183 21137
rect 32125 21128 32137 21131
rect 31343 21100 32137 21128
rect 31343 21097 31355 21100
rect 31297 21091 31355 21097
rect 32125 21097 32137 21100
rect 32171 21097 32183 21131
rect 32125 21091 32183 21097
rect 32306 21088 32312 21140
rect 32364 21128 32370 21140
rect 35621 21131 35679 21137
rect 35621 21128 35633 21131
rect 32364 21100 35633 21128
rect 32364 21088 32370 21100
rect 35621 21097 35633 21100
rect 35667 21097 35679 21131
rect 35621 21091 35679 21097
rect 36725 21131 36783 21137
rect 36725 21097 36737 21131
rect 36771 21128 36783 21131
rect 37734 21128 37740 21140
rect 36771 21100 37740 21128
rect 36771 21097 36783 21100
rect 36725 21091 36783 21097
rect 37734 21088 37740 21100
rect 37792 21088 37798 21140
rect 40221 21131 40279 21137
rect 40221 21097 40233 21131
rect 40267 21128 40279 21131
rect 40494 21128 40500 21140
rect 40267 21100 40500 21128
rect 40267 21097 40279 21100
rect 40221 21091 40279 21097
rect 40494 21088 40500 21100
rect 40552 21088 40558 21140
rect 22278 21060 22284 21072
rect 21468 21032 22284 21060
rect 19245 20995 19303 21001
rect 17828 20964 18368 20992
rect 17828 20952 17834 20964
rect 16408 20896 17264 20921
rect 15804 20884 15810 20896
rect 17144 20893 17264 20896
rect 17328 20896 17816 20924
rect 11146 20856 11152 20868
rect 10612 20828 11152 20856
rect 11146 20816 11152 20828
rect 11204 20816 11210 20868
rect 12253 20859 12311 20865
rect 12253 20825 12265 20859
rect 12299 20856 12311 20859
rect 12805 20859 12863 20865
rect 12805 20856 12817 20859
rect 12299 20828 12817 20856
rect 12299 20825 12311 20828
rect 12253 20819 12311 20825
rect 12805 20825 12817 20828
rect 12851 20856 12863 20859
rect 15286 20856 15292 20868
rect 12851 20828 15292 20856
rect 12851 20825 12863 20828
rect 12805 20819 12863 20825
rect 15286 20816 15292 20828
rect 15344 20816 15350 20868
rect 16942 20816 16948 20868
rect 17000 20856 17006 20868
rect 17221 20859 17279 20865
rect 17221 20856 17233 20859
rect 17000 20828 17233 20856
rect 17000 20816 17006 20828
rect 17221 20825 17233 20828
rect 17267 20825 17279 20859
rect 17221 20819 17279 20825
rect 17328 20800 17356 20896
rect 17405 20859 17463 20865
rect 17405 20825 17417 20859
rect 17451 20825 17463 20859
rect 17788 20856 17816 20896
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 18049 20927 18107 20933
rect 18049 20924 18061 20927
rect 17920 20896 18061 20924
rect 17920 20884 17926 20896
rect 18049 20893 18061 20896
rect 18095 20893 18107 20927
rect 18230 20924 18236 20936
rect 18191 20896 18236 20924
rect 18049 20887 18107 20893
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 18340 20933 18368 20964
rect 19245 20961 19257 20995
rect 19291 20961 19303 20995
rect 19245 20955 19303 20961
rect 18325 20927 18383 20933
rect 18325 20893 18337 20927
rect 18371 20893 18383 20927
rect 18325 20887 18383 20893
rect 18417 20927 18475 20933
rect 18417 20893 18429 20927
rect 18463 20924 18475 20927
rect 21082 20924 21088 20936
rect 18463 20896 21088 20924
rect 18463 20893 18475 20896
rect 18417 20887 18475 20893
rect 18432 20856 18460 20887
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 21266 20924 21272 20936
rect 21227 20896 21272 20924
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 21468 20933 21496 21032
rect 22278 21020 22284 21032
rect 22336 21020 22342 21072
rect 24581 21063 24639 21069
rect 24581 21029 24593 21063
rect 24627 21060 24639 21063
rect 25590 21060 25596 21072
rect 24627 21032 25596 21060
rect 24627 21029 24639 21032
rect 24581 21023 24639 21029
rect 25590 21020 25596 21032
rect 25648 21020 25654 21072
rect 26970 21060 26976 21072
rect 26883 21032 26976 21060
rect 26970 21020 26976 21032
rect 27028 21060 27034 21072
rect 27028 21032 29776 21060
rect 27028 21020 27034 21032
rect 21726 20992 21732 21004
rect 21560 20964 21732 20992
rect 21560 20933 21588 20964
rect 21726 20952 21732 20964
rect 21784 20952 21790 21004
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 21545 20927 21603 20933
rect 21545 20893 21557 20927
rect 21591 20893 21603 20927
rect 21545 20887 21603 20893
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 17788 20828 18460 20856
rect 18693 20859 18751 20865
rect 17405 20819 17463 20825
rect 18693 20825 18705 20859
rect 18739 20856 18751 20859
rect 19490 20859 19548 20865
rect 19490 20856 19502 20859
rect 18739 20828 19502 20856
rect 18739 20825 18751 20828
rect 18693 20819 18751 20825
rect 19490 20825 19502 20828
rect 19536 20825 19548 20859
rect 21100 20856 21128 20884
rect 21652 20856 21680 20887
rect 22094 20884 22100 20936
rect 22152 20924 22158 20936
rect 22373 20927 22431 20933
rect 22373 20924 22385 20927
rect 22152 20896 22385 20924
rect 22152 20884 22158 20896
rect 22373 20893 22385 20896
rect 22419 20893 22431 20927
rect 22373 20887 22431 20893
rect 22462 20884 22468 20936
rect 22520 20924 22526 20936
rect 22629 20927 22687 20933
rect 22629 20924 22641 20927
rect 22520 20896 22641 20924
rect 22520 20884 22526 20896
rect 22629 20893 22641 20896
rect 22675 20893 22687 20927
rect 22629 20887 22687 20893
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 24176 20896 24409 20924
rect 24176 20884 24182 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 25593 20927 25651 20933
rect 25593 20893 25605 20927
rect 25639 20924 25651 20927
rect 26234 20924 26240 20936
rect 25639 20896 26240 20924
rect 25639 20893 25651 20896
rect 25593 20887 25651 20893
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 27062 20884 27068 20936
rect 27120 20924 27126 20936
rect 27801 20927 27859 20933
rect 27801 20924 27813 20927
rect 27120 20896 27813 20924
rect 27120 20884 27126 20896
rect 27801 20893 27813 20896
rect 27847 20893 27859 20927
rect 28074 20924 28080 20936
rect 28035 20896 28080 20924
rect 27801 20887 27859 20893
rect 28074 20884 28080 20896
rect 28132 20884 28138 20936
rect 28166 20884 28172 20936
rect 28224 20924 28230 20936
rect 29748 20933 29776 21032
rect 30098 21020 30104 21072
rect 30156 21060 30162 21072
rect 31110 21060 31116 21072
rect 30156 21032 31116 21060
rect 30156 21020 30162 21032
rect 31110 21020 31116 21032
rect 31168 21020 31174 21072
rect 31938 21060 31944 21072
rect 31899 21032 31944 21060
rect 31938 21020 31944 21032
rect 31996 21020 32002 21072
rect 32214 21020 32220 21072
rect 32272 21060 32278 21072
rect 34790 21060 34796 21072
rect 32272 21032 34796 21060
rect 32272 21020 32278 21032
rect 34790 21020 34796 21032
rect 34848 21020 34854 21072
rect 35894 21060 35900 21072
rect 35820 21032 35900 21060
rect 30282 20992 30288 21004
rect 29932 20964 30288 20992
rect 29733 20927 29791 20933
rect 28224 20896 28269 20924
rect 28224 20884 28230 20896
rect 29733 20893 29745 20927
rect 29779 20893 29791 20927
rect 29733 20887 29791 20893
rect 25866 20865 25872 20868
rect 21100 20828 21680 20856
rect 25838 20859 25872 20865
rect 19490 20819 19548 20825
rect 25838 20825 25850 20859
rect 25838 20819 25872 20825
rect 7926 20788 7932 20800
rect 7887 20760 7932 20788
rect 7926 20748 7932 20760
rect 7984 20748 7990 20800
rect 10410 20748 10416 20800
rect 10468 20788 10474 20800
rect 12897 20791 12955 20797
rect 12897 20788 12909 20791
rect 10468 20760 12909 20788
rect 10468 20748 10474 20760
rect 12897 20757 12909 20760
rect 12943 20788 12955 20791
rect 17310 20788 17316 20800
rect 12943 20760 17316 20788
rect 12943 20757 12955 20760
rect 12897 20751 12955 20757
rect 17310 20748 17316 20760
rect 17368 20748 17374 20800
rect 17420 20788 17448 20819
rect 25866 20816 25872 20819
rect 25924 20816 25930 20868
rect 27985 20859 28043 20865
rect 27985 20825 27997 20859
rect 28031 20856 28043 20859
rect 28994 20856 29000 20868
rect 28031 20828 29000 20856
rect 28031 20825 28043 20828
rect 27985 20819 28043 20825
rect 28994 20816 29000 20828
rect 29052 20816 29058 20868
rect 29932 20865 29960 20964
rect 30282 20952 30288 20964
rect 30340 20992 30346 21004
rect 35618 20992 35624 21004
rect 30340 20964 30972 20992
rect 30340 20952 30346 20964
rect 30098 20924 30104 20936
rect 30059 20896 30104 20924
rect 30098 20884 30104 20896
rect 30156 20884 30162 20936
rect 30190 20884 30196 20936
rect 30248 20924 30254 20936
rect 30944 20933 30972 20964
rect 32140 20964 35624 20992
rect 30745 20927 30803 20933
rect 30745 20924 30757 20927
rect 30248 20896 30757 20924
rect 30248 20884 30254 20896
rect 30745 20893 30757 20896
rect 30791 20893 30803 20927
rect 30745 20887 30803 20893
rect 30929 20927 30987 20933
rect 30929 20893 30941 20927
rect 30975 20893 30987 20927
rect 31110 20924 31116 20936
rect 31071 20896 31116 20924
rect 30929 20887 30987 20893
rect 31110 20884 31116 20896
rect 31168 20884 31174 20936
rect 32140 20933 32168 20964
rect 35618 20952 35624 20964
rect 35676 20952 35682 21004
rect 32125 20927 32183 20933
rect 32125 20893 32137 20927
rect 32171 20893 32183 20927
rect 32125 20887 32183 20893
rect 32214 20884 32220 20936
rect 32272 20924 32278 20936
rect 35820 20933 35848 21032
rect 35894 21020 35900 21032
rect 35952 21020 35958 21072
rect 40126 20992 40132 21004
rect 35912 20964 40132 20992
rect 35912 20933 35940 20964
rect 40126 20952 40132 20964
rect 40184 20952 40190 21004
rect 35805 20927 35863 20933
rect 32272 20896 32317 20924
rect 32272 20884 32278 20896
rect 35805 20893 35817 20927
rect 35851 20893 35863 20927
rect 35805 20887 35863 20893
rect 35897 20927 35955 20933
rect 35897 20893 35909 20927
rect 35943 20893 35955 20927
rect 35897 20887 35955 20893
rect 35986 20884 35992 20936
rect 36044 20924 36050 20936
rect 36173 20927 36231 20933
rect 36044 20896 36089 20924
rect 36044 20884 36050 20896
rect 36173 20893 36185 20927
rect 36219 20924 36231 20927
rect 38930 20924 38936 20936
rect 36219 20896 38936 20924
rect 36219 20893 36231 20896
rect 36173 20887 36231 20893
rect 38930 20884 38936 20896
rect 38988 20884 38994 20936
rect 40037 20927 40095 20933
rect 40037 20893 40049 20927
rect 40083 20924 40095 20927
rect 40218 20924 40224 20936
rect 40083 20896 40224 20924
rect 40083 20893 40095 20896
rect 40037 20887 40095 20893
rect 40218 20884 40224 20896
rect 40276 20884 40282 20936
rect 29917 20859 29975 20865
rect 29917 20856 29929 20859
rect 29748 20828 29929 20856
rect 29748 20800 29776 20828
rect 29917 20825 29929 20828
rect 29963 20825 29975 20859
rect 29917 20819 29975 20825
rect 30009 20859 30067 20865
rect 30009 20825 30021 20859
rect 30055 20856 30067 20859
rect 30834 20856 30840 20868
rect 30055 20828 30840 20856
rect 30055 20825 30067 20828
rect 30009 20819 30067 20825
rect 30834 20816 30840 20828
rect 30892 20816 30898 20868
rect 31021 20859 31079 20865
rect 31021 20825 31033 20859
rect 31067 20856 31079 20859
rect 31754 20856 31760 20868
rect 31067 20828 31760 20856
rect 31067 20825 31079 20828
rect 31021 20819 31079 20825
rect 31754 20816 31760 20828
rect 31812 20816 31818 20868
rect 31846 20816 31852 20868
rect 31904 20856 31910 20868
rect 32401 20859 32459 20865
rect 32401 20856 32413 20859
rect 31904 20828 32413 20856
rect 31904 20816 31910 20828
rect 32401 20825 32413 20828
rect 32447 20825 32459 20859
rect 36906 20856 36912 20868
rect 36867 20828 36912 20856
rect 32401 20819 32459 20825
rect 36906 20816 36912 20828
rect 36964 20816 36970 20868
rect 37093 20859 37151 20865
rect 37093 20825 37105 20859
rect 37139 20856 37151 20859
rect 39758 20856 39764 20868
rect 37139 20828 39764 20856
rect 37139 20825 37151 20828
rect 37093 20819 37151 20825
rect 39758 20816 39764 20828
rect 39816 20856 39822 20868
rect 39853 20859 39911 20865
rect 39853 20856 39865 20859
rect 39816 20828 39865 20856
rect 39816 20816 39822 20828
rect 39853 20825 39865 20828
rect 39899 20825 39911 20859
rect 39853 20819 39911 20825
rect 19334 20788 19340 20800
rect 17420 20760 19340 20788
rect 19334 20748 19340 20760
rect 19392 20748 19398 20800
rect 20530 20748 20536 20800
rect 20588 20788 20594 20800
rect 20625 20791 20683 20797
rect 20625 20788 20637 20791
rect 20588 20760 20637 20788
rect 20588 20748 20594 20760
rect 20625 20757 20637 20760
rect 20671 20757 20683 20791
rect 20625 20751 20683 20757
rect 21913 20791 21971 20797
rect 21913 20757 21925 20791
rect 21959 20788 21971 20791
rect 22186 20788 22192 20800
rect 21959 20760 22192 20788
rect 21959 20757 21971 20760
rect 21913 20751 21971 20757
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 23753 20791 23811 20797
rect 23753 20757 23765 20791
rect 23799 20788 23811 20791
rect 23934 20788 23940 20800
rect 23799 20760 23940 20788
rect 23799 20757 23811 20760
rect 23753 20751 23811 20757
rect 23934 20748 23940 20760
rect 23992 20748 23998 20800
rect 29730 20748 29736 20800
rect 29788 20748 29794 20800
rect 30285 20791 30343 20797
rect 30285 20757 30297 20791
rect 30331 20788 30343 20791
rect 32306 20788 32312 20800
rect 30331 20760 32312 20788
rect 30331 20757 30343 20760
rect 30285 20751 30343 20757
rect 32306 20748 32312 20760
rect 32364 20748 32370 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7653 20587 7711 20593
rect 7653 20584 7665 20587
rect 6972 20556 7665 20584
rect 6972 20544 6978 20556
rect 7653 20553 7665 20556
rect 7699 20553 7711 20587
rect 7653 20547 7711 20553
rect 10502 20544 10508 20596
rect 10560 20544 10566 20596
rect 11146 20544 11152 20596
rect 11204 20584 11210 20596
rect 11517 20587 11575 20593
rect 11517 20584 11529 20587
rect 11204 20556 11529 20584
rect 11204 20544 11210 20556
rect 11517 20553 11529 20556
rect 11563 20553 11575 20587
rect 11517 20547 11575 20553
rect 13633 20587 13691 20593
rect 13633 20553 13645 20587
rect 13679 20584 13691 20587
rect 14090 20584 14096 20596
rect 13679 20556 14096 20584
rect 13679 20553 13691 20556
rect 13633 20547 13691 20553
rect 14090 20544 14096 20556
rect 14148 20544 14154 20596
rect 17310 20544 17316 20596
rect 17368 20584 17374 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17368 20556 17601 20584
rect 17368 20544 17374 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17589 20547 17647 20553
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19521 20587 19579 20593
rect 19521 20584 19533 20587
rect 19392 20556 19533 20584
rect 19392 20544 19398 20556
rect 19521 20553 19533 20556
rect 19567 20553 19579 20587
rect 19521 20547 19579 20553
rect 20625 20587 20683 20593
rect 20625 20553 20637 20587
rect 20671 20584 20683 20587
rect 21266 20584 21272 20596
rect 20671 20556 21272 20584
rect 20671 20553 20683 20556
rect 20625 20547 20683 20553
rect 21266 20544 21272 20556
rect 21324 20544 21330 20596
rect 32125 20587 32183 20593
rect 32125 20584 32137 20587
rect 22066 20556 32137 20584
rect 6638 20476 6644 20528
rect 6696 20516 6702 20528
rect 6733 20519 6791 20525
rect 6733 20516 6745 20519
rect 6696 20488 6745 20516
rect 6696 20476 6702 20488
rect 6733 20485 6745 20488
rect 6779 20485 6791 20519
rect 6733 20479 6791 20485
rect 8564 20519 8622 20525
rect 8564 20485 8576 20519
rect 8610 20516 8622 20519
rect 10137 20519 10195 20525
rect 10137 20516 10149 20519
rect 8610 20488 10149 20516
rect 8610 20485 8622 20488
rect 8564 20479 8622 20485
rect 10137 20485 10149 20488
rect 10183 20485 10195 20519
rect 10137 20479 10195 20485
rect 7098 20448 7104 20460
rect 7059 20420 7104 20448
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 10318 20408 10324 20460
rect 10376 20457 10382 20460
rect 10520 20457 10548 20544
rect 11330 20476 11336 20528
rect 11388 20516 11394 20528
rect 11701 20519 11759 20525
rect 11701 20516 11713 20519
rect 11388 20488 11713 20516
rect 11388 20476 11394 20488
rect 11701 20485 11713 20488
rect 11747 20485 11759 20519
rect 12802 20516 12808 20528
rect 12763 20488 12808 20516
rect 11701 20479 11759 20485
rect 12802 20476 12808 20488
rect 12860 20476 12866 20528
rect 12989 20519 13047 20525
rect 12989 20485 13001 20519
rect 13035 20516 13047 20519
rect 13078 20516 13084 20528
rect 13035 20488 13084 20516
rect 13035 20485 13047 20488
rect 12989 20479 13047 20485
rect 13078 20476 13084 20488
rect 13136 20516 13142 20528
rect 13906 20516 13912 20528
rect 13136 20488 13912 20516
rect 13136 20476 13142 20488
rect 13906 20476 13912 20488
rect 13964 20476 13970 20528
rect 18408 20519 18466 20525
rect 18408 20485 18420 20519
rect 18454 20516 18466 20519
rect 18506 20516 18512 20528
rect 18454 20488 18512 20516
rect 18454 20485 18466 20488
rect 18408 20479 18466 20485
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 21082 20516 21088 20528
rect 21043 20488 21088 20516
rect 21082 20476 21088 20488
rect 21140 20476 21146 20528
rect 10376 20451 10425 20457
rect 10376 20417 10379 20451
rect 10413 20417 10425 20451
rect 10376 20411 10425 20417
rect 10505 20451 10563 20457
rect 10505 20417 10517 20451
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 10597 20454 10655 20460
rect 10597 20420 10609 20454
rect 10643 20420 10655 20454
rect 10597 20414 10655 20420
rect 10376 20408 10382 20411
rect 7742 20340 7748 20392
rect 7800 20380 7806 20392
rect 8297 20383 8355 20389
rect 8297 20380 8309 20383
rect 7800 20352 8309 20380
rect 7800 20340 7806 20352
rect 8297 20349 8309 20352
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 10612 20324 10640 20414
rect 10778 20408 10784 20460
rect 10836 20448 10842 20460
rect 11885 20451 11943 20457
rect 10836 20420 10881 20448
rect 10836 20408 10842 20420
rect 11885 20417 11897 20451
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 10594 20272 10600 20324
rect 10652 20272 10658 20324
rect 11900 20312 11928 20411
rect 13262 20408 13268 20460
rect 13320 20448 13326 20460
rect 13449 20451 13507 20457
rect 13449 20448 13461 20451
rect 13320 20420 13461 20448
rect 13320 20408 13326 20420
rect 13449 20417 13461 20420
rect 13495 20417 13507 20451
rect 13449 20411 13507 20417
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20448 13691 20451
rect 14182 20448 14188 20460
rect 13679 20420 14188 20448
rect 13679 20417 13691 20420
rect 13633 20411 13691 20417
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 14734 20448 14740 20460
rect 14695 20420 14740 20448
rect 14734 20408 14740 20420
rect 14792 20408 14798 20460
rect 18138 20448 18144 20460
rect 18099 20420 18144 20448
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 22066 20448 22094 20556
rect 32125 20553 32137 20556
rect 32171 20553 32183 20587
rect 32125 20547 32183 20553
rect 22186 20525 22192 20528
rect 22180 20479 22192 20525
rect 22244 20516 22250 20528
rect 22244 20488 22280 20516
rect 22186 20476 22192 20479
rect 22244 20476 22250 20488
rect 23474 20476 23480 20528
rect 23532 20516 23538 20528
rect 23753 20519 23811 20525
rect 23753 20516 23765 20519
rect 23532 20488 23765 20516
rect 23532 20476 23538 20488
rect 23753 20485 23765 20488
rect 23799 20485 23811 20519
rect 29546 20516 29552 20528
rect 23753 20479 23811 20485
rect 29104 20488 29552 20516
rect 23934 20448 23940 20460
rect 18248 20420 22094 20448
rect 23895 20420 23940 20448
rect 14645 20383 14703 20389
rect 14645 20349 14657 20383
rect 14691 20380 14703 20383
rect 18248 20380 18276 20420
rect 23934 20408 23940 20420
rect 23992 20408 23998 20460
rect 24118 20448 24124 20460
rect 24079 20420 24124 20448
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 29104 20457 29132 20488
rect 29546 20476 29552 20488
rect 29604 20516 29610 20528
rect 30098 20516 30104 20528
rect 29604 20488 30104 20516
rect 29604 20476 29610 20488
rect 30098 20476 30104 20488
rect 30156 20476 30162 20528
rect 31570 20476 31576 20528
rect 31628 20516 31634 20528
rect 32585 20519 32643 20525
rect 31628 20488 32444 20516
rect 31628 20476 31634 20488
rect 29089 20451 29147 20457
rect 29089 20417 29101 20451
rect 29135 20417 29147 20451
rect 29089 20411 29147 20417
rect 29730 20408 29736 20460
rect 29788 20448 29794 20460
rect 32416 20457 32444 20488
rect 32585 20485 32597 20519
rect 32631 20516 32643 20519
rect 32858 20516 32864 20528
rect 32631 20488 32864 20516
rect 32631 20485 32643 20488
rect 32585 20479 32643 20485
rect 32858 20476 32864 20488
rect 32916 20476 32922 20528
rect 35989 20519 36047 20525
rect 35989 20485 36001 20519
rect 36035 20516 36047 20519
rect 36906 20516 36912 20528
rect 36035 20488 36912 20516
rect 36035 20485 36047 20488
rect 35989 20479 36047 20485
rect 36906 20476 36912 20488
rect 36964 20476 36970 20528
rect 30377 20451 30435 20457
rect 30377 20448 30389 20451
rect 29788 20420 30389 20448
rect 29788 20408 29794 20420
rect 30377 20417 30389 20420
rect 30423 20417 30435 20451
rect 30377 20411 30435 20417
rect 32309 20451 32367 20457
rect 32309 20417 32321 20451
rect 32355 20417 32367 20451
rect 32309 20411 32367 20417
rect 32401 20451 32459 20457
rect 32401 20417 32413 20451
rect 32447 20417 32459 20451
rect 35894 20448 35900 20460
rect 35855 20420 35900 20448
rect 32401 20411 32459 20417
rect 14691 20352 18276 20380
rect 21913 20383 21971 20389
rect 14691 20349 14703 20352
rect 14645 20343 14703 20349
rect 21913 20349 21925 20383
rect 21959 20349 21971 20383
rect 21913 20343 21971 20349
rect 12802 20312 12808 20324
rect 11900 20284 12808 20312
rect 12802 20272 12808 20284
rect 12860 20312 12866 20324
rect 15746 20312 15752 20324
rect 12860 20284 15752 20312
rect 12860 20272 12866 20284
rect 15746 20272 15752 20284
rect 15804 20272 15810 20324
rect 9677 20247 9735 20253
rect 9677 20213 9689 20247
rect 9723 20244 9735 20247
rect 10134 20244 10140 20256
rect 9723 20216 10140 20244
rect 9723 20213 9735 20216
rect 9677 20207 9735 20213
rect 10134 20204 10140 20216
rect 10192 20204 10198 20256
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 14369 20247 14427 20253
rect 14369 20244 14381 20247
rect 14332 20216 14381 20244
rect 14332 20204 14338 20216
rect 14369 20213 14381 20216
rect 14415 20213 14427 20247
rect 14369 20207 14427 20213
rect 14458 20204 14464 20256
rect 14516 20244 14522 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 14516 20216 14565 20244
rect 14516 20204 14522 20216
rect 14553 20213 14565 20216
rect 14599 20244 14611 20247
rect 15197 20247 15255 20253
rect 15197 20244 15209 20247
rect 14599 20216 15209 20244
rect 14599 20213 14611 20216
rect 14553 20207 14611 20213
rect 15197 20213 15209 20216
rect 15243 20213 15255 20247
rect 21928 20244 21956 20343
rect 28166 20340 28172 20392
rect 28224 20380 28230 20392
rect 28813 20383 28871 20389
rect 28813 20380 28825 20383
rect 28224 20352 28825 20380
rect 28224 20340 28230 20352
rect 28813 20349 28825 20352
rect 28859 20349 28871 20383
rect 28813 20343 28871 20349
rect 28994 20340 29000 20392
rect 29052 20380 29058 20392
rect 30101 20383 30159 20389
rect 30101 20380 30113 20383
rect 29052 20352 30113 20380
rect 29052 20340 29058 20352
rect 30101 20349 30113 20352
rect 30147 20349 30159 20383
rect 32324 20380 32352 20411
rect 35894 20408 35900 20420
rect 35952 20408 35958 20460
rect 36078 20448 36084 20460
rect 36039 20420 36084 20448
rect 36078 20408 36084 20420
rect 36136 20408 36142 20460
rect 36265 20451 36323 20457
rect 36265 20417 36277 20451
rect 36311 20448 36323 20451
rect 36630 20448 36636 20460
rect 36311 20420 36636 20448
rect 36311 20417 36323 20420
rect 36265 20411 36323 20417
rect 36630 20408 36636 20420
rect 36688 20408 36694 20460
rect 32324 20352 35756 20380
rect 30101 20343 30159 20349
rect 35728 20321 35756 20352
rect 35713 20315 35771 20321
rect 35713 20281 35725 20315
rect 35759 20281 35771 20315
rect 35713 20275 35771 20281
rect 36446 20272 36452 20324
rect 36504 20312 36510 20324
rect 36630 20312 36636 20324
rect 36504 20284 36636 20312
rect 36504 20272 36510 20284
rect 36630 20272 36636 20284
rect 36688 20272 36694 20324
rect 22094 20244 22100 20256
rect 21928 20216 22100 20244
rect 15197 20207 15255 20213
rect 22094 20204 22100 20216
rect 22152 20204 22158 20256
rect 23293 20247 23351 20253
rect 23293 20213 23305 20247
rect 23339 20244 23351 20247
rect 23750 20244 23756 20256
rect 23339 20216 23756 20244
rect 23339 20213 23351 20216
rect 23293 20207 23351 20213
rect 23750 20204 23756 20216
rect 23808 20204 23814 20256
rect 32306 20244 32312 20256
rect 32267 20216 32312 20244
rect 32306 20204 32312 20216
rect 32364 20204 32370 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 10045 20043 10103 20049
rect 10045 20009 10057 20043
rect 10091 20040 10103 20043
rect 10594 20040 10600 20052
rect 10091 20012 10600 20040
rect 10091 20009 10103 20012
rect 10045 20003 10103 20009
rect 10594 20000 10600 20012
rect 10652 20000 10658 20052
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 11606 20040 11612 20052
rect 11204 20012 11612 20040
rect 11204 20000 11210 20012
rect 11606 20000 11612 20012
rect 11664 20040 11670 20052
rect 11885 20043 11943 20049
rect 11885 20040 11897 20043
rect 11664 20012 11897 20040
rect 11664 20000 11670 20012
rect 11885 20009 11897 20012
rect 11931 20009 11943 20043
rect 11885 20003 11943 20009
rect 12158 20000 12164 20052
rect 12216 20040 12222 20052
rect 13078 20040 13084 20052
rect 12216 20012 13084 20040
rect 12216 20000 12222 20012
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 14182 20040 14188 20052
rect 14095 20012 14188 20040
rect 14182 20000 14188 20012
rect 14240 20040 14246 20052
rect 15102 20040 15108 20052
rect 14240 20012 15108 20040
rect 14240 20000 14246 20012
rect 15102 20000 15108 20012
rect 15160 20040 15166 20052
rect 18230 20040 18236 20052
rect 15160 20012 18236 20040
rect 15160 20000 15166 20012
rect 18230 20000 18236 20012
rect 18288 20000 18294 20052
rect 21266 20000 21272 20052
rect 21324 20040 21330 20052
rect 21821 20043 21879 20049
rect 21821 20040 21833 20043
rect 21324 20012 21833 20040
rect 21324 20000 21330 20012
rect 21821 20009 21833 20012
rect 21867 20009 21879 20043
rect 21821 20003 21879 20009
rect 22278 20000 22284 20052
rect 22336 20040 22342 20052
rect 22465 20043 22523 20049
rect 22465 20040 22477 20043
rect 22336 20012 22477 20040
rect 22336 20000 22342 20012
rect 22465 20009 22477 20012
rect 22511 20009 22523 20043
rect 22465 20003 22523 20009
rect 34790 20000 34796 20052
rect 34848 20040 34854 20052
rect 35069 20043 35127 20049
rect 35069 20040 35081 20043
rect 34848 20012 35081 20040
rect 34848 20000 34854 20012
rect 35069 20009 35081 20012
rect 35115 20009 35127 20043
rect 35069 20003 35127 20009
rect 39666 20000 39672 20052
rect 39724 20040 39730 20052
rect 40221 20043 40279 20049
rect 40221 20040 40233 20043
rect 39724 20012 40233 20040
rect 39724 20000 39730 20012
rect 40221 20009 40233 20012
rect 40267 20040 40279 20043
rect 40862 20040 40868 20052
rect 40267 20012 40868 20040
rect 40267 20009 40279 20012
rect 40221 20003 40279 20009
rect 40862 20000 40868 20012
rect 40920 20000 40926 20052
rect 5718 19932 5724 19984
rect 5776 19972 5782 19984
rect 6365 19975 6423 19981
rect 6365 19972 6377 19975
rect 5776 19944 6377 19972
rect 5776 19932 5782 19944
rect 6365 19941 6377 19944
rect 6411 19972 6423 19975
rect 13354 19972 13360 19984
rect 6411 19944 13360 19972
rect 6411 19941 6423 19944
rect 6365 19935 6423 19941
rect 13354 19932 13360 19944
rect 13412 19972 13418 19984
rect 14645 19975 14703 19981
rect 14645 19972 14657 19975
rect 13412 19944 14657 19972
rect 13412 19932 13418 19944
rect 14645 19941 14657 19944
rect 14691 19941 14703 19975
rect 36354 19972 36360 19984
rect 14645 19935 14703 19941
rect 35268 19944 36360 19972
rect 5629 19907 5687 19913
rect 5629 19873 5641 19907
rect 5675 19904 5687 19907
rect 7558 19904 7564 19916
rect 5675 19876 7564 19904
rect 5675 19873 5687 19876
rect 5629 19867 5687 19873
rect 7558 19864 7564 19876
rect 7616 19904 7622 19916
rect 11333 19907 11391 19913
rect 11333 19904 11345 19907
rect 7616 19876 11345 19904
rect 7616 19864 7622 19876
rect 11333 19873 11345 19876
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 2406 19796 2412 19848
rect 2464 19836 2470 19848
rect 2501 19839 2559 19845
rect 2501 19836 2513 19839
rect 2464 19808 2513 19836
rect 2464 19796 2470 19808
rect 2501 19805 2513 19808
rect 2547 19805 2559 19839
rect 2501 19799 2559 19805
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 4890 19836 4896 19848
rect 4764 19808 4896 19836
rect 4764 19796 4770 19808
rect 4890 19796 4896 19808
rect 4948 19836 4954 19848
rect 9585 19839 9643 19845
rect 9585 19836 9597 19839
rect 4948 19808 9597 19836
rect 4948 19796 4954 19808
rect 9585 19805 9597 19808
rect 9631 19836 9643 19839
rect 10318 19836 10324 19848
rect 9631 19808 10324 19836
rect 9631 19805 9643 19808
rect 9585 19799 9643 19805
rect 10318 19796 10324 19808
rect 10376 19836 10382 19848
rect 11348 19836 11376 19867
rect 12250 19864 12256 19916
rect 12308 19904 12314 19916
rect 13170 19904 13176 19916
rect 12308 19876 13176 19904
rect 12308 19864 12314 19876
rect 12820 19845 12848 19876
rect 13170 19864 13176 19876
rect 13228 19864 13234 19916
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 10376 19808 10548 19836
rect 11348 19808 12725 19836
rect 10376 19796 10382 19808
rect 3878 19728 3884 19780
rect 3936 19768 3942 19780
rect 4433 19771 4491 19777
rect 4433 19768 4445 19771
rect 3936 19740 4445 19768
rect 3936 19728 3942 19740
rect 4433 19737 4445 19740
rect 4479 19768 4491 19771
rect 5445 19771 5503 19777
rect 5445 19768 5457 19771
rect 4479 19740 5457 19768
rect 4479 19737 4491 19740
rect 4433 19731 4491 19737
rect 5445 19737 5457 19740
rect 5491 19768 5503 19771
rect 5718 19768 5724 19780
rect 5491 19740 5724 19768
rect 5491 19737 5503 19740
rect 5445 19731 5503 19737
rect 5718 19728 5724 19740
rect 5776 19728 5782 19780
rect 6178 19768 6184 19780
rect 6139 19740 6184 19768
rect 6178 19728 6184 19740
rect 6236 19728 6242 19780
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 10229 19771 10287 19777
rect 10229 19768 10241 19771
rect 10192 19740 10241 19768
rect 10192 19728 10198 19740
rect 10229 19737 10241 19740
rect 10275 19737 10287 19771
rect 10410 19768 10416 19780
rect 10371 19740 10416 19768
rect 10229 19731 10287 19737
rect 10410 19728 10416 19740
rect 10468 19728 10474 19780
rect 10520 19768 10548 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 12713 19799 12771 19805
rect 12805 19839 12863 19845
rect 12805 19805 12817 19839
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 12728 19768 12756 19799
rect 12894 19796 12900 19848
rect 12952 19836 12958 19848
rect 12952 19808 12997 19836
rect 12952 19796 12958 19808
rect 13078 19796 13084 19848
rect 13136 19836 13142 19848
rect 14660 19836 14688 19935
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 26329 19907 26387 19913
rect 26329 19904 26341 19907
rect 26292 19876 26341 19904
rect 26292 19864 26298 19876
rect 26329 19873 26341 19876
rect 26375 19873 26387 19907
rect 26329 19867 26387 19873
rect 15427 19839 15485 19845
rect 15427 19836 15439 19839
rect 13136 19808 13181 19836
rect 14660 19808 15439 19836
rect 13136 19796 13142 19808
rect 15427 19805 15439 19808
rect 15473 19805 15485 19839
rect 15562 19836 15568 19848
rect 15523 19808 15568 19836
rect 15427 19799 15485 19805
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15657 19839 15715 19845
rect 15657 19805 15669 19839
rect 15703 19805 15715 19839
rect 15657 19799 15715 19805
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19836 15899 19839
rect 16022 19836 16028 19848
rect 15887 19808 16028 19836
rect 15887 19805 15899 19808
rect 15841 19799 15899 19805
rect 13814 19768 13820 19780
rect 10520 19740 12664 19768
rect 12728 19740 13820 19768
rect 2130 19660 2136 19712
rect 2188 19700 2194 19712
rect 2317 19703 2375 19709
rect 2317 19700 2329 19703
rect 2188 19672 2329 19700
rect 2188 19660 2194 19672
rect 2317 19669 2329 19672
rect 2363 19669 2375 19703
rect 5736 19700 5764 19728
rect 6917 19703 6975 19709
rect 6917 19700 6929 19703
rect 5736 19672 6929 19700
rect 2317 19663 2375 19669
rect 6917 19669 6929 19672
rect 6963 19700 6975 19703
rect 7098 19700 7104 19712
rect 6963 19672 7104 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 12636 19700 12664 19740
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 15286 19768 15292 19780
rect 13924 19740 15292 19768
rect 13924 19700 13952 19740
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 15672 19768 15700 19799
rect 16022 19796 16028 19808
rect 16080 19796 16086 19848
rect 22649 19839 22707 19845
rect 22649 19805 22661 19839
rect 22695 19836 22707 19839
rect 23750 19836 23756 19848
rect 22695 19808 23756 19836
rect 22695 19805 22707 19808
rect 22649 19799 22707 19805
rect 23750 19796 23756 19808
rect 23808 19796 23814 19848
rect 30834 19796 30840 19848
rect 30892 19836 30898 19848
rect 30929 19839 30987 19845
rect 30929 19836 30941 19839
rect 30892 19808 30941 19836
rect 30892 19796 30898 19808
rect 30929 19805 30941 19808
rect 30975 19805 30987 19839
rect 30929 19799 30987 19805
rect 31754 19796 31760 19848
rect 31812 19836 31818 19848
rect 32674 19836 32680 19848
rect 31812 19808 32680 19836
rect 31812 19796 31818 19808
rect 32674 19796 32680 19808
rect 32732 19836 32738 19848
rect 35268 19845 35296 19944
rect 36354 19932 36360 19944
rect 36412 19932 36418 19984
rect 36262 19904 36268 19916
rect 35452 19876 36268 19904
rect 35452 19845 35480 19876
rect 36262 19864 36268 19876
rect 36320 19864 36326 19916
rect 32769 19839 32827 19845
rect 32769 19836 32781 19839
rect 32732 19808 32781 19836
rect 32732 19796 32738 19808
rect 32769 19805 32781 19808
rect 32815 19805 32827 19839
rect 32769 19799 32827 19805
rect 35253 19839 35311 19845
rect 35253 19805 35265 19839
rect 35299 19805 35311 19839
rect 35253 19799 35311 19805
rect 35437 19839 35495 19845
rect 35437 19805 35449 19839
rect 35483 19805 35495 19839
rect 35437 19799 35495 19805
rect 35621 19839 35679 19845
rect 35621 19805 35633 19839
rect 35667 19836 35679 19839
rect 35710 19836 35716 19848
rect 35667 19808 35716 19836
rect 35667 19805 35679 19808
rect 35621 19799 35679 19805
rect 35710 19796 35716 19808
rect 35768 19796 35774 19848
rect 58158 19836 58164 19848
rect 58119 19808 58164 19836
rect 58158 19796 58164 19808
rect 58216 19796 58222 19848
rect 16666 19768 16672 19780
rect 15672 19740 16672 19768
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 20070 19728 20076 19780
rect 20128 19768 20134 19780
rect 22833 19771 22891 19777
rect 22833 19768 22845 19771
rect 20128 19740 22845 19768
rect 20128 19728 20134 19740
rect 22833 19737 22845 19740
rect 22879 19768 22891 19771
rect 24118 19768 24124 19780
rect 22879 19740 24124 19768
rect 22879 19737 22891 19740
rect 22833 19731 22891 19737
rect 24118 19728 24124 19740
rect 24176 19728 24182 19780
rect 27614 19728 27620 19780
rect 27672 19768 27678 19780
rect 28077 19771 28135 19777
rect 28077 19768 28089 19771
rect 27672 19740 28089 19768
rect 27672 19728 27678 19740
rect 28077 19737 28089 19740
rect 28123 19768 28135 19771
rect 28537 19771 28595 19777
rect 28537 19768 28549 19771
rect 28123 19740 28549 19768
rect 28123 19737 28135 19740
rect 28077 19731 28135 19737
rect 28537 19737 28549 19740
rect 28583 19737 28595 19771
rect 31110 19768 31116 19780
rect 31071 19740 31116 19768
rect 28537 19731 28595 19737
rect 31110 19728 31116 19740
rect 31168 19768 31174 19780
rect 32582 19768 32588 19780
rect 31168 19740 32588 19768
rect 31168 19728 31174 19740
rect 32582 19728 32588 19740
rect 32640 19728 32646 19780
rect 35345 19771 35403 19777
rect 35345 19737 35357 19771
rect 35391 19737 35403 19771
rect 35345 19731 35403 19737
rect 12492 19672 12537 19700
rect 12636 19672 13952 19700
rect 15197 19703 15255 19709
rect 12492 19660 12498 19672
rect 15197 19669 15209 19703
rect 15243 19700 15255 19703
rect 17402 19700 17408 19712
rect 15243 19672 17408 19700
rect 15243 19669 15255 19672
rect 15197 19663 15255 19669
rect 17402 19660 17408 19672
rect 17460 19660 17466 19712
rect 30745 19703 30803 19709
rect 30745 19669 30757 19703
rect 30791 19700 30803 19703
rect 30834 19700 30840 19712
rect 30791 19672 30840 19700
rect 30791 19669 30803 19672
rect 30745 19663 30803 19669
rect 30834 19660 30840 19672
rect 30892 19660 30898 19712
rect 32858 19660 32864 19712
rect 32916 19700 32922 19712
rect 32953 19703 33011 19709
rect 32953 19700 32965 19703
rect 32916 19672 32965 19700
rect 32916 19660 32922 19672
rect 32953 19669 32965 19672
rect 32999 19669 33011 19703
rect 35360 19700 35388 19731
rect 38654 19700 38660 19712
rect 35360 19672 38660 19700
rect 32953 19663 33011 19669
rect 38654 19660 38660 19672
rect 38712 19660 38718 19712
rect 39850 19660 39856 19712
rect 39908 19700 39914 19712
rect 41046 19700 41052 19712
rect 39908 19672 41052 19700
rect 39908 19660 39914 19672
rect 41046 19660 41052 19672
rect 41104 19660 41110 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 2406 19496 2412 19508
rect 2367 19468 2412 19496
rect 2406 19456 2412 19468
rect 2464 19456 2470 19508
rect 3878 19496 3884 19508
rect 3839 19468 3884 19496
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 12805 19499 12863 19505
rect 10468 19468 12756 19496
rect 10468 19456 10474 19468
rect 10612 19437 10640 19468
rect 10597 19431 10655 19437
rect 10597 19397 10609 19431
rect 10643 19397 10655 19431
rect 10597 19391 10655 19397
rect 10781 19431 10839 19437
rect 10781 19397 10793 19431
rect 10827 19428 10839 19431
rect 10962 19428 10968 19440
rect 10827 19400 10968 19428
rect 10827 19397 10839 19400
rect 10781 19391 10839 19397
rect 10962 19388 10968 19400
rect 11020 19388 11026 19440
rect 12250 19428 12256 19440
rect 11900 19400 12256 19428
rect 2593 19363 2651 19369
rect 2593 19329 2605 19363
rect 2639 19360 2651 19363
rect 3786 19360 3792 19372
rect 2639 19332 3792 19360
rect 2639 19329 2651 19332
rect 2593 19323 2651 19329
rect 3786 19320 3792 19332
rect 3844 19320 3850 19372
rect 7926 19320 7932 19372
rect 7984 19320 7990 19372
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19360 10103 19363
rect 11514 19360 11520 19372
rect 10091 19332 11520 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11790 19360 11796 19372
rect 11751 19332 11796 19360
rect 11790 19320 11796 19332
rect 11848 19320 11854 19372
rect 11900 19369 11928 19400
rect 12250 19388 12256 19400
rect 12308 19388 12314 19440
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 12158 19360 12164 19372
rect 12119 19332 12164 19360
rect 11977 19323 12035 19329
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 2866 19292 2872 19304
rect 2823 19264 2872 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 3973 19295 4031 19301
rect 3973 19261 3985 19295
rect 4019 19261 4031 19295
rect 3973 19255 4031 19261
rect 3878 19184 3884 19236
rect 3936 19224 3942 19236
rect 3988 19224 4016 19255
rect 4062 19252 4068 19304
rect 4120 19292 4126 19304
rect 4120 19264 4165 19292
rect 4120 19252 4126 19264
rect 3936 19196 4016 19224
rect 3936 19184 3942 19196
rect 2590 19116 2596 19168
rect 2648 19156 2654 19168
rect 3513 19159 3571 19165
rect 3513 19156 3525 19159
rect 2648 19128 3525 19156
rect 2648 19116 2654 19128
rect 3513 19125 3525 19128
rect 3559 19125 3571 19159
rect 3513 19119 3571 19125
rect 4706 19116 4712 19168
rect 4764 19156 4770 19168
rect 5169 19159 5227 19165
rect 5169 19156 5181 19159
rect 4764 19128 5181 19156
rect 4764 19116 4770 19128
rect 5169 19125 5181 19128
rect 5215 19125 5227 19159
rect 5718 19156 5724 19168
rect 5679 19128 5724 19156
rect 5169 19119 5227 19125
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 6178 19116 6184 19168
rect 6236 19156 6242 19168
rect 6549 19159 6607 19165
rect 6549 19156 6561 19159
rect 6236 19128 6561 19156
rect 6236 19116 6242 19128
rect 6549 19125 6561 19128
rect 6595 19156 6607 19159
rect 7944 19156 7972 19320
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 10965 19295 11023 19301
rect 10965 19261 10977 19295
rect 11011 19292 11023 19295
rect 11992 19292 12020 19323
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 12728 19360 12756 19468
rect 12805 19465 12817 19499
rect 12851 19496 12863 19499
rect 12894 19496 12900 19508
rect 12851 19468 12900 19496
rect 12851 19465 12863 19468
rect 12805 19459 12863 19465
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 15562 19456 15568 19508
rect 15620 19456 15626 19508
rect 17770 19456 17776 19508
rect 17828 19496 17834 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 17828 19468 18337 19496
rect 17828 19456 17834 19468
rect 18325 19465 18337 19468
rect 18371 19496 18383 19499
rect 21726 19496 21732 19508
rect 18371 19468 21732 19496
rect 18371 19465 18383 19468
rect 18325 19459 18383 19465
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 27157 19499 27215 19505
rect 27157 19465 27169 19499
rect 27203 19496 27215 19499
rect 27706 19496 27712 19508
rect 27203 19468 27712 19496
rect 27203 19465 27215 19468
rect 27157 19459 27215 19465
rect 27706 19456 27712 19468
rect 27764 19456 27770 19508
rect 32674 19456 32680 19508
rect 32732 19496 32738 19508
rect 32769 19499 32827 19505
rect 32769 19496 32781 19499
rect 32732 19468 32781 19496
rect 32732 19456 32738 19468
rect 32769 19465 32781 19468
rect 32815 19465 32827 19499
rect 32769 19459 32827 19465
rect 38565 19499 38623 19505
rect 38565 19465 38577 19499
rect 38611 19496 38623 19499
rect 38654 19496 38660 19508
rect 38611 19468 38660 19496
rect 38611 19465 38623 19468
rect 38565 19459 38623 19465
rect 38654 19456 38660 19468
rect 38712 19456 38718 19508
rect 40494 19456 40500 19508
rect 40552 19456 40558 19508
rect 41046 19496 41052 19508
rect 41007 19468 41052 19496
rect 41046 19456 41052 19468
rect 41104 19456 41110 19508
rect 15580 19428 15608 19456
rect 16758 19428 16764 19440
rect 15488 19400 16764 19428
rect 12802 19360 12808 19372
rect 12728 19332 12808 19360
rect 11011 19264 12020 19292
rect 12728 19292 12756 19332
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 12989 19363 13047 19369
rect 12989 19329 13001 19363
rect 13035 19360 13047 19363
rect 13078 19360 13084 19372
rect 13035 19332 13084 19360
rect 13035 19329 13047 19332
rect 12989 19323 13047 19329
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19360 13231 19363
rect 13219 19332 13253 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 13188 19292 13216 19323
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 15488 19369 15516 19400
rect 16758 19388 16764 19400
rect 16816 19428 16822 19440
rect 16816 19400 17540 19428
rect 16816 19388 16822 19400
rect 15381 19363 15439 19369
rect 15381 19360 15393 19363
rect 13872 19332 15393 19360
rect 13872 19320 13878 19332
rect 14660 19301 14688 19332
rect 15381 19329 15393 19332
rect 15427 19329 15439 19363
rect 15381 19323 15439 19329
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 15749 19363 15807 19369
rect 15620 19332 15665 19360
rect 15620 19320 15626 19332
rect 15749 19329 15761 19363
rect 15795 19360 15807 19363
rect 16022 19360 16028 19372
rect 15795 19332 16028 19360
rect 15795 19329 15807 19332
rect 15749 19323 15807 19329
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 17512 19369 17540 19400
rect 17586 19388 17592 19440
rect 17644 19428 17650 19440
rect 29365 19431 29423 19437
rect 17644 19400 29224 19428
rect 17644 19388 17650 19400
rect 17497 19363 17555 19369
rect 17497 19329 17509 19363
rect 17543 19329 17555 19363
rect 18046 19360 18052 19372
rect 17497 19323 17555 19329
rect 17604 19332 18052 19360
rect 12728 19264 13216 19292
rect 14645 19295 14703 19301
rect 11011 19261 11023 19264
rect 10965 19255 11023 19261
rect 14645 19261 14657 19295
rect 14691 19261 14703 19295
rect 14645 19255 14703 19261
rect 9490 19184 9496 19236
rect 9548 19224 9554 19236
rect 9968 19224 9996 19255
rect 16482 19252 16488 19304
rect 16540 19292 16546 19304
rect 17604 19292 17632 19332
rect 18046 19320 18052 19332
rect 18104 19320 18110 19372
rect 18230 19360 18236 19372
rect 18143 19332 18236 19360
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 18417 19363 18475 19369
rect 18417 19329 18429 19363
rect 18463 19360 18475 19363
rect 18506 19360 18512 19372
rect 18463 19332 18512 19360
rect 18463 19329 18475 19332
rect 18417 19323 18475 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 20346 19320 20352 19372
rect 20404 19360 20410 19372
rect 29196 19369 29224 19400
rect 29365 19397 29377 19431
rect 29411 19428 29423 19431
rect 29730 19428 29736 19440
rect 29411 19400 29736 19428
rect 29411 19397 29423 19400
rect 29365 19391 29423 19397
rect 29730 19388 29736 19400
rect 29788 19388 29794 19440
rect 31297 19431 31355 19437
rect 30668 19400 31248 19428
rect 26973 19363 27031 19369
rect 26973 19360 26985 19363
rect 20404 19332 26985 19360
rect 20404 19320 20410 19332
rect 26973 19329 26985 19332
rect 27019 19329 27031 19363
rect 26973 19323 27031 19329
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19329 29239 19363
rect 29454 19360 29460 19372
rect 29415 19332 29460 19360
rect 29181 19323 29239 19329
rect 29454 19320 29460 19332
rect 29512 19320 29518 19372
rect 29546 19320 29552 19372
rect 29604 19360 29610 19372
rect 30668 19369 30696 19400
rect 30653 19363 30711 19369
rect 29604 19332 29649 19360
rect 29604 19320 29610 19332
rect 30653 19329 30665 19363
rect 30699 19329 30711 19363
rect 30834 19360 30840 19372
rect 30795 19332 30840 19360
rect 30653 19323 30711 19329
rect 30834 19320 30840 19332
rect 30892 19320 30898 19372
rect 30929 19363 30987 19369
rect 30929 19329 30941 19363
rect 30975 19329 30987 19363
rect 30929 19323 30987 19329
rect 17770 19292 17776 19304
rect 16540 19264 17632 19292
rect 17731 19264 17776 19292
rect 16540 19252 16546 19264
rect 17770 19252 17776 19264
rect 17828 19252 17834 19304
rect 18248 19292 18276 19320
rect 18877 19295 18935 19301
rect 18877 19292 18889 19295
rect 18248 19264 18889 19292
rect 18877 19261 18889 19264
rect 18923 19261 18935 19295
rect 18877 19255 18935 19261
rect 10226 19224 10232 19236
rect 9548 19196 9904 19224
rect 9968 19196 10232 19224
rect 9548 19184 9554 19196
rect 8478 19156 8484 19168
rect 6595 19128 8484 19156
rect 6595 19125 6607 19128
rect 6549 19119 6607 19125
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8570 19116 8576 19168
rect 8628 19156 8634 19168
rect 9876 19165 9904 19196
rect 10226 19184 10232 19196
rect 10284 19224 10290 19236
rect 30282 19224 30288 19236
rect 10284 19196 30288 19224
rect 10284 19184 10290 19196
rect 30282 19184 30288 19196
rect 30340 19184 30346 19236
rect 30944 19224 30972 19323
rect 31018 19320 31024 19372
rect 31076 19360 31082 19372
rect 31220 19360 31248 19400
rect 31297 19397 31309 19431
rect 31343 19428 31355 19431
rect 31938 19428 31944 19440
rect 31343 19400 31944 19428
rect 31343 19397 31355 19400
rect 31297 19391 31355 19397
rect 31938 19388 31944 19400
rect 31996 19388 32002 19440
rect 39700 19431 39758 19437
rect 39700 19397 39712 19431
rect 39746 19428 39758 19431
rect 39850 19428 39856 19440
rect 39746 19400 39856 19428
rect 39746 19397 39758 19400
rect 39700 19391 39758 19397
rect 39850 19388 39856 19400
rect 39908 19388 39914 19440
rect 32306 19360 32312 19372
rect 31076 19332 31121 19360
rect 31220 19332 32312 19360
rect 31076 19320 31082 19332
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 33318 19320 33324 19372
rect 33376 19360 33382 19372
rect 33882 19363 33940 19369
rect 33882 19360 33894 19363
rect 33376 19332 33894 19360
rect 33376 19320 33382 19332
rect 33882 19329 33894 19332
rect 33928 19329 33940 19363
rect 33882 19323 33940 19329
rect 34149 19363 34207 19369
rect 34149 19329 34161 19363
rect 34195 19360 34207 19363
rect 35342 19360 35348 19372
rect 34195 19332 35348 19360
rect 34195 19329 34207 19332
rect 34149 19323 34207 19329
rect 35342 19320 35348 19332
rect 35400 19320 35406 19372
rect 35897 19363 35955 19369
rect 35897 19329 35909 19363
rect 35943 19360 35955 19363
rect 35986 19360 35992 19372
rect 35943 19332 35992 19360
rect 35943 19329 35955 19332
rect 35897 19323 35955 19329
rect 35986 19320 35992 19332
rect 36044 19320 36050 19372
rect 39945 19363 40003 19369
rect 39945 19329 39957 19363
rect 39991 19360 40003 19363
rect 40034 19360 40040 19372
rect 39991 19332 40040 19360
rect 39991 19329 40003 19332
rect 39945 19323 40003 19329
rect 40034 19320 40040 19332
rect 40092 19320 40098 19372
rect 40402 19360 40408 19372
rect 40363 19332 40408 19360
rect 40402 19320 40408 19332
rect 40460 19320 40466 19372
rect 40512 19366 40540 19456
rect 40568 19369 40626 19375
rect 40568 19366 40580 19369
rect 40512 19338 40580 19366
rect 40568 19335 40580 19338
rect 40614 19335 40626 19369
rect 40568 19329 40626 19335
rect 40668 19369 40726 19375
rect 40668 19335 40680 19369
rect 40714 19335 40726 19369
rect 40668 19329 40726 19335
rect 40773 19363 40831 19369
rect 40773 19329 40785 19363
rect 40819 19360 40831 19363
rect 40862 19360 40868 19372
rect 40819 19332 40868 19360
rect 40819 19329 40831 19332
rect 31036 19292 31064 19320
rect 32122 19292 32128 19304
rect 31036 19264 32128 19292
rect 32122 19252 32128 19264
rect 32180 19252 32186 19304
rect 36173 19295 36231 19301
rect 36173 19261 36185 19295
rect 36219 19292 36231 19295
rect 36262 19292 36268 19304
rect 36219 19264 36268 19292
rect 36219 19261 36231 19264
rect 36173 19255 36231 19261
rect 36262 19252 36268 19264
rect 36320 19252 36326 19304
rect 40696 19236 40724 19329
rect 40773 19323 40831 19329
rect 40862 19320 40868 19332
rect 40920 19320 40926 19372
rect 31662 19224 31668 19236
rect 30944 19196 31668 19224
rect 31662 19184 31668 19196
rect 31720 19184 31726 19236
rect 40678 19184 40684 19236
rect 40736 19184 40742 19236
rect 9677 19159 9735 19165
rect 9677 19156 9689 19159
rect 8628 19128 9689 19156
rect 8628 19116 8634 19128
rect 9677 19125 9689 19128
rect 9723 19125 9735 19159
rect 9677 19119 9735 19125
rect 9861 19159 9919 19165
rect 9861 19125 9873 19159
rect 9907 19125 9919 19159
rect 11514 19156 11520 19168
rect 11475 19128 11520 19156
rect 9861 19119 9919 19125
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 15105 19159 15163 19165
rect 15105 19125 15117 19159
rect 15151 19156 15163 19159
rect 15378 19156 15384 19168
rect 15151 19128 15384 19156
rect 15151 19125 15163 19128
rect 15105 19119 15163 19125
rect 15378 19116 15384 19128
rect 15436 19116 15442 19168
rect 17218 19116 17224 19168
rect 17276 19156 17282 19168
rect 18874 19156 18880 19168
rect 17276 19128 18880 19156
rect 17276 19116 17282 19128
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 19150 19116 19156 19168
rect 19208 19156 19214 19168
rect 25774 19156 25780 19168
rect 19208 19128 25780 19156
rect 19208 19116 19214 19128
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 29638 19116 29644 19168
rect 29696 19156 29702 19168
rect 29733 19159 29791 19165
rect 29733 19156 29745 19159
rect 29696 19128 29745 19156
rect 29696 19116 29702 19128
rect 29733 19125 29745 19128
rect 29779 19125 29791 19159
rect 29733 19119 29791 19125
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 3786 18952 3792 18964
rect 3747 18924 3792 18952
rect 3786 18912 3792 18924
rect 3844 18912 3850 18964
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 5721 18955 5779 18961
rect 4120 18924 4384 18952
rect 4120 18912 4126 18924
rect 3237 18887 3295 18893
rect 3237 18853 3249 18887
rect 3283 18884 3295 18887
rect 3283 18856 4292 18884
rect 3283 18853 3295 18856
rect 3237 18847 3295 18853
rect 4264 18828 4292 18856
rect 4246 18816 4252 18828
rect 4159 18788 4252 18816
rect 4246 18776 4252 18788
rect 4304 18776 4310 18828
rect 4356 18825 4384 18924
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 9030 18952 9036 18964
rect 5767 18924 9036 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 10226 18952 10232 18964
rect 10187 18924 10232 18952
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 13078 18912 13084 18964
rect 13136 18952 13142 18964
rect 13354 18952 13360 18964
rect 13136 18924 13360 18952
rect 13136 18912 13142 18924
rect 13354 18912 13360 18924
rect 13412 18952 13418 18964
rect 13541 18955 13599 18961
rect 13541 18952 13553 18955
rect 13412 18924 13553 18952
rect 13412 18912 13418 18924
rect 13541 18921 13553 18924
rect 13587 18921 13599 18955
rect 13541 18915 13599 18921
rect 16669 18955 16727 18961
rect 16669 18921 16681 18955
rect 16715 18952 16727 18955
rect 16942 18952 16948 18964
rect 16715 18924 16948 18952
rect 16715 18921 16727 18924
rect 16669 18915 16727 18921
rect 16942 18912 16948 18924
rect 17000 18952 17006 18964
rect 17494 18952 17500 18964
rect 17000 18924 17500 18952
rect 17000 18912 17006 18924
rect 17494 18912 17500 18924
rect 17552 18912 17558 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 24302 18952 24308 18964
rect 17828 18924 24308 18952
rect 17828 18912 17834 18924
rect 24302 18912 24308 18924
rect 24360 18912 24366 18964
rect 30837 18955 30895 18961
rect 30837 18921 30849 18955
rect 30883 18952 30895 18955
rect 30926 18952 30932 18964
rect 30883 18924 30932 18952
rect 30883 18921 30895 18924
rect 30837 18915 30895 18921
rect 30926 18912 30932 18924
rect 30984 18912 30990 18964
rect 33318 18952 33324 18964
rect 33279 18924 33324 18952
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 40221 18955 40279 18961
rect 40221 18921 40233 18955
rect 40267 18952 40279 18955
rect 40494 18952 40500 18964
rect 40267 18924 40500 18952
rect 40267 18921 40279 18924
rect 40221 18915 40279 18921
rect 40494 18912 40500 18924
rect 40552 18912 40558 18964
rect 19978 18844 19984 18896
rect 20036 18884 20042 18896
rect 20438 18884 20444 18896
rect 20036 18856 20444 18884
rect 20036 18844 20042 18856
rect 20438 18844 20444 18856
rect 20496 18844 20502 18896
rect 28994 18884 29000 18896
rect 24596 18856 29000 18884
rect 4341 18819 4399 18825
rect 4341 18785 4353 18819
rect 4387 18785 4399 18819
rect 7742 18816 7748 18828
rect 7703 18788 7748 18816
rect 4341 18779 4399 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 18874 18776 18880 18828
rect 18932 18816 18938 18828
rect 19242 18816 19248 18828
rect 18932 18788 19248 18816
rect 18932 18776 18938 18788
rect 19242 18776 19248 18788
rect 19300 18776 19306 18828
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19392 18788 20392 18816
rect 19392 18776 19398 18788
rect 1854 18748 1860 18760
rect 1815 18720 1860 18748
rect 1854 18708 1860 18720
rect 1912 18708 1918 18760
rect 2130 18757 2136 18760
rect 2124 18748 2136 18757
rect 2091 18720 2136 18748
rect 2124 18711 2136 18720
rect 2130 18708 2136 18711
rect 2188 18708 2194 18760
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 12161 18751 12219 18757
rect 12161 18748 12173 18751
rect 9640 18720 12173 18748
rect 9640 18708 9646 18720
rect 12161 18717 12173 18720
rect 12207 18748 12219 18751
rect 13538 18748 13544 18760
rect 12207 18720 13544 18748
rect 12207 18717 12219 18720
rect 12161 18711 12219 18717
rect 13538 18708 13544 18720
rect 13596 18748 13602 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 13596 18720 15301 18748
rect 13596 18708 13602 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 15378 18708 15384 18760
rect 15436 18748 15442 18760
rect 15545 18751 15603 18757
rect 15545 18748 15557 18751
rect 15436 18720 15557 18748
rect 15436 18708 15442 18720
rect 15545 18717 15557 18720
rect 15591 18717 15603 18751
rect 15545 18711 15603 18717
rect 16482 18708 16488 18760
rect 16540 18748 16546 18760
rect 17402 18757 17408 18760
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 16540 18720 17141 18748
rect 16540 18708 16546 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17396 18748 17408 18757
rect 17363 18720 17408 18748
rect 17129 18711 17187 18717
rect 17396 18711 17408 18720
rect 17402 18708 17408 18711
rect 17460 18708 17466 18760
rect 19978 18757 19984 18760
rect 19976 18748 19984 18757
rect 19939 18720 19984 18748
rect 19976 18711 19984 18720
rect 19978 18708 19984 18711
rect 20036 18708 20042 18760
rect 20364 18757 20392 18788
rect 20073 18751 20131 18757
rect 20073 18717 20085 18751
rect 20119 18717 20131 18751
rect 20073 18711 20131 18717
rect 20348 18751 20406 18757
rect 20348 18717 20360 18751
rect 20394 18717 20406 18751
rect 20348 18711 20406 18717
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18748 20499 18751
rect 20990 18748 20996 18760
rect 20487 18720 20996 18748
rect 20487 18717 20499 18720
rect 20441 18711 20499 18717
rect 4706 18640 4712 18692
rect 4764 18680 4770 18692
rect 5813 18683 5871 18689
rect 5813 18680 5825 18683
rect 4764 18652 5825 18680
rect 4764 18640 4770 18652
rect 5813 18649 5825 18652
rect 5859 18649 5871 18683
rect 5813 18643 5871 18649
rect 6822 18640 6828 18692
rect 6880 18680 6886 18692
rect 12434 18689 12440 18692
rect 7478 18683 7536 18689
rect 7478 18680 7490 18683
rect 6880 18652 7490 18680
rect 6880 18640 6886 18652
rect 7478 18649 7490 18652
rect 7524 18649 7536 18683
rect 7478 18643 7536 18649
rect 12428 18643 12440 18689
rect 12492 18680 12498 18692
rect 12492 18652 12528 18680
rect 12434 18640 12440 18643
rect 12492 18640 12498 18652
rect 17586 18640 17592 18692
rect 17644 18680 17650 18692
rect 19334 18680 19340 18692
rect 17644 18652 19340 18680
rect 17644 18640 17650 18652
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 19886 18640 19892 18692
rect 19944 18680 19950 18692
rect 20079 18680 20107 18711
rect 20990 18708 20996 18720
rect 21048 18708 21054 18760
rect 23934 18708 23940 18760
rect 23992 18748 23998 18760
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 23992 18720 24409 18748
rect 23992 18708 23998 18720
rect 24397 18717 24409 18720
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 19944 18652 20107 18680
rect 20165 18683 20223 18689
rect 19944 18640 19950 18652
rect 20165 18649 20177 18683
rect 20211 18680 20223 18683
rect 20254 18680 20260 18692
rect 20211 18652 20260 18680
rect 20211 18649 20223 18652
rect 20165 18643 20223 18649
rect 20254 18640 20260 18652
rect 20312 18640 20318 18692
rect 24596 18689 24624 18856
rect 28994 18844 29000 18856
rect 29052 18844 29058 18896
rect 29546 18844 29552 18896
rect 29604 18844 29610 18896
rect 28166 18816 28172 18828
rect 24780 18788 28172 18816
rect 24780 18760 24808 18788
rect 28166 18776 28172 18788
rect 28224 18776 28230 18828
rect 29564 18816 29592 18844
rect 32217 18819 32275 18825
rect 29564 18788 29960 18816
rect 24762 18748 24768 18760
rect 24723 18720 24768 18748
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 25774 18708 25780 18760
rect 25832 18748 25838 18760
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 25832 18720 29561 18748
rect 25832 18708 25838 18720
rect 29549 18717 29561 18720
rect 29595 18717 29607 18751
rect 29730 18748 29736 18760
rect 29691 18720 29736 18748
rect 29549 18711 29607 18717
rect 29730 18708 29736 18720
rect 29788 18708 29794 18760
rect 29932 18757 29960 18788
rect 32217 18785 32229 18819
rect 32263 18816 32275 18819
rect 32766 18816 32772 18828
rect 32263 18788 32772 18816
rect 32263 18785 32275 18788
rect 32217 18779 32275 18785
rect 32766 18776 32772 18788
rect 32824 18816 32830 18828
rect 35342 18816 35348 18828
rect 32824 18788 35348 18816
rect 32824 18776 32830 18788
rect 35342 18776 35348 18788
rect 35400 18776 35406 18828
rect 35894 18776 35900 18828
rect 35952 18816 35958 18828
rect 36081 18819 36139 18825
rect 36081 18816 36093 18819
rect 35952 18788 36093 18816
rect 35952 18776 35958 18788
rect 36081 18785 36093 18788
rect 36127 18816 36139 18819
rect 36127 18788 37044 18816
rect 36127 18785 36139 18788
rect 36081 18779 36139 18785
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18717 29975 18751
rect 31938 18748 31944 18760
rect 31996 18757 32002 18760
rect 31908 18720 31944 18748
rect 29917 18711 29975 18717
rect 31938 18708 31944 18720
rect 31996 18711 32008 18757
rect 31996 18708 32002 18711
rect 32306 18708 32312 18760
rect 32364 18748 32370 18760
rect 32677 18751 32735 18757
rect 32677 18748 32689 18751
rect 32364 18720 32689 18748
rect 32364 18708 32370 18720
rect 32677 18717 32689 18720
rect 32723 18717 32735 18751
rect 32858 18748 32864 18760
rect 32819 18720 32864 18748
rect 32677 18711 32735 18717
rect 32858 18708 32864 18720
rect 32916 18708 32922 18760
rect 32953 18751 33011 18757
rect 32953 18717 32965 18751
rect 32999 18717 33011 18751
rect 32953 18711 33011 18717
rect 24581 18683 24639 18689
rect 24581 18680 24593 18683
rect 23952 18652 24593 18680
rect 23952 18624 23980 18652
rect 24581 18649 24593 18652
rect 24627 18649 24639 18683
rect 24581 18643 24639 18649
rect 24673 18683 24731 18689
rect 24673 18649 24685 18683
rect 24719 18680 24731 18683
rect 25038 18680 25044 18692
rect 24719 18652 25044 18680
rect 24719 18649 24731 18652
rect 24673 18643 24731 18649
rect 25038 18640 25044 18652
rect 25096 18680 25102 18692
rect 26145 18683 26203 18689
rect 26145 18680 26157 18683
rect 25096 18652 26157 18680
rect 25096 18640 25102 18652
rect 26145 18649 26157 18652
rect 26191 18649 26203 18683
rect 26145 18643 26203 18649
rect 26329 18683 26387 18689
rect 26329 18649 26341 18683
rect 26375 18680 26387 18683
rect 26375 18652 26924 18680
rect 26375 18649 26387 18652
rect 26329 18643 26387 18649
rect 4154 18612 4160 18624
rect 4115 18584 4160 18612
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 6178 18572 6184 18624
rect 6236 18612 6242 18624
rect 6365 18615 6423 18621
rect 6365 18612 6377 18615
rect 6236 18584 6377 18612
rect 6236 18572 6242 18584
rect 6365 18581 6377 18584
rect 6411 18581 6423 18615
rect 6365 18575 6423 18581
rect 8297 18615 8355 18621
rect 8297 18581 8309 18615
rect 8343 18612 8355 18615
rect 8386 18612 8392 18624
rect 8343 18584 8392 18612
rect 8343 18581 8355 18584
rect 8297 18575 8355 18581
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11333 18615 11391 18621
rect 11333 18612 11345 18615
rect 11112 18584 11345 18612
rect 11112 18572 11118 18584
rect 11333 18581 11345 18584
rect 11379 18612 11391 18615
rect 11790 18612 11796 18624
rect 11379 18584 11796 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11790 18572 11796 18584
rect 11848 18572 11854 18624
rect 18230 18572 18236 18624
rect 18288 18612 18294 18624
rect 18509 18615 18567 18621
rect 18509 18612 18521 18615
rect 18288 18584 18521 18612
rect 18288 18572 18294 18584
rect 18509 18581 18521 18584
rect 18555 18612 18567 18615
rect 19150 18612 19156 18624
rect 18555 18584 19156 18612
rect 18555 18581 18567 18584
rect 18509 18575 18567 18581
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 19426 18572 19432 18624
rect 19484 18612 19490 18624
rect 19797 18615 19855 18621
rect 19797 18612 19809 18615
rect 19484 18584 19809 18612
rect 19484 18572 19490 18584
rect 19797 18581 19809 18584
rect 19843 18581 19855 18615
rect 19797 18575 19855 18581
rect 20990 18572 20996 18624
rect 21048 18612 21054 18624
rect 21453 18615 21511 18621
rect 21453 18612 21465 18615
rect 21048 18584 21465 18612
rect 21048 18572 21054 18584
rect 21453 18581 21465 18584
rect 21499 18581 21511 18615
rect 23658 18612 23664 18624
rect 23619 18584 23664 18612
rect 21453 18575 21511 18581
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 23934 18572 23940 18624
rect 23992 18572 23998 18624
rect 24946 18612 24952 18624
rect 24907 18584 24952 18612
rect 24946 18572 24952 18584
rect 25004 18572 25010 18624
rect 25961 18615 26019 18621
rect 25961 18581 25973 18615
rect 26007 18612 26019 18615
rect 26050 18612 26056 18624
rect 26007 18584 26056 18612
rect 26007 18581 26019 18584
rect 25961 18575 26019 18581
rect 26050 18572 26056 18584
rect 26108 18572 26114 18624
rect 26786 18612 26792 18624
rect 26747 18584 26792 18612
rect 26786 18572 26792 18584
rect 26844 18572 26850 18624
rect 26896 18612 26924 18652
rect 26970 18640 26976 18692
rect 27028 18680 27034 18692
rect 27157 18683 27215 18689
rect 27028 18652 27073 18680
rect 27028 18640 27034 18652
rect 27157 18649 27169 18683
rect 27203 18680 27215 18683
rect 27430 18680 27436 18692
rect 27203 18652 27436 18680
rect 27203 18649 27215 18652
rect 27157 18643 27215 18649
rect 27172 18612 27200 18643
rect 27430 18640 27436 18652
rect 27488 18640 27494 18692
rect 29822 18640 29828 18692
rect 29880 18680 29886 18692
rect 29880 18652 29925 18680
rect 29880 18640 29886 18652
rect 31662 18640 31668 18692
rect 31720 18680 31726 18692
rect 32968 18680 32996 18711
rect 33042 18708 33048 18760
rect 33100 18748 33106 18760
rect 36354 18748 36360 18760
rect 33100 18720 33145 18748
rect 36315 18720 36360 18748
rect 33100 18708 33106 18720
rect 36354 18708 36360 18720
rect 36412 18708 36418 18760
rect 37016 18757 37044 18788
rect 37001 18751 37059 18757
rect 37001 18717 37013 18751
rect 37047 18717 37059 18751
rect 37001 18711 37059 18717
rect 37369 18751 37427 18757
rect 37369 18717 37381 18751
rect 37415 18748 37427 18751
rect 37642 18748 37648 18760
rect 37415 18720 37648 18748
rect 37415 18717 37427 18720
rect 37369 18711 37427 18717
rect 37642 18708 37648 18720
rect 37700 18708 37706 18760
rect 38654 18708 38660 18760
rect 38712 18748 38718 18760
rect 40037 18751 40095 18757
rect 40037 18748 40049 18751
rect 38712 18720 40049 18748
rect 38712 18708 38718 18720
rect 40037 18717 40049 18720
rect 40083 18717 40095 18751
rect 58158 18748 58164 18760
rect 58119 18720 58164 18748
rect 40037 18711 40095 18717
rect 58158 18708 58164 18720
rect 58216 18708 58222 18760
rect 31720 18652 32996 18680
rect 31720 18640 31726 18652
rect 36078 18640 36084 18692
rect 36136 18680 36142 18692
rect 36372 18680 36400 18708
rect 37093 18683 37151 18689
rect 37093 18680 37105 18683
rect 36136 18652 36400 18680
rect 37016 18652 37105 18680
rect 36136 18640 36142 18652
rect 37016 18624 37044 18652
rect 37093 18649 37105 18652
rect 37139 18649 37151 18683
rect 37093 18643 37151 18649
rect 37182 18640 37188 18692
rect 37240 18680 37246 18692
rect 37240 18652 37285 18680
rect 37240 18640 37246 18652
rect 39758 18640 39764 18692
rect 39816 18680 39822 18692
rect 39853 18683 39911 18689
rect 39853 18680 39865 18683
rect 39816 18652 39865 18680
rect 39816 18640 39822 18652
rect 39853 18649 39865 18652
rect 39899 18649 39911 18683
rect 39853 18643 39911 18649
rect 26896 18584 27200 18612
rect 30101 18615 30159 18621
rect 30101 18581 30113 18615
rect 30147 18612 30159 18615
rect 30466 18612 30472 18624
rect 30147 18584 30472 18612
rect 30147 18581 30159 18584
rect 30101 18575 30159 18581
rect 30466 18572 30472 18584
rect 30524 18572 30530 18624
rect 36814 18612 36820 18624
rect 36775 18584 36820 18612
rect 36814 18572 36820 18584
rect 36872 18572 36878 18624
rect 36998 18572 37004 18624
rect 37056 18572 37062 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 4617 18411 4675 18417
rect 4617 18408 4629 18411
rect 4212 18380 4629 18408
rect 4212 18368 4218 18380
rect 4617 18377 4629 18380
rect 4663 18408 4675 18411
rect 6086 18408 6092 18420
rect 4663 18380 6092 18408
rect 4663 18377 4675 18380
rect 4617 18371 4675 18377
rect 6086 18368 6092 18380
rect 6144 18368 6150 18420
rect 6822 18408 6828 18420
rect 6783 18380 6828 18408
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 8113 18411 8171 18417
rect 8113 18377 8125 18411
rect 8159 18408 8171 18411
rect 10042 18408 10048 18420
rect 8159 18380 10048 18408
rect 8159 18377 8171 18380
rect 8113 18371 8171 18377
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 12250 18368 12256 18420
rect 12308 18408 12314 18420
rect 16114 18408 16120 18420
rect 12308 18380 16120 18408
rect 12308 18368 12314 18380
rect 16114 18368 16120 18380
rect 16172 18368 16178 18420
rect 16666 18408 16672 18420
rect 16627 18380 16672 18408
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 17034 18368 17040 18420
rect 17092 18408 17098 18420
rect 17218 18408 17224 18420
rect 17092 18380 17224 18408
rect 17092 18368 17098 18380
rect 17218 18368 17224 18380
rect 17276 18368 17282 18420
rect 18325 18411 18383 18417
rect 18325 18377 18337 18411
rect 18371 18408 18383 18411
rect 18966 18408 18972 18420
rect 18371 18380 18972 18408
rect 18371 18377 18383 18380
rect 18325 18371 18383 18377
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 20346 18408 20352 18420
rect 19628 18380 20352 18408
rect 1854 18300 1860 18352
rect 1912 18340 1918 18352
rect 2774 18340 2780 18352
rect 1912 18312 2780 18340
rect 1912 18300 1918 18312
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 2424 18281 2452 18312
rect 2774 18300 2780 18312
rect 2832 18300 2838 18352
rect 8570 18340 8576 18352
rect 7392 18312 8576 18340
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18241 2467 18275
rect 2665 18275 2723 18281
rect 2665 18272 2677 18275
rect 2409 18235 2467 18241
rect 2516 18244 2677 18272
rect 2516 18204 2544 18244
rect 2665 18241 2677 18244
rect 2711 18241 2723 18275
rect 2665 18235 2723 18241
rect 4246 18232 4252 18284
rect 4304 18272 4310 18284
rect 5445 18275 5503 18281
rect 5445 18272 5457 18275
rect 4304 18244 5457 18272
rect 4304 18232 4310 18244
rect 5445 18241 5457 18244
rect 5491 18241 5503 18275
rect 5445 18235 5503 18241
rect 6178 18232 6184 18284
rect 6236 18272 6242 18284
rect 7392 18281 7420 18312
rect 8570 18300 8576 18312
rect 8628 18300 8634 18352
rect 9852 18343 9910 18349
rect 9852 18309 9864 18343
rect 9898 18340 9910 18343
rect 11514 18340 11520 18352
rect 9898 18312 11520 18340
rect 9898 18309 9910 18312
rect 9852 18303 9910 18309
rect 11514 18300 11520 18312
rect 11572 18300 11578 18352
rect 15562 18300 15568 18352
rect 15620 18340 15626 18352
rect 15749 18343 15807 18349
rect 15749 18340 15761 18343
rect 15620 18312 15761 18340
rect 15620 18300 15626 18312
rect 15749 18309 15761 18312
rect 15795 18309 15807 18343
rect 18598 18340 18604 18352
rect 15749 18303 15807 18309
rect 15856 18312 18604 18340
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 6236 18244 7021 18272
rect 6236 18232 6242 18244
rect 7009 18241 7021 18244
rect 7055 18241 7067 18275
rect 7009 18235 7067 18241
rect 7377 18275 7435 18281
rect 7377 18241 7389 18275
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18272 7619 18275
rect 7926 18272 7932 18284
rect 7607 18244 7932 18272
rect 7607 18241 7619 18244
rect 7561 18235 7619 18241
rect 7926 18232 7932 18244
rect 7984 18232 7990 18284
rect 8386 18272 8392 18284
rect 8347 18244 8392 18272
rect 8386 18232 8392 18244
rect 8444 18232 8450 18284
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 15856 18272 15884 18312
rect 18598 18300 18604 18312
rect 18656 18300 18662 18352
rect 19426 18340 19432 18352
rect 18708 18312 19432 18340
rect 9364 18244 15884 18272
rect 15933 18275 15991 18281
rect 9364 18232 9370 18244
rect 15933 18241 15945 18275
rect 15979 18272 15991 18275
rect 16117 18275 16175 18281
rect 15979 18244 16068 18272
rect 15979 18241 15991 18244
rect 15933 18235 15991 18241
rect 1964 18176 2544 18204
rect 5077 18207 5135 18213
rect 1964 18145 1992 18176
rect 5077 18173 5089 18207
rect 5123 18204 5135 18207
rect 5166 18204 5172 18216
rect 5123 18176 5172 18204
rect 5123 18173 5135 18176
rect 5077 18167 5135 18173
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 5534 18204 5540 18216
rect 5495 18176 5540 18204
rect 5534 18164 5540 18176
rect 5592 18164 5598 18216
rect 7098 18164 7104 18216
rect 7156 18204 7162 18216
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 7156 18176 7205 18204
rect 7156 18164 7162 18176
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 7193 18167 7251 18173
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 1949 18139 2007 18145
rect 1949 18105 1961 18139
rect 1995 18105 2007 18139
rect 1949 18099 2007 18105
rect 5721 18139 5779 18145
rect 5721 18105 5733 18139
rect 5767 18136 5779 18139
rect 7300 18136 7328 18167
rect 5767 18108 7328 18136
rect 5767 18105 5779 18108
rect 5721 18099 5779 18105
rect 3786 18068 3792 18080
rect 3747 18040 3792 18068
rect 3786 18028 3792 18040
rect 3844 18028 3850 18080
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 8404 18068 8432 18232
rect 9582 18204 9588 18216
rect 9543 18176 9588 18204
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 16040 18136 16068 18244
rect 16117 18241 16129 18275
rect 16163 18241 16175 18275
rect 16850 18272 16856 18284
rect 16811 18244 16856 18272
rect 16117 18235 16175 18241
rect 16132 18204 16160 18235
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 17034 18272 17040 18284
rect 16995 18244 17040 18272
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 17770 18272 17776 18284
rect 17731 18244 17776 18272
rect 17770 18232 17776 18244
rect 17828 18232 17834 18284
rect 18708 18281 18736 18312
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 19521 18343 19579 18349
rect 19521 18309 19533 18343
rect 19567 18340 19579 18343
rect 19628 18340 19656 18380
rect 20346 18368 20352 18380
rect 20404 18368 20410 18420
rect 20530 18368 20536 18420
rect 20588 18368 20594 18420
rect 21913 18411 21971 18417
rect 21913 18377 21925 18411
rect 21959 18408 21971 18411
rect 24210 18408 24216 18420
rect 21959 18380 24216 18408
rect 21959 18377 21971 18380
rect 21913 18371 21971 18377
rect 24210 18368 24216 18380
rect 24268 18368 24274 18420
rect 25038 18408 25044 18420
rect 24999 18380 25044 18408
rect 25038 18368 25044 18380
rect 25096 18368 25102 18420
rect 29181 18411 29239 18417
rect 29181 18408 29193 18411
rect 25148 18380 29193 18408
rect 19567 18312 19656 18340
rect 19567 18309 19579 18312
rect 19521 18303 19579 18309
rect 19702 18300 19708 18352
rect 19760 18340 19766 18352
rect 19760 18312 20392 18340
rect 19760 18300 19766 18312
rect 17865 18275 17923 18281
rect 17865 18241 17877 18275
rect 17911 18241 17923 18275
rect 17865 18235 17923 18241
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18241 18751 18275
rect 19242 18272 19248 18284
rect 19203 18244 19248 18272
rect 18693 18235 18751 18241
rect 17052 18204 17080 18232
rect 16132 18176 17080 18204
rect 16942 18136 16948 18148
rect 16040 18108 16948 18136
rect 16942 18096 16948 18108
rect 17000 18096 17006 18148
rect 17880 18136 17908 18235
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 19337 18275 19395 18281
rect 19337 18241 19349 18275
rect 19383 18272 19395 18275
rect 19978 18272 19984 18284
rect 19383 18244 19984 18272
rect 19383 18241 19395 18244
rect 19337 18235 19395 18241
rect 19978 18232 19984 18244
rect 20036 18272 20042 18284
rect 20121 18275 20179 18281
rect 20121 18272 20133 18275
rect 20036 18244 20133 18272
rect 20036 18232 20042 18244
rect 20121 18241 20133 18244
rect 20167 18241 20179 18275
rect 20254 18272 20260 18284
rect 20215 18244 20260 18272
rect 20121 18235 20179 18241
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 20364 18281 20392 18312
rect 20547 18281 20575 18368
rect 25148 18340 25176 18380
rect 29181 18377 29193 18380
rect 29227 18377 29239 18411
rect 32582 18408 32588 18420
rect 32495 18380 32588 18408
rect 29181 18371 29239 18377
rect 32582 18368 32588 18380
rect 32640 18408 32646 18420
rect 33042 18408 33048 18420
rect 32640 18380 33048 18408
rect 32640 18368 32646 18380
rect 33042 18368 33048 18380
rect 33100 18368 33106 18420
rect 35253 18411 35311 18417
rect 35253 18377 35265 18411
rect 35299 18408 35311 18411
rect 35342 18408 35348 18420
rect 35299 18380 35348 18408
rect 35299 18377 35311 18380
rect 35253 18371 35311 18377
rect 35342 18368 35348 18380
rect 35400 18368 35406 18420
rect 38010 18408 38016 18420
rect 37292 18380 38016 18408
rect 20925 18312 25176 18340
rect 20349 18275 20407 18281
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 20532 18275 20590 18281
rect 20532 18241 20544 18275
rect 20578 18241 20590 18275
rect 20532 18235 20590 18241
rect 20622 18232 20628 18284
rect 20680 18272 20686 18284
rect 20680 18244 20725 18272
rect 20680 18232 20686 18244
rect 18601 18207 18659 18213
rect 18601 18173 18613 18207
rect 18647 18204 18659 18207
rect 20806 18204 20812 18216
rect 18647 18176 20812 18204
rect 18647 18173 18659 18176
rect 18601 18167 18659 18173
rect 20806 18164 20812 18176
rect 20864 18164 20870 18216
rect 19981 18139 20039 18145
rect 19981 18136 19993 18139
rect 17880 18108 19993 18136
rect 19981 18105 19993 18108
rect 20027 18105 20039 18139
rect 19981 18099 20039 18105
rect 10962 18068 10968 18080
rect 4672 18040 8432 18068
rect 10923 18040 10968 18068
rect 4672 18028 4678 18040
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11698 18068 11704 18080
rect 11659 18040 11704 18068
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 17402 18028 17408 18080
rect 17460 18068 17466 18080
rect 17497 18071 17555 18077
rect 17497 18068 17509 18071
rect 17460 18040 17509 18068
rect 17460 18028 17466 18040
rect 17497 18037 17509 18040
rect 17543 18037 17555 18071
rect 17678 18068 17684 18080
rect 17639 18040 17684 18068
rect 17497 18031 17555 18037
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 18414 18028 18420 18080
rect 18472 18068 18478 18080
rect 18509 18071 18567 18077
rect 18509 18068 18521 18071
rect 18472 18040 18521 18068
rect 18472 18028 18478 18040
rect 18509 18037 18521 18040
rect 18555 18037 18567 18071
rect 18509 18031 18567 18037
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 20925 18068 20953 18312
rect 25774 18300 25780 18352
rect 25832 18340 25838 18352
rect 27338 18340 27344 18352
rect 25832 18312 27344 18340
rect 25832 18300 25838 18312
rect 27338 18300 27344 18312
rect 27396 18340 27402 18352
rect 27890 18340 27896 18352
rect 27396 18312 27896 18340
rect 27396 18300 27402 18312
rect 27890 18300 27896 18312
rect 27948 18340 27954 18352
rect 27948 18312 30144 18340
rect 27948 18300 27954 18312
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21048 18244 21833 18272
rect 21048 18232 21054 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22005 18275 22063 18281
rect 22005 18241 22017 18275
rect 22051 18241 22063 18275
rect 23750 18272 23756 18284
rect 23711 18244 23756 18272
rect 22005 18235 22063 18241
rect 21726 18204 21732 18216
rect 21192 18176 21732 18204
rect 21192 18080 21220 18176
rect 21726 18164 21732 18176
rect 21784 18204 21790 18216
rect 22020 18204 22048 18235
rect 23750 18232 23756 18244
rect 23808 18232 23814 18284
rect 23934 18272 23940 18284
rect 23847 18244 23940 18272
rect 23934 18232 23940 18244
rect 23992 18232 23998 18284
rect 24029 18275 24087 18281
rect 24029 18241 24041 18275
rect 24075 18241 24087 18275
rect 24029 18235 24087 18241
rect 24121 18275 24179 18281
rect 24121 18241 24133 18275
rect 24167 18272 24179 18275
rect 24670 18272 24676 18284
rect 24167 18244 24676 18272
rect 24167 18241 24179 18244
rect 24121 18235 24179 18241
rect 22462 18204 22468 18216
rect 21784 18176 22048 18204
rect 22423 18176 22468 18204
rect 21784 18164 21790 18176
rect 22462 18164 22468 18176
rect 22520 18164 22526 18216
rect 22741 18207 22799 18213
rect 22741 18173 22753 18207
rect 22787 18204 22799 18207
rect 23952 18204 23980 18232
rect 22787 18176 23980 18204
rect 22787 18173 22799 18176
rect 22741 18167 22799 18173
rect 24044 18136 24072 18235
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 25682 18232 25688 18284
rect 25740 18272 25746 18284
rect 26154 18275 26212 18281
rect 26154 18272 26166 18275
rect 25740 18244 26166 18272
rect 25740 18232 25746 18244
rect 26154 18241 26166 18244
rect 26200 18241 26212 18275
rect 26154 18235 26212 18241
rect 26326 18232 26332 18284
rect 26384 18272 26390 18284
rect 26421 18275 26479 18281
rect 26421 18272 26433 18275
rect 26384 18244 26433 18272
rect 26384 18232 26390 18244
rect 26421 18241 26433 18244
rect 26467 18272 26479 18275
rect 26973 18275 27031 18281
rect 26973 18272 26985 18275
rect 26467 18244 26985 18272
rect 26467 18241 26479 18244
rect 26421 18235 26479 18241
rect 26973 18241 26985 18244
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 27062 18232 27068 18284
rect 27120 18272 27126 18284
rect 30116 18281 30144 18312
rect 35986 18300 35992 18352
rect 36044 18340 36050 18352
rect 36541 18343 36599 18349
rect 36541 18340 36553 18343
rect 36044 18312 36553 18340
rect 36044 18300 36050 18312
rect 36541 18309 36553 18312
rect 36587 18340 36599 18343
rect 37182 18340 37188 18352
rect 36587 18312 37188 18340
rect 36587 18309 36599 18312
rect 36541 18303 36599 18309
rect 37182 18300 37188 18312
rect 37240 18300 37246 18352
rect 27240 18275 27298 18281
rect 27240 18272 27252 18275
rect 27120 18244 27252 18272
rect 27120 18232 27126 18244
rect 27240 18241 27252 18244
rect 27286 18241 27298 18275
rect 27240 18235 27298 18241
rect 29365 18275 29423 18281
rect 29365 18241 29377 18275
rect 29411 18241 29423 18275
rect 29365 18235 29423 18241
rect 29641 18275 29699 18281
rect 29641 18241 29653 18275
rect 29687 18272 29699 18275
rect 30101 18275 30159 18281
rect 29687 18244 30052 18272
rect 29687 18241 29699 18244
rect 29641 18235 29699 18241
rect 29380 18136 29408 18235
rect 29549 18207 29607 18213
rect 29549 18173 29561 18207
rect 29595 18204 29607 18207
rect 29730 18204 29736 18216
rect 29595 18176 29736 18204
rect 29595 18173 29607 18176
rect 29549 18167 29607 18173
rect 29730 18164 29736 18176
rect 29788 18164 29794 18216
rect 30024 18204 30052 18244
rect 30101 18241 30113 18275
rect 30147 18241 30159 18275
rect 31202 18272 31208 18284
rect 30101 18235 30159 18241
rect 30300 18244 31208 18272
rect 30300 18204 30328 18244
rect 31202 18232 31208 18244
rect 31260 18232 31266 18284
rect 33502 18232 33508 18284
rect 33560 18272 33566 18284
rect 33965 18275 34023 18281
rect 33965 18272 33977 18275
rect 33560 18244 33977 18272
rect 33560 18232 33566 18244
rect 33965 18241 33977 18244
rect 34011 18241 34023 18275
rect 33965 18235 34023 18241
rect 35894 18232 35900 18284
rect 35952 18272 35958 18284
rect 36357 18275 36415 18281
rect 36357 18272 36369 18275
rect 35952 18244 36369 18272
rect 35952 18232 35958 18244
rect 36357 18241 36369 18244
rect 36403 18241 36415 18275
rect 36357 18235 36415 18241
rect 36446 18232 36452 18284
rect 36504 18272 36510 18284
rect 36725 18275 36783 18281
rect 36504 18244 36549 18272
rect 36504 18232 36510 18244
rect 36725 18241 36737 18275
rect 36771 18272 36783 18275
rect 37292 18272 37320 18380
rect 38010 18368 38016 18380
rect 38068 18368 38074 18420
rect 39758 18300 39764 18352
rect 39816 18340 39822 18352
rect 40957 18343 41015 18349
rect 40957 18340 40969 18343
rect 39816 18312 40969 18340
rect 39816 18300 39822 18312
rect 40957 18309 40969 18312
rect 41003 18309 41015 18343
rect 40957 18303 41015 18309
rect 36771 18244 37320 18272
rect 37369 18275 37427 18281
rect 36771 18241 36783 18244
rect 36725 18235 36783 18241
rect 37369 18241 37381 18275
rect 37415 18241 37427 18275
rect 39850 18272 39856 18284
rect 39908 18281 39914 18284
rect 39820 18244 39856 18272
rect 37369 18235 37427 18241
rect 30024 18176 30328 18204
rect 30377 18207 30435 18213
rect 30377 18173 30389 18207
rect 30423 18204 30435 18207
rect 31662 18204 31668 18216
rect 30423 18176 31668 18204
rect 30423 18173 30435 18176
rect 30377 18167 30435 18173
rect 31662 18164 31668 18176
rect 31720 18164 31726 18216
rect 36173 18139 36231 18145
rect 36173 18136 36185 18139
rect 24044 18108 25544 18136
rect 29380 18108 36185 18136
rect 21174 18068 21180 18080
rect 18656 18040 20953 18068
rect 21135 18040 21180 18068
rect 18656 18028 18662 18040
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 24305 18071 24363 18077
rect 24305 18037 24317 18071
rect 24351 18068 24363 18071
rect 24578 18068 24584 18080
rect 24351 18040 24584 18068
rect 24351 18037 24363 18040
rect 24305 18031 24363 18037
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 25516 18068 25544 18108
rect 36173 18105 36185 18108
rect 36219 18105 36231 18139
rect 36173 18099 36231 18105
rect 37090 18096 37096 18148
rect 37148 18136 37154 18148
rect 37384 18136 37412 18235
rect 39850 18232 39856 18244
rect 39908 18235 39920 18281
rect 39908 18232 39914 18235
rect 40034 18232 40040 18284
rect 40092 18272 40098 18284
rect 40129 18275 40187 18281
rect 40129 18272 40141 18275
rect 40092 18244 40141 18272
rect 40092 18232 40098 18244
rect 40129 18241 40141 18244
rect 40175 18241 40187 18275
rect 40773 18275 40831 18281
rect 40773 18272 40785 18275
rect 40129 18235 40187 18241
rect 40236 18244 40785 18272
rect 37550 18136 37556 18148
rect 37148 18108 37412 18136
rect 37511 18108 37556 18136
rect 37148 18096 37154 18108
rect 37550 18096 37556 18108
rect 37608 18096 37614 18148
rect 39022 18136 39028 18148
rect 38580 18108 39028 18136
rect 26970 18068 26976 18080
rect 25516 18040 26976 18068
rect 26970 18028 26976 18040
rect 27028 18068 27034 18080
rect 28353 18071 28411 18077
rect 28353 18068 28365 18071
rect 27028 18040 28365 18068
rect 27028 18028 27034 18040
rect 28353 18037 28365 18040
rect 28399 18037 28411 18071
rect 29638 18068 29644 18080
rect 29599 18040 29644 18068
rect 28353 18031 28411 18037
rect 29638 18028 29644 18040
rect 29696 18028 29702 18080
rect 33502 18068 33508 18080
rect 33463 18040 33508 18068
rect 33502 18028 33508 18040
rect 33560 18068 33566 18080
rect 38580 18068 38608 18108
rect 39022 18096 39028 18108
rect 39080 18096 39086 18148
rect 38746 18068 38752 18080
rect 33560 18040 38608 18068
rect 38707 18040 38752 18068
rect 33560 18028 33566 18040
rect 38746 18028 38752 18040
rect 38804 18068 38810 18080
rect 40236 18068 40264 18244
rect 40773 18241 40785 18244
rect 40819 18241 40831 18275
rect 40773 18235 40831 18241
rect 40586 18068 40592 18080
rect 38804 18040 40264 18068
rect 40547 18040 40592 18068
rect 38804 18028 38810 18040
rect 40586 18028 40592 18040
rect 40644 18028 40650 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2409 17867 2467 17873
rect 2409 17864 2421 17867
rect 1820 17836 2421 17864
rect 1820 17824 1826 17836
rect 2409 17833 2421 17836
rect 2455 17833 2467 17867
rect 4614 17864 4620 17876
rect 4575 17836 4620 17864
rect 2409 17827 2467 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 9214 17864 9220 17876
rect 9175 17836 9220 17864
rect 9214 17824 9220 17836
rect 9272 17824 9278 17876
rect 11241 17867 11299 17873
rect 11241 17833 11253 17867
rect 11287 17864 11299 17867
rect 11422 17864 11428 17876
rect 11287 17836 11428 17864
rect 11287 17833 11299 17836
rect 11241 17827 11299 17833
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 18601 17867 18659 17873
rect 18601 17833 18613 17867
rect 18647 17864 18659 17867
rect 20070 17864 20076 17876
rect 18647 17836 20076 17864
rect 18647 17833 18659 17836
rect 18601 17827 18659 17833
rect 18616 17796 18644 17827
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 21174 17864 21180 17876
rect 20456 17836 21180 17864
rect 20456 17796 20484 17836
rect 21174 17824 21180 17836
rect 21232 17824 21238 17876
rect 25682 17864 25688 17876
rect 25643 17836 25688 17864
rect 25682 17824 25688 17836
rect 25740 17824 25746 17876
rect 27062 17824 27068 17876
rect 27120 17864 27126 17876
rect 27433 17867 27491 17873
rect 27433 17864 27445 17867
rect 27120 17836 27445 17864
rect 27120 17824 27126 17836
rect 27433 17833 27445 17836
rect 27479 17833 27491 17867
rect 30282 17864 30288 17876
rect 30243 17836 30288 17864
rect 27433 17827 27491 17833
rect 30282 17824 30288 17836
rect 30340 17824 30346 17876
rect 30466 17864 30472 17876
rect 30427 17836 30472 17864
rect 30466 17824 30472 17836
rect 30524 17824 30530 17876
rect 31726 17836 35296 17864
rect 22462 17796 22468 17808
rect 17788 17768 18644 17796
rect 19720 17768 20484 17796
rect 20548 17768 22468 17796
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17728 2835 17731
rect 2866 17728 2872 17740
rect 2823 17700 2872 17728
rect 2823 17697 2835 17700
rect 2777 17691 2835 17697
rect 2866 17688 2872 17700
rect 2924 17728 2930 17740
rect 2924 17700 3648 17728
rect 2924 17688 2930 17700
rect 2590 17660 2596 17672
rect 2551 17632 2596 17660
rect 2590 17620 2596 17632
rect 2648 17620 2654 17672
rect 3620 17660 3648 17700
rect 3786 17688 3792 17740
rect 3844 17728 3850 17740
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 3844 17700 5457 17728
rect 3844 17688 3850 17700
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 5445 17691 5503 17697
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17728 8447 17731
rect 9582 17728 9588 17740
rect 8435 17700 9588 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 9582 17688 9588 17700
rect 9640 17688 9646 17740
rect 10226 17688 10232 17740
rect 10284 17728 10290 17740
rect 13538 17728 13544 17740
rect 10284 17700 13436 17728
rect 13499 17700 13544 17728
rect 10284 17688 10290 17700
rect 3878 17660 3884 17672
rect 3620 17632 3884 17660
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 5534 17660 5540 17672
rect 5447 17632 5540 17660
rect 5534 17620 5540 17632
rect 5592 17660 5598 17672
rect 5902 17660 5908 17672
rect 5592 17632 5908 17660
rect 5592 17620 5598 17632
rect 5902 17620 5908 17632
rect 5960 17620 5966 17672
rect 9306 17660 9312 17672
rect 9267 17632 9312 17660
rect 9306 17620 9312 17632
rect 9364 17620 9370 17672
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 9456 17632 9501 17660
rect 9456 17620 9462 17632
rect 10502 17620 10508 17672
rect 10560 17660 10566 17672
rect 11256 17669 11284 17700
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 10560 17632 11069 17660
rect 10560 17620 10566 17632
rect 11057 17629 11069 17632
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 13408 17660 13436 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 17494 17660 17500 17672
rect 13408 17632 17500 17660
rect 11241 17623 11299 17629
rect 17494 17620 17500 17632
rect 17552 17620 17558 17672
rect 17788 17669 17816 17768
rect 18046 17688 18052 17740
rect 18104 17728 18110 17740
rect 19720 17728 19748 17768
rect 18104 17700 19748 17728
rect 19797 17731 19855 17737
rect 18104 17688 18110 17700
rect 19797 17697 19809 17731
rect 19843 17728 19855 17731
rect 19978 17728 19984 17740
rect 19843 17700 19984 17728
rect 19843 17697 19855 17700
rect 19797 17691 19855 17697
rect 19978 17688 19984 17700
rect 20036 17688 20042 17740
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18230 17660 18236 17672
rect 18012 17632 18236 17660
rect 18012 17620 18018 17632
rect 18230 17620 18236 17632
rect 18288 17620 18294 17672
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 18506 17660 18512 17672
rect 18463 17632 18512 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 20070 17660 20076 17672
rect 20031 17632 20076 17660
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20548 17669 20576 17768
rect 22462 17756 22468 17768
rect 22520 17756 22526 17808
rect 24210 17756 24216 17808
rect 24268 17796 24274 17808
rect 28718 17796 28724 17808
rect 24268 17768 28724 17796
rect 24268 17756 24274 17768
rect 28718 17756 28724 17768
rect 28776 17756 28782 17808
rect 29733 17799 29791 17805
rect 29733 17765 29745 17799
rect 29779 17796 29791 17799
rect 31110 17796 31116 17808
rect 29779 17768 31116 17796
rect 29779 17765 29791 17768
rect 29733 17759 29791 17765
rect 31110 17756 31116 17768
rect 31168 17756 31174 17808
rect 27614 17728 27620 17740
rect 23676 17700 27620 17728
rect 23676 17672 23704 17700
rect 27614 17688 27620 17700
rect 27672 17688 27678 17740
rect 31726 17728 31754 17836
rect 35268 17796 35296 17836
rect 35342 17824 35348 17876
rect 35400 17864 35406 17876
rect 38746 17864 38752 17876
rect 35400 17836 38752 17864
rect 35400 17824 35406 17836
rect 38746 17824 38752 17836
rect 38804 17824 38810 17876
rect 39850 17864 39856 17876
rect 39811 17836 39856 17864
rect 39850 17824 39856 17836
rect 39908 17824 39914 17876
rect 36814 17796 36820 17808
rect 35268 17768 36820 17796
rect 36814 17756 36820 17768
rect 36872 17756 36878 17808
rect 37918 17728 37924 17740
rect 30484 17700 31754 17728
rect 35452 17700 37924 17728
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17629 20591 17663
rect 20809 17663 20867 17669
rect 20809 17660 20821 17663
rect 20533 17623 20591 17629
rect 20640 17632 20821 17660
rect 5721 17595 5779 17601
rect 5721 17561 5733 17595
rect 5767 17592 5779 17595
rect 5767 17564 7236 17592
rect 5767 17561 5779 17564
rect 5721 17555 5779 17561
rect 5077 17527 5135 17533
rect 5077 17493 5089 17527
rect 5123 17524 5135 17527
rect 5166 17524 5172 17536
rect 5123 17496 5172 17524
rect 5123 17493 5135 17496
rect 5077 17487 5135 17493
rect 5166 17484 5172 17496
rect 5224 17484 5230 17536
rect 6178 17484 6184 17536
rect 6236 17524 6242 17536
rect 6457 17527 6515 17533
rect 6457 17524 6469 17527
rect 6236 17496 6469 17524
rect 6236 17484 6242 17496
rect 6457 17493 6469 17496
rect 6503 17493 6515 17527
rect 6457 17487 6515 17493
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 7009 17527 7067 17533
rect 7009 17524 7021 17527
rect 6696 17496 7021 17524
rect 6696 17484 6702 17496
rect 7009 17493 7021 17496
rect 7055 17493 7067 17527
rect 7208 17524 7236 17564
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 8122 17595 8180 17601
rect 8122 17592 8134 17595
rect 7340 17564 8134 17592
rect 7340 17552 7346 17564
rect 8122 17561 8134 17564
rect 8168 17561 8180 17595
rect 8122 17555 8180 17561
rect 10042 17552 10048 17604
rect 10100 17592 10106 17604
rect 11330 17592 11336 17604
rect 10100 17564 11336 17592
rect 10100 17552 10106 17564
rect 11330 17552 11336 17564
rect 11388 17552 11394 17604
rect 11698 17552 11704 17604
rect 11756 17592 11762 17604
rect 11793 17595 11851 17601
rect 11793 17592 11805 17595
rect 11756 17564 11805 17592
rect 11756 17552 11762 17564
rect 11793 17561 11805 17564
rect 11839 17592 11851 17595
rect 12250 17592 12256 17604
rect 11839 17564 12256 17592
rect 11839 17561 11851 17564
rect 11793 17555 11851 17561
rect 12250 17552 12256 17564
rect 12308 17552 12314 17604
rect 12710 17552 12716 17604
rect 12768 17592 12774 17604
rect 20548 17592 20576 17623
rect 12768 17564 20576 17592
rect 12768 17552 12774 17564
rect 7650 17524 7656 17536
rect 7208 17496 7656 17524
rect 7009 17487 7067 17493
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 7800 17496 9045 17524
rect 7800 17484 7806 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 9033 17487 9091 17493
rect 9953 17527 10011 17533
rect 9953 17493 9965 17527
rect 9999 17524 10011 17527
rect 10226 17524 10232 17536
rect 9999 17496 10232 17524
rect 9999 17493 10011 17496
rect 9953 17487 10011 17493
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 10502 17524 10508 17536
rect 10463 17496 10508 17524
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 17034 17484 17040 17536
rect 17092 17524 17098 17536
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 17092 17496 17601 17524
rect 17092 17484 17098 17496
rect 17589 17493 17601 17496
rect 17635 17524 17647 17527
rect 17770 17524 17776 17536
rect 17635 17496 17776 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 17770 17484 17776 17496
rect 17828 17484 17834 17536
rect 18506 17484 18512 17536
rect 18564 17524 18570 17536
rect 20640 17524 20668 17632
rect 20809 17629 20821 17632
rect 20855 17660 20867 17663
rect 21082 17660 21088 17672
rect 20855 17632 21088 17660
rect 20855 17629 20867 17632
rect 20809 17623 20867 17629
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17660 23627 17663
rect 23658 17660 23664 17672
rect 23615 17632 23664 17660
rect 23615 17629 23627 17632
rect 23569 17623 23627 17629
rect 23658 17620 23664 17632
rect 23716 17620 23722 17672
rect 24394 17660 24400 17672
rect 24355 17632 24400 17660
rect 24394 17620 24400 17632
rect 24452 17620 24458 17672
rect 24670 17660 24676 17672
rect 24631 17632 24676 17660
rect 24670 17620 24676 17632
rect 24728 17620 24734 17672
rect 25866 17620 25872 17672
rect 25924 17654 25930 17672
rect 25961 17663 26019 17669
rect 25961 17654 25973 17663
rect 25924 17629 25973 17654
rect 26007 17629 26019 17663
rect 25924 17626 26019 17629
rect 25924 17620 25930 17626
rect 25961 17623 26019 17626
rect 26053 17663 26111 17669
rect 26053 17629 26065 17663
rect 26099 17629 26111 17663
rect 26053 17623 26111 17629
rect 26145 17663 26203 17669
rect 26145 17629 26157 17663
rect 26191 17660 26203 17663
rect 26234 17660 26240 17672
rect 26191 17632 26240 17660
rect 26191 17629 26203 17632
rect 26145 17623 26203 17629
rect 18564 17496 20668 17524
rect 18564 17484 18570 17496
rect 22094 17484 22100 17536
rect 22152 17524 22158 17536
rect 22152 17496 22197 17524
rect 22152 17484 22158 17496
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 26077 17524 26105 17623
rect 26234 17620 26240 17632
rect 26292 17620 26298 17672
rect 26329 17663 26387 17669
rect 26329 17629 26341 17663
rect 26375 17660 26387 17663
rect 26510 17660 26516 17672
rect 26375 17632 26516 17660
rect 26375 17629 26387 17632
rect 26329 17623 26387 17629
rect 26510 17620 26516 17632
rect 26568 17660 26574 17672
rect 26789 17663 26847 17669
rect 26789 17660 26801 17663
rect 26568 17632 26801 17660
rect 26568 17620 26574 17632
rect 26789 17629 26801 17632
rect 26835 17629 26847 17663
rect 26789 17623 26847 17629
rect 26878 17620 26884 17672
rect 26936 17660 26942 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26936 17632 26985 17660
rect 26936 17620 26942 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 26973 17623 27031 17629
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17629 27123 17663
rect 27065 17623 27123 17629
rect 27157 17663 27215 17669
rect 27157 17629 27169 17663
rect 27203 17662 27215 17663
rect 27246 17662 27252 17672
rect 27203 17634 27252 17662
rect 27203 17629 27215 17634
rect 27157 17623 27215 17629
rect 25832 17496 26105 17524
rect 27080 17524 27108 17623
rect 27246 17620 27252 17634
rect 27304 17620 27310 17672
rect 27430 17620 27436 17672
rect 27488 17660 27494 17672
rect 30484 17669 30512 17700
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 27488 17632 29561 17660
rect 27488 17620 27494 17632
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 29549 17623 29607 17629
rect 30469 17663 30527 17669
rect 30469 17629 30481 17663
rect 30515 17629 30527 17663
rect 30469 17623 30527 17629
rect 30558 17620 30564 17672
rect 30616 17660 30622 17672
rect 30742 17660 30748 17672
rect 30616 17632 30661 17660
rect 30703 17632 30748 17660
rect 30616 17620 30622 17632
rect 30742 17620 30748 17632
rect 30800 17620 30806 17672
rect 35069 17663 35127 17669
rect 35069 17629 35081 17663
rect 35115 17629 35127 17663
rect 35069 17623 35127 17629
rect 35161 17663 35219 17669
rect 35161 17629 35173 17663
rect 35207 17660 35219 17663
rect 35342 17660 35348 17672
rect 35207 17632 35348 17660
rect 35207 17629 35219 17632
rect 35161 17623 35219 17629
rect 27982 17552 27988 17604
rect 28040 17592 28046 17604
rect 34974 17592 34980 17604
rect 28040 17564 34980 17592
rect 28040 17552 28046 17564
rect 34974 17552 34980 17564
rect 35032 17552 35038 17604
rect 27338 17524 27344 17536
rect 27080 17496 27344 17524
rect 25832 17484 25838 17496
rect 27338 17484 27344 17496
rect 27396 17484 27402 17536
rect 29914 17484 29920 17536
rect 29972 17524 29978 17536
rect 34885 17527 34943 17533
rect 34885 17524 34897 17527
rect 29972 17496 34897 17524
rect 29972 17484 29978 17496
rect 34885 17493 34897 17496
rect 34931 17493 34943 17527
rect 35084 17524 35112 17623
rect 35342 17620 35348 17632
rect 35400 17620 35406 17672
rect 35452 17669 35480 17700
rect 37918 17688 37924 17700
rect 37976 17728 37982 17740
rect 40957 17731 41015 17737
rect 40957 17728 40969 17731
rect 37976 17700 38792 17728
rect 37976 17688 37982 17700
rect 35437 17663 35495 17669
rect 35437 17629 35449 17663
rect 35483 17629 35495 17663
rect 36078 17660 36084 17672
rect 35437 17623 35495 17629
rect 35544 17632 36084 17660
rect 35250 17552 35256 17604
rect 35308 17592 35314 17604
rect 35308 17564 35353 17592
rect 35308 17552 35314 17564
rect 35544 17524 35572 17632
rect 36078 17620 36084 17632
rect 36136 17620 36142 17672
rect 36354 17620 36360 17672
rect 36412 17660 36418 17672
rect 36449 17663 36507 17669
rect 36449 17660 36461 17663
rect 36412 17632 36461 17660
rect 36412 17620 36418 17632
rect 36449 17629 36461 17632
rect 36495 17629 36507 17663
rect 37093 17663 37151 17669
rect 37093 17660 37105 17663
rect 36449 17623 36507 17629
rect 36556 17632 37105 17660
rect 36170 17592 36176 17604
rect 36131 17564 36176 17592
rect 36170 17552 36176 17564
rect 36228 17552 36234 17604
rect 36262 17552 36268 17604
rect 36320 17592 36326 17604
rect 36320 17564 36365 17592
rect 36320 17552 36326 17564
rect 35894 17524 35900 17536
rect 35084 17496 35572 17524
rect 35855 17496 35900 17524
rect 34885 17487 34943 17493
rect 35894 17484 35900 17496
rect 35952 17484 35958 17536
rect 36078 17484 36084 17536
rect 36136 17524 36142 17536
rect 36556 17524 36584 17632
rect 37093 17629 37105 17632
rect 37139 17629 37151 17663
rect 37274 17660 37280 17672
rect 37235 17632 37280 17660
rect 37093 17623 37151 17629
rect 37274 17620 37280 17632
rect 37332 17620 37338 17672
rect 37458 17660 37464 17672
rect 37419 17632 37464 17660
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 38764 17669 38792 17700
rect 40144 17700 40969 17728
rect 38749 17663 38807 17669
rect 38749 17629 38761 17663
rect 38795 17629 38807 17663
rect 38749 17623 38807 17629
rect 38838 17620 38844 17672
rect 38896 17660 38902 17672
rect 40144 17669 40172 17700
rect 40957 17697 40969 17700
rect 41003 17697 41015 17731
rect 40957 17691 41015 17697
rect 40129 17663 40187 17669
rect 40129 17660 40141 17663
rect 38896 17632 40141 17660
rect 38896 17620 38902 17632
rect 40129 17629 40141 17632
rect 40175 17629 40187 17663
rect 40129 17623 40187 17629
rect 40218 17657 40276 17663
rect 40218 17623 40230 17657
rect 40264 17623 40276 17657
rect 40218 17617 40276 17623
rect 40313 17660 40371 17666
rect 40313 17626 40325 17660
rect 40359 17626 40371 17660
rect 40313 17620 40371 17626
rect 40494 17620 40500 17672
rect 40552 17660 40558 17672
rect 40552 17632 40597 17660
rect 40552 17620 40558 17632
rect 37185 17595 37243 17601
rect 37185 17561 37197 17595
rect 37231 17561 37243 17595
rect 38562 17592 38568 17604
rect 38523 17564 38568 17592
rect 37185 17555 37243 17561
rect 36906 17524 36912 17536
rect 36136 17496 36584 17524
rect 36867 17496 36912 17524
rect 36136 17484 36142 17496
rect 36906 17484 36912 17496
rect 36964 17484 36970 17536
rect 37200 17524 37228 17555
rect 38562 17552 38568 17564
rect 38620 17552 38626 17604
rect 37826 17524 37832 17536
rect 37200 17496 37832 17524
rect 37826 17484 37832 17496
rect 37884 17484 37890 17536
rect 38933 17527 38991 17533
rect 38933 17493 38945 17527
rect 38979 17524 38991 17527
rect 39206 17524 39212 17536
rect 38979 17496 39212 17524
rect 38979 17493 38991 17496
rect 38933 17487 38991 17493
rect 39206 17484 39212 17496
rect 39264 17484 39270 17536
rect 40236 17524 40264 17617
rect 40328 17592 40356 17620
rect 40586 17592 40592 17604
rect 40328 17564 40592 17592
rect 40586 17552 40592 17564
rect 40644 17552 40650 17604
rect 40678 17524 40684 17536
rect 40236 17496 40684 17524
rect 40678 17484 40684 17496
rect 40736 17484 40742 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 3881 17323 3939 17329
rect 3881 17289 3893 17323
rect 3927 17320 3939 17323
rect 4890 17320 4896 17332
rect 3927 17292 4896 17320
rect 3927 17289 3939 17292
rect 3881 17283 3939 17289
rect 4890 17280 4896 17292
rect 4948 17280 4954 17332
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5445 17323 5503 17329
rect 5445 17320 5457 17323
rect 5316 17292 5457 17320
rect 5316 17280 5322 17292
rect 5445 17289 5457 17292
rect 5491 17289 5503 17323
rect 5445 17283 5503 17289
rect 7193 17323 7251 17329
rect 7193 17289 7205 17323
rect 7239 17320 7251 17323
rect 7282 17320 7288 17332
rect 7239 17292 7288 17320
rect 7239 17289 7251 17292
rect 7193 17283 7251 17289
rect 7282 17280 7288 17292
rect 7340 17280 7346 17332
rect 9306 17320 9312 17332
rect 9267 17292 9312 17320
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 9398 17280 9404 17332
rect 9456 17320 9462 17332
rect 12897 17323 12955 17329
rect 12897 17320 12909 17323
rect 9456 17292 12909 17320
rect 9456 17280 9462 17292
rect 12897 17289 12909 17292
rect 12943 17289 12955 17323
rect 19978 17320 19984 17332
rect 12897 17283 12955 17289
rect 13096 17292 19984 17320
rect 10229 17255 10287 17261
rect 10229 17221 10241 17255
rect 10275 17252 10287 17255
rect 10686 17252 10692 17264
rect 10275 17224 10692 17252
rect 10275 17221 10287 17224
rect 10229 17215 10287 17221
rect 10686 17212 10692 17224
rect 10744 17212 10750 17264
rect 11609 17255 11667 17261
rect 11609 17221 11621 17255
rect 11655 17252 11667 17255
rect 11882 17252 11888 17264
rect 11655 17224 11888 17252
rect 11655 17221 11667 17224
rect 11609 17215 11667 17221
rect 11882 17212 11888 17224
rect 11940 17212 11946 17264
rect 13096 17252 13124 17292
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20625 17323 20683 17329
rect 20625 17320 20637 17323
rect 20220 17292 20637 17320
rect 20220 17280 20226 17292
rect 20625 17289 20637 17292
rect 20671 17289 20683 17323
rect 20625 17283 20683 17289
rect 21913 17323 21971 17329
rect 21913 17289 21925 17323
rect 21959 17320 21971 17323
rect 24210 17320 24216 17332
rect 21959 17292 24216 17320
rect 21959 17289 21971 17292
rect 21913 17283 21971 17289
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 24489 17323 24547 17329
rect 24489 17289 24501 17323
rect 24535 17289 24547 17323
rect 26602 17320 26608 17332
rect 24489 17283 24547 17289
rect 24596 17292 26608 17320
rect 13262 17252 13268 17264
rect 11992 17224 13124 17252
rect 13223 17224 13268 17252
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4614 17184 4620 17196
rect 4479 17156 4620 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 3237 17119 3295 17125
rect 3237 17085 3249 17119
rect 3283 17116 3295 17119
rect 3712 17116 3740 17147
rect 4614 17144 4620 17156
rect 4672 17184 4678 17196
rect 4890 17184 4896 17196
rect 4672 17156 4896 17184
rect 4672 17144 4678 17156
rect 4890 17144 4896 17156
rect 4948 17144 4954 17196
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5316 17156 5733 17184
rect 5316 17144 5322 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 5721 17147 5779 17153
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 7377 17187 7435 17193
rect 7377 17184 7389 17187
rect 6696 17156 7389 17184
rect 6696 17144 6702 17156
rect 7377 17153 7389 17156
rect 7423 17153 7435 17187
rect 7742 17184 7748 17196
rect 7703 17156 7748 17184
rect 7377 17147 7435 17153
rect 7742 17144 7748 17156
rect 7800 17144 7806 17196
rect 7926 17184 7932 17196
rect 7887 17156 7932 17184
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 10042 17193 10048 17196
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9824 17156 9873 17184
rect 9824 17144 9830 17156
rect 9861 17153 9873 17156
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 10009 17187 10048 17193
rect 10009 17153 10021 17187
rect 10009 17147 10048 17153
rect 10042 17144 10048 17147
rect 10100 17144 10106 17196
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 10326 17187 10384 17193
rect 10326 17153 10338 17187
rect 10372 17153 10384 17187
rect 10326 17147 10384 17153
rect 4706 17116 4712 17128
rect 3283 17088 4712 17116
rect 3283 17085 3295 17088
rect 3237 17079 3295 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 7098 17076 7104 17128
rect 7156 17116 7162 17128
rect 7282 17116 7288 17128
rect 7156 17088 7288 17116
rect 7156 17076 7162 17088
rect 7282 17076 7288 17088
rect 7340 17116 7346 17128
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 7340 17088 7573 17116
rect 7340 17076 7346 17088
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 7650 17076 7656 17128
rect 7708 17116 7714 17128
rect 7708 17088 7753 17116
rect 7708 17076 7714 17088
rect 4617 17051 4675 17057
rect 4617 17017 4629 17051
rect 4663 17048 4675 17051
rect 4798 17048 4804 17060
rect 4663 17020 4804 17048
rect 4663 17017 4675 17020
rect 4617 17011 4675 17017
rect 4798 17008 4804 17020
rect 4856 17048 4862 17060
rect 9674 17048 9680 17060
rect 4856 17020 9680 17048
rect 4856 17008 4862 17020
rect 9674 17008 9680 17020
rect 9732 17008 9738 17060
rect 10152 17048 10180 17147
rect 10341 17116 10369 17147
rect 11330 17144 11336 17196
rect 11388 17184 11394 17196
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11388 17156 11529 17184
rect 11388 17144 11394 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 11517 17147 11575 17153
rect 11698 17144 11704 17156
rect 11756 17184 11762 17196
rect 11992 17184 12020 17224
rect 13262 17212 13268 17224
rect 13320 17212 13326 17264
rect 18414 17212 18420 17264
rect 18472 17252 18478 17264
rect 18782 17252 18788 17264
rect 18472 17224 18788 17252
rect 18472 17212 18478 17224
rect 18782 17212 18788 17224
rect 18840 17212 18846 17264
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 24504 17252 24532 17283
rect 20864 17224 24532 17252
rect 20864 17212 20870 17224
rect 11756 17156 12020 17184
rect 13037 17187 13095 17193
rect 11756 17144 11762 17156
rect 13037 17153 13049 17187
rect 13083 17153 13095 17187
rect 13037 17147 13095 17153
rect 10410 17116 10416 17128
rect 10323 17088 10416 17116
rect 10410 17076 10416 17088
rect 10468 17116 10474 17128
rect 11790 17116 11796 17128
rect 10468 17088 11796 17116
rect 10468 17076 10474 17088
rect 11790 17076 11796 17088
rect 11848 17116 11854 17128
rect 13052 17116 13080 17147
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 13228 17156 13273 17184
rect 13228 17144 13234 17156
rect 13354 17144 13360 17196
rect 13412 17193 13418 17196
rect 13412 17187 13451 17193
rect 13439 17153 13451 17187
rect 13412 17147 13451 17153
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 13998 17184 14004 17196
rect 13587 17156 14004 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 13412 17144 13418 17147
rect 13998 17144 14004 17156
rect 14056 17144 14062 17196
rect 20530 17184 20536 17196
rect 20491 17156 20536 17184
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 20990 17184 20996 17196
rect 20763 17156 20996 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 21726 17144 21732 17196
rect 21784 17184 21790 17196
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21784 17156 21833 17184
rect 21784 17144 21790 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 21910 17144 21916 17196
rect 21968 17184 21974 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21968 17156 22017 17184
rect 21968 17144 21974 17156
rect 22005 17153 22017 17156
rect 22051 17184 22063 17187
rect 22465 17187 22523 17193
rect 22465 17184 22477 17187
rect 22051 17156 22477 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 22465 17153 22477 17156
rect 22511 17153 22523 17187
rect 22646 17184 22652 17196
rect 22607 17156 22652 17184
rect 22465 17147 22523 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 23753 17187 23811 17193
rect 23753 17153 23765 17187
rect 23799 17184 23811 17187
rect 24596 17184 24624 17292
rect 26602 17280 26608 17292
rect 26660 17280 26666 17332
rect 27065 17323 27123 17329
rect 27065 17289 27077 17323
rect 27111 17320 27123 17323
rect 27246 17320 27252 17332
rect 27111 17292 27252 17320
rect 27111 17289 27123 17292
rect 27065 17283 27123 17289
rect 27246 17280 27252 17292
rect 27304 17280 27310 17332
rect 34011 17323 34069 17329
rect 34011 17289 34023 17323
rect 34057 17320 34069 17323
rect 35250 17320 35256 17332
rect 34057 17292 35256 17320
rect 34057 17289 34069 17292
rect 34011 17283 34069 17289
rect 35250 17280 35256 17292
rect 35308 17320 35314 17332
rect 36262 17320 36268 17332
rect 35308 17292 36268 17320
rect 35308 17280 35314 17292
rect 36262 17280 36268 17292
rect 36320 17320 36326 17332
rect 37182 17320 37188 17332
rect 36320 17292 37188 17320
rect 36320 17280 36326 17292
rect 37182 17280 37188 17292
rect 37240 17280 37246 17332
rect 39022 17320 39028 17332
rect 38983 17292 39028 17320
rect 39022 17280 39028 17292
rect 39080 17280 39086 17332
rect 39040 17252 39068 17280
rect 39577 17255 39635 17261
rect 39577 17252 39589 17255
rect 24688 17224 31754 17252
rect 39040 17224 39589 17252
rect 24688 17193 24716 17224
rect 23799 17156 24624 17184
rect 24673 17187 24731 17193
rect 23799 17153 23811 17156
rect 23753 17147 23811 17153
rect 24673 17153 24685 17187
rect 24719 17153 24731 17187
rect 24673 17147 24731 17153
rect 24949 17187 25007 17193
rect 24949 17153 24961 17187
rect 24995 17184 25007 17187
rect 25314 17184 25320 17196
rect 24995 17156 25320 17184
rect 24995 17153 25007 17156
rect 24949 17147 25007 17153
rect 25314 17144 25320 17156
rect 25372 17144 25378 17196
rect 31726 17184 31754 17224
rect 39577 17221 39589 17224
rect 39623 17221 39635 17255
rect 39577 17215 39635 17221
rect 35894 17184 35900 17196
rect 31726 17156 35900 17184
rect 35894 17144 35900 17156
rect 35952 17144 35958 17196
rect 36722 17144 36728 17196
rect 36780 17184 36786 17196
rect 37553 17187 37611 17193
rect 37553 17184 37565 17187
rect 36780 17156 37565 17184
rect 36780 17144 36786 17156
rect 37553 17153 37565 17156
rect 37599 17184 37611 17187
rect 38562 17184 38568 17196
rect 37599 17156 38568 17184
rect 37599 17153 37611 17156
rect 37553 17147 37611 17153
rect 38562 17144 38568 17156
rect 38620 17144 38626 17196
rect 19702 17116 19708 17128
rect 11848 17088 13124 17116
rect 11848 17076 11854 17088
rect 10778 17048 10784 17060
rect 10152 17020 10784 17048
rect 10778 17008 10784 17020
rect 10836 17008 10842 17060
rect 13096 17048 13124 17088
rect 13372 17088 19708 17116
rect 13372 17048 13400 17088
rect 19702 17076 19708 17088
rect 19760 17076 19766 17128
rect 20548 17116 20576 17144
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 20548 17088 21189 17116
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 24394 17116 24400 17128
rect 24075 17088 24400 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 13096 17020 13400 17048
rect 19242 17008 19248 17060
rect 19300 17048 19306 17060
rect 19300 17020 19932 17048
rect 19300 17008 19306 17020
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 6638 16980 6644 16992
rect 6052 16952 6644 16980
rect 6052 16940 6058 16952
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 10505 16983 10563 16989
rect 10505 16980 10517 16983
rect 9456 16952 10517 16980
rect 9456 16940 9462 16952
rect 10505 16949 10517 16952
rect 10551 16949 10563 16983
rect 10505 16943 10563 16949
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 13630 16980 13636 16992
rect 12483 16952 13636 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 18141 16983 18199 16989
rect 18141 16949 18153 16983
rect 18187 16980 18199 16983
rect 18230 16980 18236 16992
rect 18187 16952 18236 16980
rect 18187 16949 18199 16952
rect 18141 16943 18199 16949
rect 18230 16940 18236 16952
rect 18288 16980 18294 16992
rect 18782 16980 18788 16992
rect 18288 16952 18788 16980
rect 18288 16940 18294 16952
rect 18782 16940 18788 16952
rect 18840 16940 18846 16992
rect 19518 16980 19524 16992
rect 19479 16952 19524 16980
rect 19518 16940 19524 16952
rect 19576 16940 19582 16992
rect 19904 16980 19932 17020
rect 19978 17008 19984 17060
rect 20036 17048 20042 17060
rect 21910 17048 21916 17060
rect 20036 17020 21916 17048
rect 20036 17008 20042 17020
rect 21910 17008 21916 17020
rect 21968 17008 21974 17060
rect 22649 17051 22707 17057
rect 22649 17017 22661 17051
rect 22695 17048 22707 17051
rect 24044 17048 24072 17079
rect 24394 17076 24400 17088
rect 24452 17076 24458 17128
rect 24765 17119 24823 17125
rect 24765 17085 24777 17119
rect 24811 17085 24823 17119
rect 24765 17079 24823 17085
rect 22695 17020 24072 17048
rect 22695 17017 22707 17020
rect 22649 17011 22707 17017
rect 24118 17008 24124 17060
rect 24176 17048 24182 17060
rect 24780 17048 24808 17079
rect 25222 17076 25228 17128
rect 25280 17116 25286 17128
rect 25593 17119 25651 17125
rect 25593 17116 25605 17119
rect 25280 17088 25605 17116
rect 25280 17076 25286 17088
rect 25593 17085 25605 17088
rect 25639 17116 25651 17119
rect 25866 17116 25872 17128
rect 25639 17088 25872 17116
rect 25639 17085 25651 17088
rect 25593 17079 25651 17085
rect 25866 17076 25872 17088
rect 25924 17116 25930 17128
rect 33778 17116 33784 17128
rect 25924 17088 31754 17116
rect 33739 17088 33784 17116
rect 25924 17076 25930 17088
rect 24176 17020 24808 17048
rect 24176 17008 24182 17020
rect 27154 17008 27160 17060
rect 27212 17048 27218 17060
rect 29546 17048 29552 17060
rect 27212 17020 29552 17048
rect 27212 17008 27218 17020
rect 29546 17008 29552 17020
rect 29604 17008 29610 17060
rect 31726 17048 31754 17088
rect 33778 17076 33784 17088
rect 33836 17076 33842 17128
rect 34606 17076 34612 17128
rect 34664 17116 34670 17128
rect 34974 17116 34980 17128
rect 34664 17088 34980 17116
rect 34664 17076 34670 17088
rect 34974 17076 34980 17088
rect 35032 17116 35038 17128
rect 35069 17119 35127 17125
rect 35069 17116 35081 17119
rect 35032 17088 35081 17116
rect 35032 17076 35038 17088
rect 35069 17085 35081 17088
rect 35115 17085 35127 17119
rect 35069 17079 35127 17085
rect 35345 17119 35403 17125
rect 35345 17085 35357 17119
rect 35391 17116 35403 17119
rect 36078 17116 36084 17128
rect 35391 17088 36084 17116
rect 35391 17085 35403 17088
rect 35345 17079 35403 17085
rect 36078 17076 36084 17088
rect 36136 17076 36142 17128
rect 36814 17076 36820 17128
rect 36872 17116 36878 17128
rect 37277 17119 37335 17125
rect 37277 17116 37289 17119
rect 36872 17088 37289 17116
rect 36872 17076 36878 17088
rect 37277 17085 37289 17088
rect 37323 17085 37335 17119
rect 37277 17079 37335 17085
rect 38194 17076 38200 17128
rect 38252 17116 38258 17128
rect 40494 17116 40500 17128
rect 38252 17088 40500 17116
rect 38252 17076 38258 17088
rect 40494 17076 40500 17088
rect 40552 17076 40558 17128
rect 58158 17048 58164 17060
rect 31726 17020 32904 17048
rect 58119 17020 58164 17048
rect 32876 16992 32904 17020
rect 58158 17008 58164 17020
rect 58216 17008 58222 17060
rect 24762 16980 24768 16992
rect 19904 16952 24768 16980
rect 24762 16940 24768 16952
rect 24820 16940 24826 16992
rect 24946 16980 24952 16992
rect 24907 16952 24952 16980
rect 24946 16940 24952 16952
rect 25004 16940 25010 16992
rect 32858 16940 32864 16992
rect 32916 16980 32922 16992
rect 35526 16980 35532 16992
rect 32916 16952 35532 16980
rect 32916 16940 32922 16952
rect 35526 16940 35532 16952
rect 35584 16940 35590 16992
rect 37734 16940 37740 16992
rect 37792 16980 37798 16992
rect 39758 16980 39764 16992
rect 37792 16952 39764 16980
rect 37792 16940 37798 16952
rect 39758 16940 39764 16952
rect 39816 16940 39822 16992
rect 40034 16940 40040 16992
rect 40092 16980 40098 16992
rect 40865 16983 40923 16989
rect 40865 16980 40877 16983
rect 40092 16952 40877 16980
rect 40092 16940 40098 16952
rect 40865 16949 40877 16952
rect 40911 16949 40923 16983
rect 40865 16943 40923 16949
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 5258 16776 5264 16788
rect 5219 16748 5264 16776
rect 5258 16736 5264 16748
rect 5316 16736 5322 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 12710 16776 12716 16788
rect 9732 16748 12434 16776
rect 12671 16748 12716 16776
rect 9732 16736 9738 16748
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 11885 16711 11943 16717
rect 11885 16708 11897 16711
rect 8352 16680 11897 16708
rect 8352 16668 8358 16680
rect 11885 16677 11897 16680
rect 11931 16677 11943 16711
rect 12406 16708 12434 16748
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 13446 16736 13452 16788
rect 13504 16776 13510 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 13504 16748 13553 16776
rect 13504 16736 13510 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 13541 16739 13599 16745
rect 14016 16748 16405 16776
rect 14016 16708 14044 16748
rect 16393 16745 16405 16748
rect 16439 16776 16451 16779
rect 17310 16776 17316 16788
rect 16439 16748 17316 16776
rect 16439 16745 16451 16748
rect 16393 16739 16451 16745
rect 17310 16736 17316 16748
rect 17368 16736 17374 16788
rect 17494 16776 17500 16788
rect 17455 16748 17500 16776
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 18233 16779 18291 16785
rect 18233 16745 18245 16779
rect 18279 16776 18291 16779
rect 18690 16776 18696 16788
rect 18279 16748 18696 16776
rect 18279 16745 18291 16748
rect 18233 16739 18291 16745
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19702 16776 19708 16788
rect 19484 16748 19708 16776
rect 19484 16736 19490 16748
rect 19702 16736 19708 16748
rect 19760 16736 19766 16788
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 20349 16779 20407 16785
rect 20349 16776 20361 16779
rect 20128 16748 20361 16776
rect 20128 16736 20134 16748
rect 20349 16745 20361 16748
rect 20395 16745 20407 16779
rect 21910 16776 21916 16788
rect 21871 16748 21916 16776
rect 20349 16739 20407 16745
rect 21910 16736 21916 16748
rect 21968 16736 21974 16788
rect 22649 16779 22707 16785
rect 22649 16745 22661 16779
rect 22695 16776 22707 16779
rect 24578 16776 24584 16788
rect 22695 16748 24440 16776
rect 24539 16748 24584 16776
rect 22695 16745 22707 16748
rect 22649 16739 22707 16745
rect 12406 16680 14044 16708
rect 11885 16671 11943 16677
rect 14090 16668 14096 16720
rect 14148 16708 14154 16720
rect 24412 16708 24440 16748
rect 24578 16736 24584 16748
rect 24636 16736 24642 16788
rect 25314 16776 25320 16788
rect 25275 16748 25320 16776
rect 25314 16736 25320 16748
rect 25372 16736 25378 16788
rect 26234 16736 26240 16788
rect 26292 16776 26298 16788
rect 26697 16779 26755 16785
rect 26697 16776 26709 16779
rect 26292 16748 26709 16776
rect 26292 16736 26298 16748
rect 26697 16745 26709 16748
rect 26743 16776 26755 16779
rect 27430 16776 27436 16788
rect 26743 16748 27436 16776
rect 26743 16745 26755 16748
rect 26697 16739 26755 16745
rect 27430 16736 27436 16748
rect 27488 16736 27494 16788
rect 27706 16736 27712 16788
rect 27764 16776 27770 16788
rect 34054 16776 34060 16788
rect 27764 16748 34060 16776
rect 27764 16736 27770 16748
rect 34054 16736 34060 16748
rect 34112 16736 34118 16788
rect 35894 16776 35900 16788
rect 35807 16748 35900 16776
rect 35894 16736 35900 16748
rect 35952 16776 35958 16788
rect 36354 16776 36360 16788
rect 35952 16748 36360 16776
rect 35952 16736 35958 16748
rect 36354 16736 36360 16748
rect 36412 16736 36418 16788
rect 37292 16748 39344 16776
rect 27798 16708 27804 16720
rect 14148 16680 23336 16708
rect 24412 16680 27660 16708
rect 27759 16680 27804 16708
rect 14148 16668 14154 16680
rect 10778 16640 10784 16652
rect 10244 16612 10784 16640
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16572 4491 16575
rect 5350 16572 5356 16584
rect 4479 16544 5356 16572
rect 4479 16541 4491 16544
rect 4433 16535 4491 16541
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 9950 16572 9956 16584
rect 9911 16544 9956 16572
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10134 16581 10140 16584
rect 10101 16575 10140 16581
rect 10101 16541 10113 16575
rect 10101 16535 10140 16541
rect 10134 16532 10140 16535
rect 10192 16532 10198 16584
rect 10244 16581 10272 16612
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 14108 16640 14136 16668
rect 15286 16640 15292 16652
rect 12912 16612 14136 16640
rect 15247 16612 15292 16640
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 10410 16532 10416 16584
rect 10468 16581 10474 16584
rect 10468 16572 10476 16581
rect 11238 16572 11244 16584
rect 10468 16544 10513 16572
rect 11199 16544 11244 16572
rect 10468 16535 10476 16544
rect 10468 16532 10474 16535
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 11790 16581 11796 16584
rect 11334 16575 11392 16581
rect 11334 16541 11346 16575
rect 11380 16541 11392 16575
rect 11334 16535 11392 16541
rect 11747 16575 11796 16581
rect 11747 16541 11759 16575
rect 11793 16541 11796 16575
rect 11747 16535 11796 16541
rect 10318 16504 10324 16516
rect 10279 16476 10324 16504
rect 10318 16464 10324 16476
rect 10376 16464 10382 16516
rect 10962 16464 10968 16516
rect 11020 16504 11026 16516
rect 11348 16504 11376 16535
rect 11790 16532 11796 16535
rect 11848 16532 11854 16584
rect 12158 16532 12164 16584
rect 12216 16572 12222 16584
rect 12912 16581 12940 16612
rect 13372 16581 13400 16612
rect 15286 16600 15292 16612
rect 15344 16640 15350 16652
rect 15930 16640 15936 16652
rect 15344 16612 15936 16640
rect 15344 16600 15350 16612
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 16942 16640 16948 16652
rect 16903 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 21361 16643 21419 16649
rect 21361 16640 21373 16643
rect 18064 16612 21373 16640
rect 12713 16575 12771 16581
rect 12713 16572 12725 16575
rect 12216 16544 12725 16572
rect 12216 16532 12222 16544
rect 12713 16541 12725 16544
rect 12759 16541 12771 16575
rect 12713 16535 12771 16541
rect 12897 16575 12955 16581
rect 12897 16541 12909 16575
rect 12943 16541 12955 16575
rect 12897 16535 12955 16541
rect 13357 16575 13415 16581
rect 13357 16541 13369 16575
rect 13403 16541 13415 16575
rect 13357 16535 13415 16541
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16572 13599 16575
rect 13630 16572 13636 16584
rect 13587 16544 13636 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 11020 16476 11376 16504
rect 11517 16507 11575 16513
rect 11020 16464 11026 16476
rect 11517 16473 11529 16507
rect 11563 16473 11575 16507
rect 11517 16467 11575 16473
rect 3878 16396 3884 16448
rect 3936 16436 3942 16448
rect 4249 16439 4307 16445
rect 4249 16436 4261 16439
rect 3936 16408 4261 16436
rect 3936 16396 3942 16408
rect 4249 16405 4261 16408
rect 4295 16405 4307 16439
rect 10594 16436 10600 16448
rect 10555 16408 10600 16436
rect 4249 16399 4307 16405
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 11532 16436 11560 16467
rect 11606 16464 11612 16516
rect 11664 16504 11670 16516
rect 11664 16476 11709 16504
rect 11664 16464 11670 16476
rect 11882 16464 11888 16516
rect 11940 16504 11946 16516
rect 12912 16504 12940 16535
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 14737 16575 14795 16581
rect 14737 16541 14749 16575
rect 14783 16572 14795 16575
rect 15194 16572 15200 16584
rect 14783 16544 15200 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 15194 16532 15200 16544
rect 15252 16532 15258 16584
rect 17494 16532 17500 16584
rect 17552 16572 17558 16584
rect 18064 16581 18092 16612
rect 21361 16609 21373 16612
rect 21407 16640 21419 16643
rect 23198 16640 23204 16652
rect 21407 16612 22508 16640
rect 23159 16612 23204 16640
rect 21407 16609 21419 16612
rect 21361 16603 21419 16609
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17552 16544 18061 16572
rect 17552 16532 17558 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18230 16572 18236 16584
rect 18191 16544 18236 16572
rect 18049 16535 18107 16541
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 19518 16572 19524 16584
rect 18340 16544 19524 16572
rect 14550 16504 14556 16516
rect 11940 16476 12940 16504
rect 14511 16476 14556 16504
rect 11940 16464 11946 16476
rect 14550 16464 14556 16476
rect 14608 16464 14614 16516
rect 12710 16436 12716 16448
rect 10836 16408 12716 16436
rect 10836 16396 10842 16408
rect 12710 16396 12716 16408
rect 12768 16396 12774 16448
rect 13722 16396 13728 16448
rect 13780 16436 13786 16448
rect 18340 16436 18368 16544
rect 19518 16532 19524 16544
rect 19576 16532 19582 16584
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16572 19855 16575
rect 20070 16572 20076 16584
rect 19843 16544 20076 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 20070 16532 20076 16544
rect 20128 16532 20134 16584
rect 20162 16532 20168 16584
rect 20220 16572 20226 16584
rect 22480 16581 22508 16612
rect 23198 16600 23204 16612
rect 23256 16600 23262 16652
rect 23308 16640 23336 16680
rect 23753 16643 23811 16649
rect 23753 16640 23765 16643
rect 23308 16612 23765 16640
rect 20349 16575 20407 16581
rect 20349 16572 20361 16575
rect 20220 16544 20361 16572
rect 20220 16532 20226 16544
rect 20349 16541 20361 16544
rect 20395 16541 20407 16575
rect 20349 16535 20407 16541
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22646 16572 22652 16584
rect 22607 16544 22652 16572
rect 22465 16535 22523 16541
rect 13780 16408 18368 16436
rect 13780 16396 13786 16408
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 20548 16436 20576 16535
rect 22646 16532 22652 16544
rect 22704 16572 22710 16584
rect 23308 16581 23336 16612
rect 23753 16609 23765 16612
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 24486 16600 24492 16652
rect 24544 16640 24550 16652
rect 24544 16612 24624 16640
rect 24544 16600 24550 16612
rect 24596 16581 24624 16612
rect 24762 16600 24768 16652
rect 24820 16640 24826 16652
rect 26145 16643 26203 16649
rect 26145 16640 26157 16643
rect 24820 16612 26157 16640
rect 24820 16600 24826 16612
rect 26145 16609 26157 16612
rect 26191 16640 26203 16643
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 26191 16612 27077 16640
rect 26191 16609 26203 16612
rect 26145 16603 26203 16609
rect 27065 16609 27077 16612
rect 27111 16609 27123 16643
rect 27632 16640 27660 16680
rect 27798 16668 27804 16680
rect 27856 16668 27862 16720
rect 33778 16708 33784 16720
rect 28966 16680 33784 16708
rect 28966 16640 28994 16680
rect 29546 16640 29552 16652
rect 27632 16612 28994 16640
rect 29507 16612 29552 16640
rect 27065 16603 27123 16609
rect 23109 16575 23167 16581
rect 23109 16572 23121 16575
rect 22704 16544 23121 16572
rect 22704 16532 22710 16544
rect 23109 16541 23121 16544
rect 23155 16541 23167 16575
rect 23109 16535 23167 16541
rect 23293 16575 23351 16581
rect 23293 16541 23305 16575
rect 23339 16541 23351 16575
rect 23293 16535 23351 16541
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24670 16532 24676 16584
rect 24728 16572 24734 16584
rect 24857 16575 24915 16581
rect 24728 16544 24773 16572
rect 24728 16532 24734 16544
rect 24857 16541 24869 16575
rect 24903 16572 24915 16575
rect 25038 16572 25044 16584
rect 24903 16544 25044 16572
rect 24903 16541 24915 16544
rect 24857 16535 24915 16541
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 26602 16532 26608 16584
rect 26660 16572 26666 16584
rect 26881 16575 26939 16581
rect 26881 16572 26893 16575
rect 26660 16544 26893 16572
rect 26660 16532 26666 16544
rect 26881 16541 26893 16544
rect 26927 16541 26939 16575
rect 27080 16572 27108 16603
rect 29546 16600 29552 16612
rect 29604 16640 29610 16652
rect 29914 16640 29920 16652
rect 29604 16612 29920 16640
rect 29604 16600 29610 16612
rect 29914 16600 29920 16612
rect 29972 16640 29978 16652
rect 30377 16643 30435 16649
rect 29972 16612 30236 16640
rect 29972 16600 29978 16612
rect 27706 16572 27712 16584
rect 27080 16544 27712 16572
rect 26881 16535 26939 16541
rect 27706 16532 27712 16544
rect 27764 16532 27770 16584
rect 30208 16581 30236 16612
rect 30377 16609 30389 16643
rect 30423 16640 30435 16643
rect 32033 16643 32091 16649
rect 32033 16640 32045 16643
rect 30423 16612 32045 16640
rect 30423 16609 30435 16612
rect 30377 16603 30435 16609
rect 32033 16609 32045 16612
rect 32079 16640 32091 16643
rect 32582 16640 32588 16652
rect 32079 16612 32588 16640
rect 32079 16609 32091 16612
rect 32033 16603 32091 16609
rect 32582 16600 32588 16612
rect 32640 16600 32646 16652
rect 32858 16640 32864 16652
rect 32819 16612 32864 16640
rect 32858 16600 32864 16612
rect 32916 16600 32922 16652
rect 33336 16649 33364 16680
rect 33778 16668 33784 16680
rect 33836 16668 33842 16720
rect 33321 16643 33379 16649
rect 33321 16609 33333 16643
rect 33367 16609 33379 16643
rect 33321 16603 33379 16609
rect 33597 16643 33655 16649
rect 33597 16609 33609 16643
rect 33643 16640 33655 16643
rect 34698 16640 34704 16652
rect 33643 16612 33824 16640
rect 33643 16609 33655 16612
rect 33597 16603 33655 16609
rect 30193 16575 30251 16581
rect 30193 16541 30205 16575
rect 30239 16541 30251 16575
rect 30193 16535 30251 16541
rect 20622 16464 20628 16516
rect 20680 16504 20686 16516
rect 27617 16507 27675 16513
rect 27617 16504 27629 16507
rect 20680 16476 27629 16504
rect 20680 16464 20686 16476
rect 27617 16473 27629 16476
rect 27663 16473 27675 16507
rect 33796 16504 33824 16612
rect 34072 16612 34704 16640
rect 34072 16504 34100 16612
rect 34698 16600 34704 16612
rect 34756 16600 34762 16652
rect 37292 16649 37320 16748
rect 37918 16708 37924 16720
rect 37879 16680 37924 16708
rect 37918 16668 37924 16680
rect 37976 16668 37982 16720
rect 39316 16649 39344 16748
rect 37277 16643 37335 16649
rect 37277 16609 37289 16643
rect 37323 16609 37335 16643
rect 37277 16603 37335 16609
rect 39301 16643 39359 16649
rect 39301 16609 39313 16643
rect 39347 16640 39359 16643
rect 40034 16640 40040 16652
rect 39347 16612 40040 16640
rect 39347 16609 39359 16612
rect 39301 16603 39359 16609
rect 40034 16600 40040 16612
rect 40092 16600 40098 16652
rect 34793 16575 34851 16581
rect 34793 16572 34805 16575
rect 33796 16476 34100 16504
rect 34716 16544 34805 16572
rect 27617 16467 27675 16473
rect 34716 16448 34744 16544
rect 34793 16541 34805 16544
rect 34839 16541 34851 16575
rect 34974 16572 34980 16584
rect 34935 16544 34980 16572
rect 34793 16535 34851 16541
rect 34974 16532 34980 16544
rect 35032 16532 35038 16584
rect 35069 16575 35127 16581
rect 35069 16541 35081 16575
rect 35115 16541 35127 16575
rect 35069 16535 35127 16541
rect 35161 16575 35219 16581
rect 35161 16541 35173 16575
rect 35207 16572 35219 16575
rect 35526 16572 35532 16584
rect 35207 16544 35532 16572
rect 35207 16541 35219 16544
rect 35161 16535 35219 16541
rect 35084 16504 35112 16535
rect 35526 16532 35532 16544
rect 35584 16532 35590 16584
rect 35437 16507 35495 16513
rect 35084 16476 35204 16504
rect 20806 16436 20812 16448
rect 19576 16408 20812 16436
rect 19576 16396 19582 16408
rect 20806 16396 20812 16408
rect 20864 16436 20870 16448
rect 20990 16436 20996 16448
rect 20864 16408 20996 16436
rect 20864 16396 20870 16408
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 24302 16396 24308 16448
rect 24360 16436 24366 16448
rect 24397 16439 24455 16445
rect 24397 16436 24409 16439
rect 24360 16408 24409 16436
rect 24360 16396 24366 16408
rect 24397 16405 24409 16408
rect 24443 16405 24455 16439
rect 24397 16399 24455 16405
rect 34698 16396 34704 16448
rect 34756 16396 34762 16448
rect 35176 16436 35204 16476
rect 35437 16473 35449 16507
rect 35483 16504 35495 16507
rect 37010 16507 37068 16513
rect 37010 16504 37022 16507
rect 35483 16476 37022 16504
rect 35483 16473 35495 16476
rect 35437 16467 35495 16473
rect 37010 16473 37022 16476
rect 37056 16473 37068 16507
rect 37010 16467 37068 16473
rect 38654 16464 38660 16516
rect 38712 16504 38718 16516
rect 39034 16507 39092 16513
rect 39034 16504 39046 16507
rect 38712 16476 39046 16504
rect 38712 16464 38718 16476
rect 39034 16473 39046 16476
rect 39080 16473 39092 16507
rect 39034 16467 39092 16473
rect 37090 16436 37096 16448
rect 35176 16408 37096 16436
rect 37090 16396 37096 16408
rect 37148 16396 37154 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 5442 16232 5448 16244
rect 3160 16204 5448 16232
rect 3160 16173 3188 16204
rect 5442 16192 5448 16204
rect 5500 16232 5506 16244
rect 6914 16232 6920 16244
rect 5500 16204 6920 16232
rect 5500 16192 5506 16204
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 10505 16235 10563 16241
rect 10505 16201 10517 16235
rect 10551 16232 10563 16235
rect 10870 16232 10876 16244
rect 10551 16204 10876 16232
rect 10551 16201 10563 16204
rect 10505 16195 10563 16201
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11974 16192 11980 16244
rect 12032 16232 12038 16244
rect 15378 16232 15384 16244
rect 12032 16204 15384 16232
rect 12032 16192 12038 16204
rect 15378 16192 15384 16204
rect 15436 16192 15442 16244
rect 17218 16232 17224 16244
rect 15488 16204 17224 16232
rect 3145 16167 3203 16173
rect 3145 16133 3157 16167
rect 3191 16133 3203 16167
rect 3145 16127 3203 16133
rect 10318 16124 10324 16176
rect 10376 16164 10382 16176
rect 11790 16164 11796 16176
rect 10376 16136 11796 16164
rect 10376 16124 10382 16136
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 12161 16167 12219 16173
rect 12161 16133 12173 16167
rect 12207 16164 12219 16167
rect 12207 16136 13584 16164
rect 12207 16133 12219 16136
rect 12161 16127 12219 16133
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2498 16096 2504 16108
rect 2455 16068 2504 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2498 16056 2504 16068
rect 2556 16056 2562 16108
rect 7650 16096 7656 16108
rect 7611 16068 7656 16096
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16096 7803 16099
rect 9398 16096 9404 16108
rect 7791 16068 9404 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 10042 16056 10048 16108
rect 10100 16096 10106 16108
rect 10226 16096 10232 16108
rect 10100 16068 10232 16096
rect 10100 16056 10106 16068
rect 10226 16056 10232 16068
rect 10284 16096 10290 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 10284 16068 10425 16096
rect 10284 16056 10290 16068
rect 10413 16065 10425 16068
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 10597 16099 10655 16105
rect 10597 16065 10609 16099
rect 10643 16096 10655 16099
rect 11330 16096 11336 16108
rect 10643 16068 11336 16096
rect 10643 16065 10655 16068
rect 10597 16059 10655 16065
rect 11330 16056 11336 16068
rect 11388 16096 11394 16108
rect 12069 16099 12127 16105
rect 12069 16096 12081 16099
rect 11388 16068 12081 16096
rect 11388 16056 11394 16068
rect 12069 16065 12081 16068
rect 12115 16065 12127 16099
rect 12069 16059 12127 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 12434 16096 12440 16108
rect 12299 16068 12440 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 3970 15988 3976 16040
rect 4028 16028 4034 16040
rect 11054 16028 11060 16040
rect 4028 16000 11060 16028
rect 4028 15988 4034 16000
rect 11054 15988 11060 16000
rect 11112 16028 11118 16040
rect 12084 16028 12112 16059
rect 12434 16056 12440 16068
rect 12492 16096 12498 16108
rect 12492 16068 12664 16096
rect 12492 16056 12498 16068
rect 12158 16028 12164 16040
rect 11112 16000 12020 16028
rect 12084 16000 12164 16028
rect 11112 15988 11118 16000
rect 4982 15920 4988 15972
rect 5040 15960 5046 15972
rect 5040 15932 7604 15960
rect 5040 15920 5046 15932
rect 2222 15892 2228 15904
rect 2183 15864 2228 15892
rect 2222 15852 2228 15864
rect 2280 15852 2286 15904
rect 4614 15892 4620 15904
rect 4575 15864 4620 15892
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 6638 15852 6644 15904
rect 6696 15892 6702 15904
rect 7576 15901 7604 15932
rect 7377 15895 7435 15901
rect 7377 15892 7389 15895
rect 6696 15864 7389 15892
rect 6696 15852 6702 15864
rect 7377 15861 7389 15864
rect 7423 15861 7435 15895
rect 7377 15855 7435 15861
rect 7561 15895 7619 15901
rect 7561 15861 7573 15895
rect 7607 15861 7619 15895
rect 7561 15855 7619 15861
rect 9953 15895 10011 15901
rect 9953 15861 9965 15895
rect 9999 15892 10011 15895
rect 10042 15892 10048 15904
rect 9999 15864 10048 15892
rect 9999 15861 10011 15864
rect 9953 15855 10011 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 11609 15895 11667 15901
rect 11609 15861 11621 15895
rect 11655 15892 11667 15895
rect 11698 15892 11704 15904
rect 11655 15864 11704 15892
rect 11655 15861 11667 15864
rect 11609 15855 11667 15861
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 11992 15892 12020 16000
rect 12158 15988 12164 16000
rect 12216 15988 12222 16040
rect 12636 16028 12664 16068
rect 12710 16056 12716 16108
rect 12768 16096 12774 16108
rect 13262 16096 13268 16108
rect 12768 16068 13268 16096
rect 12768 16056 12774 16068
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 13556 16105 13584 16136
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16096 13599 16099
rect 14550 16096 14556 16108
rect 13587 16068 14556 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 14645 16099 14703 16105
rect 14645 16065 14657 16099
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16065 14795 16099
rect 14737 16059 14795 16065
rect 13722 16028 13728 16040
rect 12636 16000 13728 16028
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 14182 15960 14188 15972
rect 12406 15932 14188 15960
rect 12406 15892 12434 15932
rect 14182 15920 14188 15932
rect 14240 15960 14246 15972
rect 14660 15960 14688 16059
rect 14752 16028 14780 16059
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 15488 16105 15516 16204
rect 16758 16164 16764 16176
rect 15580 16136 16764 16164
rect 15013 16099 15071 16105
rect 14884 16068 14929 16096
rect 14884 16056 14890 16068
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15059 16068 15485 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15473 16065 15485 16068
rect 15519 16065 15531 16099
rect 15473 16059 15531 16065
rect 15580 16028 15608 16136
rect 15764 16105 15792 16136
rect 16758 16124 16764 16136
rect 16816 16124 16822 16176
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 15841 16099 15899 16105
rect 15841 16065 15853 16099
rect 15887 16096 15899 16099
rect 15930 16096 15936 16108
rect 15887 16068 15936 16096
rect 15887 16065 15899 16068
rect 15841 16059 15899 16065
rect 14752 16000 15608 16028
rect 15672 16028 15700 16059
rect 15930 16056 15936 16068
rect 15988 16056 15994 16108
rect 16666 16028 16672 16040
rect 15672 16000 16672 16028
rect 16666 15988 16672 16000
rect 16724 15988 16730 16040
rect 16776 16028 16804 16124
rect 16960 16105 16988 16204
rect 17218 16192 17224 16204
rect 17276 16192 17282 16244
rect 19337 16235 19395 16241
rect 19337 16201 19349 16235
rect 19383 16232 19395 16235
rect 20622 16232 20628 16244
rect 19383 16204 20628 16232
rect 19383 16201 19395 16204
rect 19337 16195 19395 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20806 16232 20812 16244
rect 20767 16204 20812 16232
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 21726 16192 21732 16244
rect 21784 16232 21790 16244
rect 21821 16235 21879 16241
rect 21821 16232 21833 16235
rect 21784 16204 21833 16232
rect 21784 16192 21790 16204
rect 21821 16201 21833 16204
rect 21867 16201 21879 16235
rect 21821 16195 21879 16201
rect 22646 16192 22652 16244
rect 22704 16232 22710 16244
rect 22741 16235 22799 16241
rect 22741 16232 22753 16235
rect 22704 16204 22753 16232
rect 22704 16192 22710 16204
rect 22741 16201 22753 16204
rect 22787 16201 22799 16235
rect 22741 16195 22799 16201
rect 24486 16192 24492 16244
rect 24544 16232 24550 16244
rect 24544 16204 34376 16232
rect 24544 16192 24550 16204
rect 18417 16167 18475 16173
rect 18417 16164 18429 16167
rect 17144 16136 18429 16164
rect 17144 16105 17172 16136
rect 18417 16133 18429 16136
rect 18463 16133 18475 16167
rect 18417 16127 18475 16133
rect 31573 16167 31631 16173
rect 31573 16133 31585 16167
rect 31619 16164 31631 16167
rect 34348 16164 34376 16204
rect 34974 16192 34980 16244
rect 35032 16232 35038 16244
rect 35161 16235 35219 16241
rect 35161 16232 35173 16235
rect 35032 16204 35173 16232
rect 35032 16192 35038 16204
rect 35161 16201 35173 16204
rect 35207 16201 35219 16235
rect 36906 16232 36912 16244
rect 35161 16195 35219 16201
rect 35268 16204 36912 16232
rect 35268 16164 35296 16204
rect 36906 16192 36912 16204
rect 36964 16192 36970 16244
rect 37461 16235 37519 16241
rect 37461 16201 37473 16235
rect 37507 16232 37519 16235
rect 37734 16232 37740 16244
rect 37507 16204 37740 16232
rect 37507 16201 37519 16204
rect 37461 16195 37519 16201
rect 37734 16192 37740 16204
rect 37792 16192 37798 16244
rect 38838 16232 38844 16244
rect 38212 16204 38844 16232
rect 31619 16136 32352 16164
rect 34348 16136 35296 16164
rect 35345 16167 35403 16173
rect 31619 16133 31631 16136
rect 31573 16127 31631 16133
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16065 17187 16099
rect 17129 16059 17187 16065
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16065 17279 16099
rect 17221 16059 17279 16065
rect 17236 16028 17264 16059
rect 17310 16056 17316 16108
rect 17368 16096 17374 16108
rect 17368 16068 17413 16096
rect 17368 16056 17374 16068
rect 17770 16056 17776 16108
rect 17828 16096 17834 16108
rect 18049 16099 18107 16105
rect 18049 16096 18061 16099
rect 17828 16068 18061 16096
rect 17828 16056 17834 16068
rect 18049 16065 18061 16068
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 18233 16099 18291 16105
rect 18233 16065 18245 16099
rect 18279 16065 18291 16099
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 18233 16059 18291 16065
rect 16776 16000 17264 16028
rect 18248 16028 18276 16059
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19426 16096 19432 16108
rect 19387 16068 19432 16096
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 26234 16096 26240 16108
rect 26195 16068 26240 16096
rect 26234 16056 26240 16068
rect 26292 16056 26298 16108
rect 27801 16099 27859 16105
rect 27801 16065 27813 16099
rect 27847 16096 27859 16099
rect 27890 16096 27896 16108
rect 27847 16068 27896 16096
rect 27847 16065 27859 16068
rect 27801 16059 27859 16065
rect 27890 16056 27896 16068
rect 27948 16056 27954 16108
rect 30742 16056 30748 16108
rect 30800 16096 30806 16108
rect 31205 16099 31263 16105
rect 31205 16096 31217 16099
rect 30800 16068 31217 16096
rect 30800 16056 30806 16068
rect 31205 16065 31217 16068
rect 31251 16065 31263 16099
rect 31205 16059 31263 16065
rect 31389 16099 31447 16105
rect 31389 16065 31401 16099
rect 31435 16096 31447 16099
rect 32030 16096 32036 16108
rect 31435 16068 32036 16096
rect 31435 16065 31447 16068
rect 31389 16059 31447 16065
rect 32030 16056 32036 16068
rect 32088 16056 32094 16108
rect 32324 16105 32352 16136
rect 35345 16133 35357 16167
rect 35391 16164 35403 16167
rect 35894 16164 35900 16176
rect 35391 16136 35900 16164
rect 35391 16133 35403 16136
rect 35345 16127 35403 16133
rect 35894 16124 35900 16136
rect 35952 16124 35958 16176
rect 36354 16124 36360 16176
rect 36412 16164 36418 16176
rect 36538 16164 36544 16176
rect 36412 16136 36544 16164
rect 36412 16124 36418 16136
rect 36538 16124 36544 16136
rect 36596 16124 36602 16176
rect 38212 16173 38240 16204
rect 38825 16192 38844 16204
rect 38896 16192 38902 16244
rect 39022 16192 39028 16244
rect 39080 16232 39086 16244
rect 39080 16204 39252 16232
rect 39080 16192 39086 16204
rect 38197 16167 38255 16173
rect 38197 16133 38209 16167
rect 38243 16133 38255 16167
rect 38197 16127 38255 16133
rect 32125 16099 32183 16105
rect 32125 16065 32137 16099
rect 32171 16065 32183 16099
rect 32125 16059 32183 16065
rect 32309 16099 32367 16105
rect 32309 16065 32321 16099
rect 32355 16065 32367 16099
rect 32309 16059 32367 16065
rect 32401 16099 32459 16105
rect 32401 16065 32413 16099
rect 32447 16065 32459 16099
rect 32401 16059 32459 16065
rect 32493 16099 32551 16105
rect 32493 16065 32505 16099
rect 32539 16096 32551 16099
rect 32582 16096 32588 16108
rect 32539 16068 32588 16096
rect 32539 16065 32551 16068
rect 32493 16059 32551 16065
rect 19334 16028 19340 16040
rect 18248 16000 19340 16028
rect 19334 15988 19340 16000
rect 19392 15988 19398 16040
rect 25038 16028 25044 16040
rect 24999 16000 25044 16028
rect 25038 15988 25044 16000
rect 25096 15988 25102 16040
rect 27430 15988 27436 16040
rect 27488 16028 27494 16040
rect 27525 16031 27583 16037
rect 27525 16028 27537 16031
rect 27488 16000 27537 16028
rect 27488 15988 27494 16000
rect 27525 15997 27537 16000
rect 27571 15997 27583 16031
rect 27525 15991 27583 15997
rect 30374 15988 30380 16040
rect 30432 16028 30438 16040
rect 32140 16028 32168 16059
rect 30432 16000 32168 16028
rect 30432 15988 30438 16000
rect 14240 15932 14688 15960
rect 14240 15920 14246 15932
rect 15378 15920 15384 15972
rect 15436 15960 15442 15972
rect 20165 15963 20223 15969
rect 20165 15960 20177 15963
rect 15436 15932 20177 15960
rect 15436 15920 15442 15932
rect 20165 15929 20177 15932
rect 20211 15960 20223 15963
rect 20530 15960 20536 15972
rect 20211 15932 20536 15960
rect 20211 15929 20223 15932
rect 20165 15923 20223 15929
rect 20530 15920 20536 15932
rect 20588 15920 20594 15972
rect 31846 15920 31852 15972
rect 31904 15960 31910 15972
rect 32416 15960 32444 16059
rect 32582 16056 32588 16068
rect 32640 16056 32646 16108
rect 34606 16096 34612 16108
rect 34567 16068 34612 16096
rect 34606 16056 34612 16068
rect 34664 16056 34670 16108
rect 35529 16099 35587 16105
rect 35529 16065 35541 16099
rect 35575 16096 35587 16099
rect 36814 16096 36820 16108
rect 35575 16068 36820 16096
rect 35575 16065 35587 16068
rect 35529 16059 35587 16065
rect 36814 16056 36820 16068
rect 36872 16056 36878 16108
rect 37182 16056 37188 16108
rect 37240 16096 37246 16108
rect 37277 16099 37335 16105
rect 37277 16096 37289 16099
rect 37240 16068 37289 16096
rect 37240 16056 37246 16068
rect 37277 16065 37289 16068
rect 37323 16065 37335 16099
rect 37277 16059 37335 16065
rect 34333 16031 34391 16037
rect 34333 15997 34345 16031
rect 34379 16028 34391 16031
rect 34514 16028 34520 16040
rect 34379 16000 34520 16028
rect 34379 15997 34391 16000
rect 34333 15991 34391 15997
rect 34514 15988 34520 16000
rect 34572 15988 34578 16040
rect 38212 16028 38240 16127
rect 38825 16080 38853 16192
rect 39224 16164 39252 16204
rect 39224 16136 39344 16164
rect 38913 16099 38971 16105
rect 38913 16096 38925 16099
rect 38902 16080 38925 16096
rect 38825 16065 38925 16080
rect 38959 16065 38971 16099
rect 38825 16059 38971 16065
rect 39025 16099 39083 16105
rect 39025 16065 39037 16099
rect 39071 16065 39083 16099
rect 39025 16059 39083 16065
rect 39117 16099 39175 16105
rect 39117 16065 39129 16099
rect 39163 16096 39175 16099
rect 39206 16096 39212 16108
rect 39163 16068 39212 16096
rect 39163 16065 39175 16068
rect 39117 16059 39175 16065
rect 38825 16052 38930 16059
rect 37246 16000 38240 16028
rect 31904 15932 32444 15960
rect 31904 15920 31910 15932
rect 14366 15892 14372 15904
rect 11992 15864 12434 15892
rect 14327 15864 14372 15892
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 16114 15892 16120 15904
rect 16075 15864 16120 15892
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 17589 15895 17647 15901
rect 17589 15861 17601 15895
rect 17635 15892 17647 15895
rect 18046 15892 18052 15904
rect 17635 15864 18052 15892
rect 17635 15861 17647 15864
rect 17589 15855 17647 15861
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 20714 15892 20720 15904
rect 20312 15864 20720 15892
rect 20312 15852 20318 15864
rect 20714 15852 20720 15864
rect 20772 15852 20778 15904
rect 23845 15895 23903 15901
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 24946 15892 24952 15904
rect 23891 15864 24952 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 24946 15852 24952 15864
rect 25004 15852 25010 15904
rect 25682 15852 25688 15904
rect 25740 15892 25746 15904
rect 26421 15895 26479 15901
rect 26421 15892 26433 15895
rect 25740 15864 26433 15892
rect 25740 15852 25746 15864
rect 26421 15861 26433 15864
rect 26467 15861 26479 15895
rect 26421 15855 26479 15861
rect 32769 15895 32827 15901
rect 32769 15861 32781 15895
rect 32815 15892 32827 15895
rect 33226 15892 33232 15904
rect 32815 15864 33232 15892
rect 32815 15861 32827 15864
rect 32769 15855 32827 15861
rect 33226 15852 33232 15864
rect 33284 15852 33290 15904
rect 36630 15852 36636 15904
rect 36688 15892 36694 15904
rect 36906 15892 36912 15904
rect 36688 15864 36912 15892
rect 36688 15852 36694 15864
rect 36906 15852 36912 15864
rect 36964 15892 36970 15904
rect 37246 15892 37274 16000
rect 38654 15988 38660 16040
rect 38712 16028 38718 16040
rect 38712 16000 38757 16028
rect 38712 15988 38718 16000
rect 36964 15864 37274 15892
rect 36964 15852 36970 15864
rect 37550 15852 37556 15904
rect 37608 15892 37614 15904
rect 39040 15892 39068 16059
rect 39206 16056 39212 16068
rect 39264 16056 39270 16108
rect 39316 16105 39344 16136
rect 39301 16099 39359 16105
rect 39301 16065 39313 16099
rect 39347 16065 39359 16099
rect 39301 16059 39359 16065
rect 58158 15892 58164 15904
rect 37608 15864 39068 15892
rect 58119 15864 58164 15892
rect 37608 15852 37614 15864
rect 58158 15852 58164 15864
rect 58216 15852 58222 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 3970 15648 3976 15700
rect 4028 15688 4034 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 4028 15660 4077 15688
rect 4028 15648 4034 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 4065 15651 4123 15657
rect 4709 15691 4767 15697
rect 4709 15657 4721 15691
rect 4755 15688 4767 15691
rect 5258 15688 5264 15700
rect 4755 15660 5264 15688
rect 4755 15657 4767 15660
rect 4709 15651 4767 15657
rect 4724 15552 4752 15651
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7190 15688 7196 15700
rect 7151 15660 7196 15688
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 7374 15648 7380 15700
rect 7432 15688 7438 15700
rect 10413 15691 10471 15697
rect 10413 15688 10425 15691
rect 7432 15660 10425 15688
rect 7432 15648 7438 15660
rect 10413 15657 10425 15660
rect 10459 15657 10471 15691
rect 10413 15651 10471 15657
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 12066 15688 12072 15700
rect 11296 15660 12072 15688
rect 11296 15648 11302 15660
rect 12066 15648 12072 15660
rect 12124 15648 12130 15700
rect 12897 15691 12955 15697
rect 12897 15657 12909 15691
rect 12943 15688 12955 15691
rect 23198 15688 23204 15700
rect 12943 15660 22094 15688
rect 23159 15660 23204 15688
rect 12943 15657 12955 15660
rect 12897 15651 12955 15657
rect 7926 15580 7932 15632
rect 7984 15620 7990 15632
rect 22066 15620 22094 15660
rect 23198 15648 23204 15660
rect 23256 15648 23262 15700
rect 23290 15648 23296 15700
rect 23348 15688 23354 15700
rect 23477 15691 23535 15697
rect 23477 15688 23489 15691
rect 23348 15660 23489 15688
rect 23348 15648 23354 15660
rect 23477 15657 23489 15660
rect 23523 15657 23535 15691
rect 23477 15651 23535 15657
rect 24854 15648 24860 15700
rect 24912 15688 24918 15700
rect 25133 15691 25191 15697
rect 25133 15688 25145 15691
rect 24912 15660 25145 15688
rect 24912 15648 24918 15660
rect 25133 15657 25145 15660
rect 25179 15688 25191 15691
rect 25590 15688 25596 15700
rect 25179 15660 25596 15688
rect 25179 15657 25191 15660
rect 25133 15651 25191 15657
rect 25590 15648 25596 15660
rect 25648 15648 25654 15700
rect 25685 15691 25743 15697
rect 25685 15657 25697 15691
rect 25731 15688 25743 15691
rect 25958 15688 25964 15700
rect 25731 15660 25964 15688
rect 25731 15657 25743 15660
rect 25685 15651 25743 15657
rect 25958 15648 25964 15660
rect 26016 15648 26022 15700
rect 26513 15691 26571 15697
rect 26513 15657 26525 15691
rect 26559 15688 26571 15691
rect 27890 15688 27896 15700
rect 26559 15660 27896 15688
rect 26559 15657 26571 15660
rect 26513 15651 26571 15657
rect 27890 15648 27896 15660
rect 27948 15648 27954 15700
rect 29270 15648 29276 15700
rect 29328 15688 29334 15700
rect 29825 15691 29883 15697
rect 29825 15688 29837 15691
rect 29328 15660 29837 15688
rect 29328 15648 29334 15660
rect 29825 15657 29837 15660
rect 29871 15657 29883 15691
rect 34054 15688 34060 15700
rect 34015 15660 34060 15688
rect 29825 15651 29883 15657
rect 23014 15620 23020 15632
rect 7984 15592 9260 15620
rect 22066 15592 23020 15620
rect 7984 15580 7990 15592
rect 3896 15524 4752 15552
rect 7285 15555 7343 15561
rect 2130 15484 2136 15496
rect 2091 15456 2136 15484
rect 2130 15444 2136 15456
rect 2188 15444 2194 15496
rect 2314 15484 2320 15496
rect 2275 15456 2320 15484
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 3050 15484 3056 15496
rect 3011 15456 3056 15484
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 3418 15444 3424 15496
rect 3476 15484 3482 15496
rect 3896 15493 3924 15524
rect 7285 15521 7297 15555
rect 7331 15552 7343 15555
rect 8202 15552 8208 15564
rect 7331 15524 8208 15552
rect 7331 15521 7343 15524
rect 7285 15515 7343 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 3881 15487 3939 15493
rect 3881 15484 3893 15487
rect 3476 15456 3893 15484
rect 3476 15444 3482 15456
rect 3881 15453 3893 15456
rect 3927 15453 3939 15487
rect 3881 15447 3939 15453
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 5537 15487 5595 15493
rect 5537 15484 5549 15487
rect 4212 15456 5549 15484
rect 4212 15444 4218 15456
rect 5537 15453 5549 15456
rect 5583 15453 5595 15487
rect 5537 15447 5595 15453
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15484 5687 15487
rect 5902 15484 5908 15496
rect 5675 15456 5908 15484
rect 5675 15453 5687 15456
rect 5629 15447 5687 15453
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15484 7435 15487
rect 8294 15484 8300 15496
rect 7423 15456 8300 15484
rect 7423 15453 7435 15456
rect 7377 15447 7435 15453
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 9232 15493 9260 15592
rect 23014 15580 23020 15592
rect 23072 15580 23078 15632
rect 24762 15620 24768 15632
rect 23400 15592 24768 15620
rect 10505 15555 10563 15561
rect 10505 15521 10517 15555
rect 10551 15552 10563 15555
rect 10870 15552 10876 15564
rect 10551 15524 10876 15552
rect 10551 15521 10563 15524
rect 10505 15515 10563 15521
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 13538 15512 13544 15564
rect 13596 15552 13602 15564
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13596 15524 14105 15552
rect 13596 15512 13602 15524
rect 14093 15521 14105 15524
rect 14139 15521 14151 15555
rect 14093 15515 14151 15521
rect 18693 15555 18751 15561
rect 18693 15521 18705 15555
rect 18739 15552 18751 15555
rect 19242 15552 19248 15564
rect 18739 15524 19248 15552
rect 18739 15521 18751 15524
rect 18693 15515 18751 15521
rect 19242 15512 19248 15524
rect 19300 15552 19306 15564
rect 23400 15552 23428 15592
rect 24762 15580 24768 15592
rect 24820 15620 24826 15632
rect 29840 15620 29868 15651
rect 34054 15648 34060 15660
rect 34112 15648 34118 15700
rect 24820 15592 26464 15620
rect 29840 15592 30052 15620
rect 24820 15580 24826 15592
rect 23566 15552 23572 15564
rect 19300 15524 23428 15552
rect 23527 15524 23572 15552
rect 19300 15512 19306 15524
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 26436 15552 26464 15592
rect 27157 15555 27215 15561
rect 27157 15552 27169 15555
rect 26436 15524 27169 15552
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 8941 15447 8999 15453
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15484 9275 15487
rect 9398 15484 9404 15496
rect 9263 15456 9404 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 5350 15376 5356 15428
rect 5408 15416 5414 15428
rect 8956 15416 8984 15447
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 14366 15493 14372 15496
rect 12713 15487 12771 15493
rect 12713 15484 12725 15487
rect 10652 15456 10697 15484
rect 11532 15456 12725 15484
rect 10652 15444 10658 15456
rect 11532 15428 11560 15456
rect 12713 15453 12725 15456
rect 12759 15453 12771 15487
rect 14360 15484 14372 15493
rect 14327 15456 14372 15484
rect 12713 15447 12771 15453
rect 14360 15447 14372 15456
rect 14366 15444 14372 15447
rect 14424 15444 14430 15496
rect 16669 15487 16727 15493
rect 16669 15453 16681 15487
rect 16715 15484 16727 15487
rect 17862 15484 17868 15496
rect 16715 15456 17868 15484
rect 16715 15453 16727 15456
rect 16669 15447 16727 15453
rect 17862 15444 17868 15456
rect 17920 15444 17926 15496
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 20438 15484 20444 15496
rect 20399 15456 20444 15484
rect 20438 15444 20444 15456
rect 20496 15444 20502 15496
rect 20530 15444 20536 15496
rect 20588 15484 20594 15496
rect 22097 15487 22155 15493
rect 22097 15484 22109 15487
rect 20588 15456 22109 15484
rect 20588 15444 20594 15456
rect 22097 15453 22109 15456
rect 22143 15484 22155 15487
rect 22646 15484 22652 15496
rect 22143 15456 22652 15484
rect 22143 15453 22155 15456
rect 22097 15447 22155 15453
rect 22646 15444 22652 15456
rect 22704 15444 22710 15496
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23658 15484 23664 15496
rect 23619 15456 23664 15484
rect 23385 15447 23443 15453
rect 11514 15416 11520 15428
rect 5408 15388 11520 15416
rect 5408 15376 5414 15388
rect 11514 15376 11520 15388
rect 11572 15376 11578 15428
rect 16114 15376 16120 15428
rect 16172 15416 16178 15428
rect 16914 15419 16972 15425
rect 16914 15416 16926 15419
rect 16172 15388 16926 15416
rect 16172 15376 16178 15388
rect 16914 15385 16926 15388
rect 16960 15385 16972 15419
rect 20272 15416 20300 15444
rect 20625 15419 20683 15425
rect 20625 15416 20637 15419
rect 20272 15388 20637 15416
rect 16914 15379 16972 15385
rect 20625 15385 20637 15388
rect 20671 15385 20683 15419
rect 23400 15416 23428 15447
rect 23658 15444 23664 15456
rect 23716 15484 23722 15496
rect 26436 15493 26464 15524
rect 27157 15521 27169 15524
rect 27203 15552 27215 15555
rect 27203 15524 29960 15552
rect 27203 15521 27215 15524
rect 27157 15515 27215 15521
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 23716 15456 24409 15484
rect 23716 15444 23722 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 24397 15447 24455 15453
rect 26421 15487 26479 15493
rect 26421 15453 26433 15487
rect 26467 15453 26479 15487
rect 26602 15484 26608 15496
rect 26563 15456 26608 15484
rect 26421 15447 26479 15453
rect 26602 15444 26608 15456
rect 26660 15444 26666 15496
rect 28261 15487 28319 15493
rect 28261 15453 28273 15487
rect 28307 15484 28319 15487
rect 29822 15484 29828 15496
rect 28307 15456 29828 15484
rect 28307 15453 28319 15456
rect 28261 15447 28319 15453
rect 29822 15444 29828 15456
rect 29880 15444 29886 15496
rect 24946 15416 24952 15428
rect 23400 15388 24952 15416
rect 20625 15379 20683 15385
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 25682 15376 25688 15428
rect 25740 15416 25746 15428
rect 28077 15419 28135 15425
rect 28077 15416 28089 15419
rect 25740 15388 28089 15416
rect 25740 15376 25746 15388
rect 28077 15385 28089 15388
rect 28123 15416 28135 15419
rect 28718 15416 28724 15428
rect 28123 15388 28724 15416
rect 28123 15385 28135 15388
rect 28077 15379 28135 15385
rect 28718 15376 28724 15388
rect 28776 15376 28782 15428
rect 3237 15351 3295 15357
rect 3237 15317 3249 15351
rect 3283 15348 3295 15351
rect 3510 15348 3516 15360
rect 3283 15320 3516 15348
rect 3283 15317 3295 15320
rect 3237 15311 3295 15317
rect 3510 15308 3516 15320
rect 3568 15308 3574 15360
rect 5166 15348 5172 15360
rect 5127 15320 5172 15348
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 5810 15348 5816 15360
rect 5771 15320 5816 15348
rect 5810 15308 5816 15320
rect 5868 15308 5874 15360
rect 7006 15348 7012 15360
rect 6967 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 9950 15308 9956 15360
rect 10008 15348 10014 15360
rect 10229 15351 10287 15357
rect 10229 15348 10241 15351
rect 10008 15320 10241 15348
rect 10008 15308 10014 15320
rect 10229 15317 10241 15320
rect 10275 15317 10287 15351
rect 10229 15311 10287 15317
rect 11882 15308 11888 15360
rect 11940 15348 11946 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 11940 15320 12173 15348
rect 11940 15308 11946 15320
rect 12161 15317 12173 15320
rect 12207 15317 12219 15351
rect 12161 15311 12219 15317
rect 15286 15308 15292 15360
rect 15344 15348 15350 15360
rect 15473 15351 15531 15357
rect 15473 15348 15485 15351
rect 15344 15320 15485 15348
rect 15344 15308 15350 15320
rect 15473 15317 15485 15320
rect 15519 15317 15531 15351
rect 15473 15311 15531 15317
rect 18049 15351 18107 15357
rect 18049 15317 18061 15351
rect 18095 15348 18107 15351
rect 18138 15348 18144 15360
rect 18095 15320 18144 15348
rect 18095 15317 18107 15320
rect 18049 15311 18107 15317
rect 18138 15308 18144 15320
rect 18196 15308 18202 15360
rect 19797 15351 19855 15357
rect 19797 15317 19809 15351
rect 19843 15348 19855 15351
rect 20070 15348 20076 15360
rect 19843 15320 20076 15348
rect 19843 15317 19855 15320
rect 19797 15311 19855 15317
rect 20070 15308 20076 15320
rect 20128 15308 20134 15360
rect 20257 15351 20315 15357
rect 20257 15317 20269 15351
rect 20303 15348 20315 15351
rect 20346 15348 20352 15360
rect 20303 15320 20352 15348
rect 20303 15317 20315 15320
rect 20257 15311 20315 15317
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 27982 15308 27988 15360
rect 28040 15348 28046 15360
rect 28445 15351 28503 15357
rect 28445 15348 28457 15351
rect 28040 15320 28457 15348
rect 28040 15308 28046 15320
rect 28445 15317 28457 15320
rect 28491 15317 28503 15351
rect 29932 15348 29960 15524
rect 30024 15416 30052 15592
rect 31846 15552 31852 15564
rect 30668 15524 31852 15552
rect 30374 15484 30380 15496
rect 30335 15456 30380 15484
rect 30374 15444 30380 15456
rect 30432 15444 30438 15496
rect 30466 15444 30472 15496
rect 30524 15484 30530 15496
rect 30668 15493 30696 15524
rect 31846 15512 31852 15524
rect 31904 15512 31910 15564
rect 35069 15555 35127 15561
rect 35069 15521 35081 15555
rect 35115 15552 35127 15555
rect 35115 15524 36860 15552
rect 35115 15521 35127 15524
rect 35069 15515 35127 15521
rect 36832 15496 36860 15524
rect 30561 15487 30619 15493
rect 30561 15484 30573 15487
rect 30524 15456 30573 15484
rect 30524 15444 30530 15456
rect 30561 15453 30573 15456
rect 30607 15453 30619 15487
rect 30561 15447 30619 15453
rect 30653 15487 30711 15493
rect 30653 15453 30665 15487
rect 30699 15453 30711 15487
rect 30653 15447 30711 15453
rect 30745 15487 30803 15493
rect 30745 15453 30757 15487
rect 30791 15453 30803 15487
rect 30745 15447 30803 15453
rect 30852 15456 32720 15484
rect 30760 15416 30788 15447
rect 30024 15388 30788 15416
rect 30852 15348 30880 15456
rect 31021 15419 31079 15425
rect 31021 15385 31033 15419
rect 31067 15416 31079 15419
rect 32594 15419 32652 15425
rect 32594 15416 32606 15419
rect 31067 15388 32606 15416
rect 31067 15385 31079 15388
rect 31021 15379 31079 15385
rect 32594 15385 32606 15388
rect 32640 15385 32652 15419
rect 32692 15416 32720 15456
rect 32766 15444 32772 15496
rect 32824 15484 32830 15496
rect 32861 15487 32919 15493
rect 32861 15484 32873 15487
rect 32824 15456 32873 15484
rect 32824 15444 32830 15456
rect 32861 15453 32873 15456
rect 32907 15453 32919 15487
rect 32861 15447 32919 15453
rect 34054 15444 34060 15496
rect 34112 15484 34118 15496
rect 34701 15487 34759 15493
rect 34701 15484 34713 15487
rect 34112 15456 34713 15484
rect 34112 15444 34118 15456
rect 34701 15453 34713 15456
rect 34747 15453 34759 15487
rect 34701 15447 34759 15453
rect 34790 15444 34796 15496
rect 34848 15484 34854 15496
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34848 15456 34897 15484
rect 34848 15444 34854 15456
rect 34885 15453 34897 15456
rect 34931 15484 34943 15487
rect 35529 15487 35587 15493
rect 35529 15484 35541 15487
rect 34931 15456 35541 15484
rect 34931 15453 34943 15456
rect 34885 15447 34943 15453
rect 35529 15453 35541 15456
rect 35575 15453 35587 15487
rect 35529 15447 35587 15453
rect 35713 15487 35771 15493
rect 35713 15453 35725 15487
rect 35759 15453 35771 15487
rect 36814 15484 36820 15496
rect 36775 15456 36820 15484
rect 35713 15447 35771 15453
rect 34606 15416 34612 15428
rect 32692 15388 34612 15416
rect 32594 15379 32652 15385
rect 34606 15376 34612 15388
rect 34664 15416 34670 15428
rect 35728 15416 35756 15447
rect 36814 15444 36820 15456
rect 36872 15444 36878 15496
rect 37182 15444 37188 15496
rect 37240 15484 37246 15496
rect 37645 15487 37703 15493
rect 37645 15484 37657 15487
rect 37240 15456 37657 15484
rect 37240 15444 37246 15456
rect 37645 15453 37657 15456
rect 37691 15453 37703 15487
rect 37826 15484 37832 15496
rect 37787 15456 37832 15484
rect 37645 15447 37703 15453
rect 37826 15444 37832 15456
rect 37884 15444 37890 15496
rect 36173 15419 36231 15425
rect 36173 15416 36185 15419
rect 34664 15388 36185 15416
rect 34664 15376 34670 15388
rect 36173 15385 36185 15388
rect 36219 15385 36231 15419
rect 36173 15379 36231 15385
rect 37001 15419 37059 15425
rect 37001 15385 37013 15419
rect 37047 15416 37059 15419
rect 37274 15416 37280 15428
rect 37047 15388 37280 15416
rect 37047 15385 37059 15388
rect 37001 15379 37059 15385
rect 37274 15376 37280 15388
rect 37332 15416 37338 15428
rect 37458 15416 37464 15428
rect 37332 15388 37464 15416
rect 37332 15376 37338 15388
rect 37458 15376 37464 15388
rect 37516 15376 37522 15428
rect 29932 15320 30880 15348
rect 28445 15311 28503 15317
rect 31294 15308 31300 15360
rect 31352 15348 31358 15360
rect 31481 15351 31539 15357
rect 31481 15348 31493 15351
rect 31352 15320 31493 15348
rect 31352 15308 31358 15320
rect 31481 15317 31493 15320
rect 31527 15317 31539 15351
rect 31481 15311 31539 15317
rect 35713 15351 35771 15357
rect 35713 15317 35725 15351
rect 35759 15348 35771 15351
rect 37090 15348 37096 15360
rect 35759 15320 37096 15348
rect 35759 15317 35771 15320
rect 35713 15311 35771 15317
rect 37090 15308 37096 15320
rect 37148 15308 37154 15360
rect 37185 15351 37243 15357
rect 37185 15317 37197 15351
rect 37231 15348 37243 15351
rect 37550 15348 37556 15360
rect 37231 15320 37556 15348
rect 37231 15317 37243 15320
rect 37185 15311 37243 15317
rect 37550 15308 37556 15320
rect 37608 15308 37614 15360
rect 38013 15351 38071 15357
rect 38013 15317 38025 15351
rect 38059 15348 38071 15351
rect 38378 15348 38384 15360
rect 38059 15320 38384 15348
rect 38059 15317 38071 15320
rect 38013 15311 38071 15317
rect 38378 15308 38384 15320
rect 38436 15308 38442 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 2958 15144 2964 15156
rect 2871 15116 2964 15144
rect 2958 15104 2964 15116
rect 3016 15144 3022 15156
rect 4154 15144 4160 15156
rect 3016 15116 4160 15144
rect 3016 15104 3022 15116
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 14182 15144 14188 15156
rect 14143 15116 14188 15144
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 14826 15104 14832 15156
rect 14884 15144 14890 15156
rect 15105 15147 15163 15153
rect 15105 15144 15117 15147
rect 14884 15116 15117 15144
rect 14884 15104 14890 15116
rect 15105 15113 15117 15116
rect 15151 15113 15163 15147
rect 16666 15144 16672 15156
rect 16627 15116 16672 15144
rect 15105 15107 15163 15113
rect 16666 15104 16672 15116
rect 16724 15104 16730 15156
rect 18138 15144 18144 15156
rect 16868 15116 18144 15144
rect 2774 15076 2780 15088
rect 1596 15048 2780 15076
rect 1596 15017 1624 15048
rect 2774 15036 2780 15048
rect 2832 15036 2838 15088
rect 4614 15076 4620 15088
rect 3436 15048 4620 15076
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 1848 15011 1906 15017
rect 1848 14977 1860 15011
rect 1894 15008 1906 15011
rect 2222 15008 2228 15020
rect 1894 14980 2228 15008
rect 1894 14977 1906 14980
rect 1848 14971 1906 14977
rect 2222 14968 2228 14980
rect 2280 14968 2286 15020
rect 2792 15008 2820 15036
rect 3436 15017 3464 15048
rect 4614 15036 4620 15048
rect 4672 15076 4678 15088
rect 16868 15085 16896 15116
rect 18138 15104 18144 15116
rect 18196 15144 18202 15156
rect 18196 15116 21036 15144
rect 18196 15104 18202 15116
rect 16853 15079 16911 15085
rect 4672 15048 6408 15076
rect 4672 15036 4678 15048
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 2792 14980 3433 15008
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 6380 15017 6408 15048
rect 16853 15045 16865 15079
rect 16899 15045 16911 15079
rect 16853 15039 16911 15045
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 20910 15079 20968 15085
rect 20910 15076 20922 15079
rect 20864 15048 20922 15076
rect 20864 15036 20870 15048
rect 20910 15045 20922 15048
rect 20956 15045 20968 15079
rect 21008 15076 21036 15116
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 22002 15144 22008 15156
rect 21140 15116 22008 15144
rect 21140 15104 21146 15116
rect 22002 15104 22008 15116
rect 22060 15144 22066 15156
rect 22833 15147 22891 15153
rect 22060 15116 22508 15144
rect 22060 15104 22066 15116
rect 22480 15085 22508 15116
rect 22833 15113 22845 15147
rect 22879 15144 22891 15147
rect 23198 15144 23204 15156
rect 22879 15116 23204 15144
rect 22879 15113 22891 15116
rect 22833 15107 22891 15113
rect 23198 15104 23204 15116
rect 23256 15104 23262 15156
rect 29822 15144 29828 15156
rect 23492 15116 25820 15144
rect 29783 15116 29828 15144
rect 22465 15079 22523 15085
rect 21008 15048 22416 15076
rect 20910 15039 20968 15045
rect 3677 15011 3735 15017
rect 3677 15008 3689 15011
rect 3568 14980 3689 15008
rect 3568 14968 3574 14980
rect 3677 14977 3689 14980
rect 3723 14977 3735 15011
rect 3677 14971 3735 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 6632 15011 6690 15017
rect 6632 14977 6644 15011
rect 6678 15008 6690 15011
rect 6914 15008 6920 15020
rect 6678 14980 6920 15008
rect 6678 14977 6690 14980
rect 6632 14971 6690 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 15286 15008 15292 15020
rect 15247 14980 15292 15008
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15473 15011 15531 15017
rect 15473 14977 15485 15011
rect 15519 15008 15531 15011
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 15519 14980 17049 15008
rect 15519 14977 15531 14980
rect 15473 14971 15531 14977
rect 17037 14977 17049 14980
rect 17083 15008 17095 15011
rect 17770 15008 17776 15020
rect 17083 14980 17776 15008
rect 17083 14977 17095 14980
rect 17037 14971 17095 14977
rect 17770 14968 17776 14980
rect 17828 14968 17834 15020
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 17957 15011 18015 15017
rect 17957 15008 17969 15011
rect 17920 14980 17969 15008
rect 17920 14968 17926 14980
rect 17957 14977 17969 14980
rect 18003 14977 18015 15011
rect 17957 14971 18015 14977
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18213 15011 18271 15017
rect 18213 15008 18225 15011
rect 18104 14980 18225 15008
rect 18104 14968 18110 14980
rect 18213 14977 18225 14980
rect 18259 14977 18271 15011
rect 20530 15008 20536 15020
rect 18213 14971 18271 14977
rect 19904 14980 20536 15008
rect 19334 14872 19340 14884
rect 19247 14844 19340 14872
rect 19334 14832 19340 14844
rect 19392 14872 19398 14884
rect 19904 14872 19932 14980
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 22281 15011 22339 15017
rect 22281 14977 22293 15011
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 21177 14943 21235 14949
rect 21177 14909 21189 14943
rect 21223 14940 21235 14943
rect 21450 14940 21456 14952
rect 21223 14912 21456 14940
rect 21223 14909 21235 14912
rect 21177 14903 21235 14909
rect 21450 14900 21456 14912
rect 21508 14940 21514 14952
rect 22094 14940 22100 14952
rect 21508 14912 22100 14940
rect 21508 14900 21514 14912
rect 22094 14900 22100 14912
rect 22152 14900 22158 14952
rect 19392 14844 19932 14872
rect 19392 14832 19398 14844
rect 4798 14804 4804 14816
rect 4759 14776 4804 14804
rect 4798 14764 4804 14776
rect 4856 14764 4862 14816
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12802 14804 12808 14816
rect 12492 14776 12808 14804
rect 12492 14764 12498 14776
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 19797 14807 19855 14813
rect 19797 14773 19809 14807
rect 19843 14804 19855 14807
rect 20438 14804 20444 14816
rect 19843 14776 20444 14804
rect 19843 14773 19855 14776
rect 19797 14767 19855 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 20530 14764 20536 14816
rect 20588 14804 20594 14816
rect 22296 14804 22324 14971
rect 22388 14872 22416 15048
rect 22465 15045 22477 15079
rect 22511 15045 22523 15079
rect 22465 15039 22523 15045
rect 22557 15079 22615 15085
rect 22557 15045 22569 15079
rect 22603 15076 22615 15079
rect 22922 15076 22928 15088
rect 22603 15048 22928 15076
rect 22603 15045 22615 15048
rect 22557 15039 22615 15045
rect 22922 15036 22928 15048
rect 22980 15076 22986 15088
rect 23492 15076 23520 15116
rect 22980 15048 23520 15076
rect 23569 15079 23627 15085
rect 22980 15036 22986 15048
rect 23569 15045 23581 15079
rect 23615 15076 23627 15079
rect 25130 15076 25136 15088
rect 23615 15048 25136 15076
rect 23615 15045 23627 15048
rect 23569 15039 23627 15045
rect 25130 15036 25136 15048
rect 25188 15036 25194 15088
rect 25792 15085 25820 15116
rect 29822 15104 29828 15116
rect 29880 15104 29886 15156
rect 30466 15104 30472 15156
rect 30524 15144 30530 15156
rect 31205 15147 31263 15153
rect 31205 15144 31217 15147
rect 30524 15116 31217 15144
rect 30524 15104 30530 15116
rect 31205 15113 31217 15116
rect 31251 15113 31263 15147
rect 34054 15144 34060 15156
rect 34015 15116 34060 15144
rect 31205 15107 31263 15113
rect 34054 15104 34060 15116
rect 34112 15104 34118 15156
rect 34977 15147 35035 15153
rect 34977 15113 34989 15147
rect 35023 15144 35035 15147
rect 35894 15144 35900 15156
rect 35023 15116 35900 15144
rect 35023 15113 35035 15116
rect 34977 15107 35035 15113
rect 35894 15104 35900 15116
rect 35952 15144 35958 15156
rect 37182 15144 37188 15156
rect 35952 15116 37188 15144
rect 35952 15104 35958 15116
rect 37182 15104 37188 15116
rect 37240 15104 37246 15156
rect 37274 15104 37280 15156
rect 37332 15144 37338 15156
rect 38657 15147 38715 15153
rect 38657 15144 38669 15147
rect 37332 15116 38669 15144
rect 37332 15104 37338 15116
rect 38657 15113 38669 15116
rect 38703 15113 38715 15147
rect 38657 15107 38715 15113
rect 25777 15079 25835 15085
rect 25777 15045 25789 15079
rect 25823 15045 25835 15079
rect 25777 15039 25835 15045
rect 30742 15036 30748 15088
rect 30800 15076 30806 15088
rect 31573 15079 31631 15085
rect 31573 15076 31585 15079
rect 30800 15048 31585 15076
rect 30800 15036 30806 15048
rect 31573 15045 31585 15048
rect 31619 15045 31631 15079
rect 31573 15039 31631 15045
rect 32766 15036 32772 15088
rect 32824 15076 32830 15088
rect 36725 15079 36783 15085
rect 32824 15048 33548 15076
rect 32824 15036 32830 15048
rect 22646 15008 22652 15020
rect 22607 14980 22652 15008
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 23293 15011 23351 15017
rect 23293 15008 23305 15011
rect 22756 14980 23305 15008
rect 22756 14872 22784 14980
rect 23293 14977 23305 14980
rect 23339 14977 23351 15011
rect 23293 14971 23351 14977
rect 23382 14968 23388 15020
rect 23440 15008 23446 15020
rect 23477 15011 23535 15017
rect 23477 15008 23489 15011
rect 23440 14980 23489 15008
rect 23440 14968 23446 14980
rect 23477 14977 23489 14980
rect 23523 14977 23535 15011
rect 23477 14971 23535 14977
rect 23658 14968 23664 15020
rect 23716 15008 23722 15020
rect 24489 15011 24547 15017
rect 23716 14980 24440 15008
rect 23716 14968 23722 14980
rect 22388 14844 22784 14872
rect 23198 14832 23204 14884
rect 23256 14872 23262 14884
rect 24305 14875 24363 14881
rect 24305 14872 24317 14875
rect 23256 14844 24317 14872
rect 23256 14832 23262 14844
rect 24305 14841 24317 14844
rect 24351 14841 24363 14875
rect 24412 14872 24440 14980
rect 24489 14977 24501 15011
rect 24535 15008 24547 15011
rect 24765 15011 24823 15017
rect 24535 14980 24716 15008
rect 24535 14977 24547 14980
rect 24489 14971 24547 14977
rect 24578 14940 24584 14952
rect 24539 14912 24584 14940
rect 24578 14900 24584 14912
rect 24636 14900 24642 14952
rect 24688 14940 24716 14980
rect 24765 14977 24777 15011
rect 24811 15008 24823 15011
rect 24854 15008 24860 15020
rect 24811 14980 24860 15008
rect 24811 14977 24823 14980
rect 24765 14971 24823 14977
rect 24854 14968 24860 14980
rect 24912 14968 24918 15020
rect 25593 15011 25651 15017
rect 25593 14977 25605 15011
rect 25639 15008 25651 15011
rect 25682 15008 25688 15020
rect 25639 14980 25688 15008
rect 25639 14977 25651 14980
rect 25593 14971 25651 14977
rect 25682 14968 25688 14980
rect 25740 14968 25746 15020
rect 28534 14968 28540 15020
rect 28592 15008 28598 15020
rect 28701 15011 28759 15017
rect 28701 15008 28713 15011
rect 28592 14980 28713 15008
rect 28592 14968 28598 14980
rect 28701 14977 28713 14980
rect 28747 14977 28759 15011
rect 28701 14971 28759 14977
rect 31294 14968 31300 15020
rect 31352 15008 31358 15020
rect 31389 15011 31447 15017
rect 31389 15008 31401 15011
rect 31352 14980 31401 15008
rect 31352 14968 31358 14980
rect 31389 14977 31401 14980
rect 31435 14977 31447 15011
rect 31389 14971 31447 14977
rect 33226 14968 33232 15020
rect 33284 15017 33290 15020
rect 33520 15017 33548 15048
rect 36725 15045 36737 15079
rect 36771 15076 36783 15079
rect 38105 15079 38163 15085
rect 36771 15048 37872 15076
rect 36771 15045 36783 15048
rect 36725 15039 36783 15045
rect 33284 15008 33296 15017
rect 33505 15011 33563 15017
rect 33284 14980 33329 15008
rect 33284 14971 33296 14980
rect 33505 14977 33517 15011
rect 33551 14977 33563 15011
rect 33505 14971 33563 14977
rect 33284 14968 33290 14971
rect 34514 14968 34520 15020
rect 34572 15008 34578 15020
rect 34793 15011 34851 15017
rect 34793 15008 34805 15011
rect 34572 14980 34805 15008
rect 34572 14968 34578 14980
rect 34793 14977 34805 14980
rect 34839 14977 34851 15011
rect 37461 15011 37519 15017
rect 37461 15008 37473 15011
rect 34793 14971 34851 14977
rect 36648 14980 37473 15008
rect 25314 14940 25320 14952
rect 24688 14912 25320 14940
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 28442 14940 28448 14952
rect 28403 14912 28448 14940
rect 28442 14900 28448 14912
rect 28500 14900 28506 14952
rect 34054 14900 34060 14952
rect 34112 14940 34118 14952
rect 34609 14943 34667 14949
rect 34609 14940 34621 14943
rect 34112 14912 34621 14940
rect 34112 14900 34118 14912
rect 34609 14909 34621 14912
rect 34655 14909 34667 14943
rect 34609 14903 34667 14909
rect 34698 14900 34704 14952
rect 34756 14940 34762 14952
rect 36648 14940 36676 14980
rect 34756 14912 36676 14940
rect 34756 14900 34762 14912
rect 26602 14872 26608 14884
rect 24412 14844 26608 14872
rect 24305 14835 24363 14841
rect 26602 14832 26608 14844
rect 26660 14832 26666 14884
rect 37016 14872 37044 14980
rect 37461 14977 37473 14980
rect 37507 14977 37519 15011
rect 37461 14971 37519 14977
rect 37550 14968 37556 15020
rect 37608 15008 37614 15020
rect 37844 15017 37872 15048
rect 38105 15045 38117 15079
rect 38151 15076 38163 15079
rect 39770 15079 39828 15085
rect 39770 15076 39782 15079
rect 38151 15048 39782 15076
rect 38151 15045 38163 15048
rect 38105 15039 38163 15045
rect 39770 15045 39782 15048
rect 39816 15045 39828 15079
rect 39770 15039 39828 15045
rect 37645 15011 37703 15017
rect 37645 15008 37657 15011
rect 37608 14980 37657 15008
rect 37608 14968 37614 14980
rect 37645 14977 37657 14980
rect 37691 14977 37703 15011
rect 37645 14971 37703 14977
rect 37737 15011 37795 15017
rect 37737 14977 37749 15011
rect 37783 14977 37795 15011
rect 37737 14971 37795 14977
rect 37829 15011 37887 15017
rect 37829 14977 37841 15011
rect 37875 15008 37887 15011
rect 38562 15008 38568 15020
rect 37875 14980 38568 15008
rect 37875 14977 37887 14980
rect 37829 14971 37887 14977
rect 37090 14900 37096 14952
rect 37148 14940 37154 14952
rect 37752 14940 37780 14971
rect 38562 14968 38568 14980
rect 38620 14968 38626 15020
rect 40034 15008 40040 15020
rect 39995 14980 40040 15008
rect 40034 14968 40040 14980
rect 40092 14968 40098 15020
rect 37148 14912 37780 14940
rect 37148 14900 37154 14912
rect 39022 14872 39028 14884
rect 37016 14844 39028 14872
rect 39022 14832 39028 14844
rect 39080 14832 39086 14884
rect 20588 14776 22324 14804
rect 20588 14764 20594 14776
rect 22646 14764 22652 14816
rect 22704 14804 22710 14816
rect 23658 14804 23664 14816
rect 22704 14776 23664 14804
rect 22704 14764 22710 14776
rect 23658 14764 23664 14776
rect 23716 14764 23722 14816
rect 23842 14804 23848 14816
rect 23803 14776 23848 14804
rect 23842 14764 23848 14776
rect 23900 14764 23906 14816
rect 24486 14804 24492 14816
rect 24447 14776 24492 14804
rect 24486 14764 24492 14776
rect 24544 14764 24550 14816
rect 25961 14807 26019 14813
rect 25961 14773 25973 14807
rect 26007 14804 26019 14807
rect 26326 14804 26332 14816
rect 26007 14776 26332 14804
rect 26007 14773 26019 14776
rect 25961 14767 26019 14773
rect 26326 14764 26332 14776
rect 26384 14764 26390 14816
rect 27154 14764 27160 14816
rect 27212 14804 27218 14816
rect 27430 14804 27436 14816
rect 27212 14776 27436 14804
rect 27212 14764 27218 14776
rect 27430 14764 27436 14776
rect 27488 14804 27494 14816
rect 28350 14804 28356 14816
rect 27488 14776 28356 14804
rect 27488 14764 27494 14776
rect 28350 14764 28356 14776
rect 28408 14764 28414 14816
rect 32030 14764 32036 14816
rect 32088 14804 32094 14816
rect 32125 14807 32183 14813
rect 32125 14804 32137 14807
rect 32088 14776 32137 14804
rect 32088 14764 32094 14776
rect 32125 14773 32137 14776
rect 32171 14773 32183 14807
rect 32125 14767 32183 14773
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 2314 14560 2320 14612
rect 2372 14600 2378 14612
rect 2501 14603 2559 14609
rect 2501 14600 2513 14603
rect 2372 14572 2513 14600
rect 2372 14560 2378 14572
rect 2501 14569 2513 14572
rect 2547 14569 2559 14603
rect 2501 14563 2559 14569
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3108 14572 3801 14600
rect 3108 14560 3114 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 6914 14600 6920 14612
rect 6875 14572 6920 14600
rect 3789 14563 3847 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 7515 14572 11621 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 11609 14563 11667 14569
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 3878 14532 3884 14544
rect 2188 14504 3884 14532
rect 2188 14492 2194 14504
rect 3878 14492 3884 14504
rect 3936 14532 3942 14544
rect 3936 14504 4200 14532
rect 3936 14492 3942 14504
rect 2958 14464 2964 14476
rect 2919 14436 2964 14464
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14464 3203 14467
rect 3602 14464 3608 14476
rect 3191 14436 3608 14464
rect 3191 14433 3203 14436
rect 3145 14427 3203 14433
rect 3602 14424 3608 14436
rect 3660 14464 3666 14476
rect 4062 14464 4068 14476
rect 3660 14436 4068 14464
rect 3660 14424 3666 14436
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 4172 14473 4200 14504
rect 6270 14492 6276 14544
rect 6328 14532 6334 14544
rect 7484 14532 7512 14563
rect 13170 14560 13176 14612
rect 13228 14600 13234 14612
rect 17310 14600 17316 14612
rect 13228 14572 17316 14600
rect 13228 14560 13234 14572
rect 17310 14560 17316 14572
rect 17368 14560 17374 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19978 14600 19984 14612
rect 19392 14572 19984 14600
rect 19392 14560 19398 14572
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 20901 14603 20959 14609
rect 20901 14600 20913 14603
rect 20864 14572 20913 14600
rect 20864 14560 20870 14572
rect 20901 14569 20913 14572
rect 20947 14569 20959 14603
rect 20901 14563 20959 14569
rect 23842 14560 23848 14612
rect 23900 14600 23906 14612
rect 24581 14603 24639 14609
rect 24581 14600 24593 14603
rect 23900 14572 24593 14600
rect 23900 14560 23906 14572
rect 24581 14569 24593 14572
rect 24627 14569 24639 14603
rect 27798 14600 27804 14612
rect 24581 14563 24639 14569
rect 25608 14572 27804 14600
rect 21726 14532 21732 14544
rect 6328 14504 7512 14532
rect 20272 14504 21732 14532
rect 6328 14492 6334 14504
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14433 4215 14467
rect 4157 14427 4215 14433
rect 4798 14424 4804 14476
rect 4856 14464 4862 14476
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 4856 14436 5457 14464
rect 4856 14424 4862 14436
rect 5445 14433 5457 14436
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 5810 14424 5816 14476
rect 5868 14464 5874 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 5868 14436 6469 14464
rect 5868 14424 5874 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14464 6607 14467
rect 7190 14464 7196 14476
rect 6595 14436 7196 14464
rect 6595 14433 6607 14436
rect 6549 14427 6607 14433
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 13538 14464 13544 14476
rect 11011 14436 13544 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 3418 14396 3424 14408
rect 2915 14368 3424 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 3418 14356 3424 14368
rect 3476 14356 3482 14408
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 5537 14399 5595 14405
rect 5537 14365 5549 14399
rect 5583 14396 5595 14399
rect 5902 14396 5908 14408
rect 5583 14368 5908 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14396 6239 14399
rect 6270 14396 6276 14408
rect 6227 14368 6276 14396
rect 6227 14365 6239 14368
rect 6181 14359 6239 14365
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 6365 14399 6423 14405
rect 6365 14365 6377 14399
rect 6411 14365 6423 14399
rect 6365 14359 6423 14365
rect 6733 14399 6791 14405
rect 6733 14365 6745 14399
rect 6779 14396 6791 14399
rect 7098 14396 7104 14408
rect 6779 14368 7104 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 5077 14331 5135 14337
rect 5077 14297 5089 14331
rect 5123 14328 5135 14331
rect 5166 14328 5172 14340
rect 5123 14300 5172 14328
rect 5123 14297 5135 14300
rect 5077 14291 5135 14297
rect 5166 14288 5172 14300
rect 5224 14328 5230 14340
rect 6086 14328 6092 14340
rect 5224 14300 6092 14328
rect 5224 14288 5230 14300
rect 6086 14288 6092 14300
rect 6144 14288 6150 14340
rect 6380 14328 6408 14359
rect 7098 14356 7104 14368
rect 7156 14396 7162 14408
rect 7742 14396 7748 14408
rect 7156 14368 7748 14396
rect 7156 14356 7162 14368
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 10226 14396 10232 14408
rect 8260 14368 10232 14396
rect 8260 14356 8266 14368
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10870 14356 10876 14408
rect 10928 14396 10934 14408
rect 20272 14405 20300 14504
rect 21726 14492 21732 14504
rect 21784 14492 21790 14544
rect 23382 14532 23388 14544
rect 23216 14504 23388 14532
rect 20257 14399 20315 14405
rect 10928 14368 12434 14396
rect 10928 14356 10934 14368
rect 7006 14328 7012 14340
rect 6380 14300 7012 14328
rect 7006 14288 7012 14300
rect 7064 14288 7070 14340
rect 10134 14288 10140 14340
rect 10192 14328 10198 14340
rect 10698 14331 10756 14337
rect 10698 14328 10710 14331
rect 10192 14300 10710 14328
rect 10192 14288 10198 14300
rect 10698 14297 10710 14300
rect 10744 14297 10756 14331
rect 11514 14328 11520 14340
rect 11475 14300 11520 14328
rect 10698 14291 10756 14297
rect 11514 14288 11520 14300
rect 11572 14288 11578 14340
rect 5721 14263 5779 14269
rect 5721 14229 5733 14263
rect 5767 14260 5779 14263
rect 7282 14260 7288 14272
rect 5767 14232 7288 14260
rect 5767 14229 5779 14232
rect 5721 14223 5779 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 9582 14260 9588 14272
rect 9543 14232 9588 14260
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 12406 14260 12434 14368
rect 20257 14365 20269 14399
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20441 14396 20499 14402
rect 20404 14368 20453 14396
rect 20404 14356 20410 14368
rect 20441 14362 20453 14368
rect 20487 14362 20499 14396
rect 20441 14356 20499 14362
rect 20530 14356 20536 14408
rect 20588 14396 20594 14408
rect 20671 14399 20729 14405
rect 20588 14368 20633 14396
rect 20588 14356 20594 14368
rect 20671 14365 20683 14399
rect 20717 14396 20729 14399
rect 21082 14396 21088 14408
rect 20717 14368 21088 14396
rect 20717 14365 20729 14368
rect 20671 14359 20729 14365
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 23017 14399 23075 14405
rect 23017 14396 23029 14399
rect 21192 14368 23029 14396
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 21192 14328 21220 14368
rect 23017 14365 23029 14368
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 15344 14300 21220 14328
rect 21453 14331 21511 14337
rect 15344 14288 15350 14300
rect 21453 14297 21465 14331
rect 21499 14328 21511 14331
rect 21726 14328 21732 14340
rect 21499 14300 21732 14328
rect 21499 14297 21511 14300
rect 21453 14291 21511 14297
rect 21726 14288 21732 14300
rect 21784 14288 21790 14340
rect 22002 14288 22008 14340
rect 22060 14328 22066 14340
rect 23216 14337 23244 14504
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 23569 14535 23627 14541
rect 23569 14501 23581 14535
rect 23615 14532 23627 14535
rect 24486 14532 24492 14544
rect 23615 14504 24492 14532
rect 23615 14501 23627 14504
rect 23569 14495 23627 14501
rect 24486 14492 24492 14504
rect 24544 14492 24550 14544
rect 25608 14532 25636 14572
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 28534 14600 28540 14612
rect 28495 14572 28540 14600
rect 28534 14560 28540 14572
rect 28592 14560 28598 14612
rect 34149 14603 34207 14609
rect 34149 14569 34161 14603
rect 34195 14600 34207 14603
rect 34606 14600 34612 14612
rect 34195 14572 34612 14600
rect 34195 14569 34207 14572
rect 34149 14563 34207 14569
rect 34606 14560 34612 14572
rect 34664 14560 34670 14612
rect 28074 14532 28080 14544
rect 24596 14504 25636 14532
rect 27816 14504 28080 14532
rect 23385 14399 23443 14405
rect 23385 14365 23397 14399
rect 23431 14396 23443 14399
rect 23658 14396 23664 14408
rect 23431 14368 23664 14396
rect 23431 14365 23443 14368
rect 23385 14359 23443 14365
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 24596 14405 24624 14504
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 24673 14399 24731 14405
rect 24673 14365 24685 14399
rect 24719 14396 24731 14399
rect 24857 14399 24915 14405
rect 24719 14368 24808 14396
rect 24719 14365 24731 14368
rect 24673 14359 24731 14365
rect 23201 14331 23259 14337
rect 23201 14328 23213 14331
rect 22060 14300 23213 14328
rect 22060 14288 22066 14300
rect 23201 14297 23213 14300
rect 23247 14297 23259 14331
rect 23201 14291 23259 14297
rect 23290 14288 23296 14340
rect 23348 14328 23354 14340
rect 23348 14300 23393 14328
rect 23348 14288 23354 14300
rect 24397 14263 24455 14269
rect 24397 14260 24409 14263
rect 12406 14232 24409 14260
rect 24397 14229 24409 14232
rect 24443 14229 24455 14263
rect 24397 14223 24455 14229
rect 24486 14220 24492 14272
rect 24544 14260 24550 14272
rect 24780 14260 24808 14368
rect 24857 14365 24869 14399
rect 24903 14396 24915 14399
rect 25958 14396 25964 14408
rect 24903 14368 25964 14396
rect 24903 14365 24915 14368
rect 24857 14359 24915 14365
rect 25958 14356 25964 14368
rect 26016 14356 26022 14408
rect 27816 14396 27844 14504
rect 28074 14492 28080 14504
rect 28132 14532 28138 14544
rect 32306 14532 32312 14544
rect 28132 14504 32312 14532
rect 28132 14492 28138 14504
rect 32306 14492 32312 14504
rect 32364 14492 32370 14544
rect 34624 14464 34652 14560
rect 36541 14467 36599 14473
rect 34624 14436 35112 14464
rect 27881 14399 27939 14405
rect 27881 14396 27893 14399
rect 27816 14368 27893 14396
rect 27881 14365 27893 14368
rect 27927 14365 27939 14399
rect 27881 14359 27939 14365
rect 27982 14356 27988 14408
rect 28040 14396 28046 14408
rect 28077 14399 28135 14405
rect 28077 14396 28089 14399
rect 28040 14368 28089 14396
rect 28040 14356 28046 14368
rect 28077 14365 28089 14368
rect 28123 14365 28135 14399
rect 28077 14359 28135 14365
rect 28169 14399 28227 14405
rect 28169 14365 28181 14399
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 25682 14288 25688 14340
rect 25740 14328 25746 14340
rect 25869 14331 25927 14337
rect 25869 14328 25881 14331
rect 25740 14300 25881 14328
rect 25740 14288 25746 14300
rect 25869 14297 25881 14300
rect 25915 14297 25927 14331
rect 25869 14291 25927 14297
rect 26050 14288 26056 14340
rect 26108 14328 26114 14340
rect 26237 14331 26295 14337
rect 26108 14300 26153 14328
rect 26108 14288 26114 14300
rect 26237 14297 26249 14331
rect 26283 14328 26295 14331
rect 27430 14328 27436 14340
rect 26283 14300 27436 14328
rect 26283 14297 26295 14300
rect 26237 14291 26295 14297
rect 27430 14288 27436 14300
rect 27488 14288 27494 14340
rect 28184 14328 28212 14359
rect 28258 14356 28264 14408
rect 28316 14396 28322 14408
rect 28316 14368 28361 14396
rect 28316 14356 28322 14368
rect 29454 14356 29460 14408
rect 29512 14396 29518 14408
rect 29733 14399 29791 14405
rect 29733 14396 29745 14399
rect 29512 14368 29745 14396
rect 29512 14356 29518 14368
rect 29733 14365 29745 14368
rect 29779 14396 29791 14399
rect 30282 14396 30288 14408
rect 29779 14368 30288 14396
rect 29779 14365 29791 14368
rect 29733 14359 29791 14365
rect 30282 14356 30288 14368
rect 30340 14356 30346 14408
rect 34514 14356 34520 14408
rect 34572 14396 34578 14408
rect 35084 14405 35112 14436
rect 36541 14433 36553 14467
rect 36587 14464 36599 14467
rect 36814 14464 36820 14476
rect 36587 14436 36820 14464
rect 36587 14433 36599 14436
rect 36541 14427 36599 14433
rect 36814 14424 36820 14436
rect 36872 14424 36878 14476
rect 38749 14467 38807 14473
rect 38749 14433 38761 14467
rect 38795 14464 38807 14467
rect 40218 14464 40224 14476
rect 38795 14436 40224 14464
rect 38795 14433 38807 14436
rect 38749 14427 38807 14433
rect 40218 14424 40224 14436
rect 40276 14424 40282 14476
rect 34885 14399 34943 14405
rect 34885 14396 34897 14399
rect 34572 14368 34897 14396
rect 34572 14356 34578 14368
rect 34885 14365 34897 14368
rect 34931 14365 34943 14399
rect 34885 14359 34943 14365
rect 35069 14399 35127 14405
rect 35069 14365 35081 14399
rect 35115 14365 35127 14399
rect 36262 14396 36268 14408
rect 36223 14368 36268 14396
rect 35069 14359 35127 14365
rect 36262 14356 36268 14368
rect 36320 14356 36326 14408
rect 37090 14356 37096 14408
rect 37148 14396 37154 14408
rect 37185 14399 37243 14405
rect 37185 14396 37197 14399
rect 37148 14368 37197 14396
rect 37148 14356 37154 14368
rect 37185 14365 37197 14368
rect 37231 14365 37243 14399
rect 37185 14359 37243 14365
rect 38194 14356 38200 14408
rect 38252 14396 38258 14408
rect 38473 14399 38531 14405
rect 38473 14396 38485 14399
rect 38252 14368 38485 14396
rect 38252 14356 38258 14368
rect 38473 14365 38485 14368
rect 38519 14365 38531 14399
rect 38473 14359 38531 14365
rect 39853 14399 39911 14405
rect 39853 14365 39865 14399
rect 39899 14365 39911 14399
rect 39853 14359 39911 14365
rect 40129 14399 40187 14405
rect 40129 14365 40141 14399
rect 40175 14396 40187 14399
rect 40678 14396 40684 14408
rect 40175 14368 40684 14396
rect 40175 14365 40187 14368
rect 40129 14359 40187 14365
rect 28350 14328 28356 14340
rect 28184 14300 28356 14328
rect 28350 14288 28356 14300
rect 28408 14288 28414 14340
rect 28718 14288 28724 14340
rect 28776 14328 28782 14340
rect 29549 14331 29607 14337
rect 29549 14328 29561 14331
rect 28776 14300 29561 14328
rect 28776 14288 28782 14300
rect 29549 14297 29561 14300
rect 29595 14297 29607 14331
rect 29549 14291 29607 14297
rect 38286 14288 38292 14340
rect 38344 14328 38350 14340
rect 39868 14328 39896 14359
rect 40678 14356 40684 14368
rect 40736 14356 40742 14408
rect 58158 14396 58164 14408
rect 58119 14368 58164 14396
rect 58158 14356 58164 14368
rect 58216 14356 58222 14408
rect 38344 14300 39896 14328
rect 38344 14288 38350 14300
rect 25314 14260 25320 14272
rect 24544 14232 24808 14260
rect 25275 14232 25320 14260
rect 24544 14220 24550 14232
rect 25314 14220 25320 14232
rect 25372 14220 25378 14272
rect 25958 14220 25964 14272
rect 26016 14260 26022 14272
rect 26697 14263 26755 14269
rect 26697 14260 26709 14263
rect 26016 14232 26709 14260
rect 26016 14220 26022 14232
rect 26697 14229 26709 14232
rect 26743 14229 26755 14263
rect 26697 14223 26755 14229
rect 27341 14263 27399 14269
rect 27341 14229 27353 14263
rect 27387 14260 27399 14263
rect 28258 14260 28264 14272
rect 27387 14232 28264 14260
rect 27387 14229 27399 14232
rect 27341 14223 27399 14229
rect 28258 14220 28264 14232
rect 28316 14220 28322 14272
rect 29914 14260 29920 14272
rect 29875 14232 29920 14260
rect 29914 14220 29920 14232
rect 29972 14220 29978 14272
rect 35069 14263 35127 14269
rect 35069 14229 35081 14263
rect 35115 14260 35127 14263
rect 35434 14260 35440 14272
rect 35115 14232 35440 14260
rect 35115 14229 35127 14232
rect 35069 14223 35127 14229
rect 35434 14220 35440 14232
rect 35492 14220 35498 14272
rect 37090 14260 37096 14272
rect 37051 14232 37096 14260
rect 37090 14220 37096 14232
rect 37148 14220 37154 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 3418 14056 3424 14068
rect 3379 14028 3424 14056
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3970 14016 3976 14068
rect 4028 14056 4034 14068
rect 5077 14059 5135 14065
rect 5077 14056 5089 14059
rect 4028 14028 5089 14056
rect 4028 14016 4034 14028
rect 5077 14025 5089 14028
rect 5123 14025 5135 14059
rect 10134 14056 10140 14068
rect 10095 14028 10140 14056
rect 5077 14019 5135 14025
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 23198 14056 23204 14068
rect 10284 14028 23204 14056
rect 10284 14016 10290 14028
rect 23198 14016 23204 14028
rect 23256 14016 23262 14068
rect 23290 14016 23296 14068
rect 23348 14056 23354 14068
rect 23477 14059 23535 14065
rect 23477 14056 23489 14059
rect 23348 14028 23489 14056
rect 23348 14016 23354 14028
rect 23477 14025 23489 14028
rect 23523 14056 23535 14059
rect 26050 14056 26056 14068
rect 23523 14028 26056 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 26050 14016 26056 14028
rect 26108 14016 26114 14068
rect 34698 14056 34704 14068
rect 27255 14028 34704 14056
rect 4798 13948 4804 14000
rect 4856 13988 4862 14000
rect 5537 13991 5595 13997
rect 5537 13988 5549 13991
rect 4856 13960 5549 13988
rect 4856 13948 4862 13960
rect 5537 13957 5549 13960
rect 5583 13957 5595 13991
rect 14274 13988 14280 14000
rect 5537 13951 5595 13957
rect 9600 13960 14280 13988
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13920 5503 13923
rect 9398 13920 9404 13932
rect 5491 13892 6500 13920
rect 9359 13892 9404 13920
rect 5491 13889 5503 13892
rect 5445 13883 5503 13889
rect 6472 13864 6500 13892
rect 9398 13880 9404 13892
rect 9456 13880 9462 13932
rect 9600 13929 9628 13960
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 16666 13948 16672 14000
rect 16724 13988 16730 14000
rect 17221 13991 17279 13997
rect 17221 13988 17233 13991
rect 16724 13960 17233 13988
rect 16724 13948 16730 13960
rect 17221 13957 17233 13960
rect 17267 13988 17279 13991
rect 19242 13988 19248 14000
rect 17267 13960 19248 13988
rect 17267 13957 17279 13960
rect 17221 13951 17279 13957
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 21082 13988 21088 14000
rect 20995 13960 21088 13988
rect 21082 13948 21088 13960
rect 21140 13988 21146 14000
rect 25222 13988 25228 14000
rect 21140 13960 25228 13988
rect 21140 13948 21146 13960
rect 25222 13948 25228 13960
rect 25280 13948 25286 14000
rect 27154 13988 27160 14000
rect 26160 13960 27160 13988
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 9953 13923 10011 13929
rect 9953 13920 9965 13923
rect 9916 13892 9965 13920
rect 9916 13880 9922 13892
rect 9953 13889 9965 13892
rect 9999 13889 10011 13923
rect 9953 13883 10011 13889
rect 13193 13923 13251 13929
rect 13193 13889 13205 13923
rect 13239 13920 13251 13923
rect 13998 13920 14004 13932
rect 13239 13892 14004 13920
rect 13239 13889 13251 13892
rect 13193 13883 13251 13889
rect 13998 13880 14004 13892
rect 14056 13880 14062 13932
rect 17310 13880 17316 13932
rect 17368 13920 17374 13932
rect 17405 13923 17463 13929
rect 17405 13920 17417 13923
rect 17368 13892 17417 13920
rect 17368 13880 17374 13892
rect 17405 13889 17417 13892
rect 17451 13889 17463 13923
rect 17405 13883 17463 13889
rect 24601 13923 24659 13929
rect 24601 13889 24613 13923
rect 24647 13920 24659 13923
rect 25590 13920 25596 13932
rect 24647 13892 25596 13920
rect 24647 13889 24659 13892
rect 24601 13883 24659 13889
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 25958 13880 25964 13932
rect 26016 13929 26022 13932
rect 26160 13929 26188 13960
rect 27154 13948 27160 13960
rect 27212 13948 27218 14000
rect 26016 13923 26065 13929
rect 26016 13889 26019 13923
rect 26053 13889 26065 13923
rect 26016 13883 26065 13889
rect 26145 13923 26203 13929
rect 26145 13889 26157 13923
rect 26191 13889 26203 13923
rect 26145 13883 26203 13889
rect 26237 13923 26295 13929
rect 26237 13889 26249 13923
rect 26283 13920 26295 13923
rect 26326 13920 26332 13932
rect 26283 13892 26332 13920
rect 26283 13889 26295 13892
rect 26237 13883 26295 13889
rect 26016 13880 26022 13883
rect 26326 13880 26332 13892
rect 26384 13880 26390 13932
rect 26418 13880 26424 13932
rect 26476 13920 26482 13932
rect 27255 13920 27283 14028
rect 34698 14016 34704 14028
rect 34756 14016 34762 14068
rect 35894 14056 35900 14068
rect 34992 14028 35900 14056
rect 27433 13991 27491 13997
rect 27433 13957 27445 13991
rect 27479 13988 27491 13991
rect 27614 13988 27620 14000
rect 27479 13960 27620 13988
rect 27479 13957 27491 13960
rect 27433 13951 27491 13957
rect 27614 13948 27620 13960
rect 27672 13988 27678 14000
rect 29546 13988 29552 14000
rect 27672 13960 29552 13988
rect 27672 13948 27678 13960
rect 29546 13948 29552 13960
rect 29604 13948 29610 14000
rect 32306 13948 32312 14000
rect 32364 13988 32370 14000
rect 32953 13991 33011 13997
rect 32953 13988 32965 13991
rect 32364 13960 32965 13988
rect 32364 13948 32370 13960
rect 32953 13957 32965 13960
rect 32999 13957 33011 13991
rect 32953 13951 33011 13957
rect 33137 13991 33195 13997
rect 33137 13957 33149 13991
rect 33183 13957 33195 13991
rect 33137 13951 33195 13957
rect 26476 13892 27283 13920
rect 26476 13880 26482 13892
rect 29270 13880 29276 13932
rect 29328 13920 29334 13932
rect 29897 13923 29955 13929
rect 29897 13920 29909 13923
rect 29328 13892 29909 13920
rect 29328 13880 29334 13892
rect 29897 13889 29909 13892
rect 29943 13889 29955 13923
rect 29897 13883 29955 13889
rect 30282 13880 30288 13932
rect 30340 13920 30346 13932
rect 30340 13892 30696 13920
rect 30340 13880 30346 13892
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13821 5779 13855
rect 6454 13852 6460 13864
rect 6415 13824 6460 13852
rect 5721 13815 5779 13821
rect 5736 13784 5764 13815
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 7340 13824 9689 13852
rect 7340 13812 7346 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 13449 13855 13507 13861
rect 9824 13824 9869 13852
rect 9824 13812 9830 13824
rect 13449 13821 13461 13855
rect 13495 13852 13507 13855
rect 14090 13852 14096 13864
rect 13495 13824 14096 13852
rect 13495 13821 13507 13824
rect 13449 13815 13507 13821
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 17589 13855 17647 13861
rect 17589 13821 17601 13855
rect 17635 13852 17647 13855
rect 17954 13852 17960 13864
rect 17635 13824 17960 13852
rect 17635 13821 17647 13824
rect 17589 13815 17647 13821
rect 17954 13812 17960 13824
rect 18012 13812 18018 13864
rect 24857 13855 24915 13861
rect 24857 13821 24869 13855
rect 24903 13852 24915 13855
rect 29641 13855 29699 13861
rect 29641 13852 29653 13855
rect 24903 13824 26096 13852
rect 24903 13821 24915 13824
rect 24857 13815 24915 13821
rect 5810 13784 5816 13796
rect 5736 13756 5816 13784
rect 5810 13744 5816 13756
rect 5868 13744 5874 13796
rect 11606 13744 11612 13796
rect 11664 13784 11670 13796
rect 12066 13784 12072 13796
rect 11664 13756 12072 13784
rect 11664 13744 11670 13756
rect 12066 13744 12072 13756
rect 12124 13744 12130 13796
rect 14366 13676 14372 13728
rect 14424 13716 14430 13728
rect 14921 13719 14979 13725
rect 14921 13716 14933 13719
rect 14424 13688 14933 13716
rect 14424 13676 14430 13688
rect 14921 13685 14933 13688
rect 14967 13685 14979 13719
rect 14921 13679 14979 13685
rect 19981 13719 20039 13725
rect 19981 13685 19993 13719
rect 20027 13716 20039 13719
rect 20162 13716 20168 13728
rect 20027 13688 20168 13716
rect 20027 13685 20039 13688
rect 19981 13679 20039 13685
rect 20162 13676 20168 13688
rect 20220 13676 20226 13728
rect 25774 13716 25780 13728
rect 25735 13688 25780 13716
rect 25774 13676 25780 13688
rect 25832 13676 25838 13728
rect 26068 13716 26096 13824
rect 28736 13824 29653 13852
rect 28736 13728 28764 13824
rect 29641 13821 29653 13824
rect 29687 13821 29699 13855
rect 30668 13852 30696 13892
rect 33152 13864 33180 13951
rect 34992 13929 35020 14028
rect 35894 14016 35900 14028
rect 35952 14016 35958 14068
rect 37366 14016 37372 14068
rect 37424 14056 37430 14068
rect 37734 14056 37740 14068
rect 37424 14028 37740 14056
rect 37424 14016 37430 14028
rect 37734 14016 37740 14028
rect 37792 14056 37798 14068
rect 37829 14059 37887 14065
rect 37829 14056 37841 14059
rect 37792 14028 37841 14056
rect 37792 14016 37798 14028
rect 37829 14025 37841 14028
rect 37875 14025 37887 14059
rect 37829 14019 37887 14025
rect 37918 14016 37924 14068
rect 37976 14056 37982 14068
rect 38749 14059 38807 14065
rect 38749 14056 38761 14059
rect 37976 14028 38761 14056
rect 37976 14016 37982 14028
rect 38749 14025 38761 14028
rect 38795 14025 38807 14059
rect 38749 14019 38807 14025
rect 35161 13991 35219 13997
rect 35161 13957 35173 13991
rect 35207 13988 35219 13991
rect 36170 13988 36176 14000
rect 35207 13960 36176 13988
rect 35207 13957 35219 13960
rect 35161 13951 35219 13957
rect 36170 13948 36176 13960
rect 36228 13948 36234 14000
rect 40218 13988 40224 14000
rect 37752 13960 40224 13988
rect 34977 13923 35035 13929
rect 34977 13889 34989 13923
rect 35023 13889 35035 13923
rect 35802 13920 35808 13932
rect 34977 13883 35035 13889
rect 35084 13892 35808 13920
rect 33134 13852 33140 13864
rect 30668 13824 31064 13852
rect 33047 13824 33140 13852
rect 29641 13815 29699 13821
rect 31036 13793 31064 13824
rect 33134 13812 33140 13824
rect 33192 13852 33198 13864
rect 35084 13852 35112 13892
rect 35802 13880 35808 13892
rect 35860 13920 35866 13932
rect 37752 13929 37780 13960
rect 40218 13948 40224 13960
rect 40276 13948 40282 14000
rect 37737 13923 37795 13929
rect 37737 13920 37749 13923
rect 35860 13892 37749 13920
rect 35860 13880 35866 13892
rect 37737 13889 37749 13892
rect 37783 13889 37795 13923
rect 37737 13883 37795 13889
rect 38838 13880 38844 13932
rect 38896 13920 38902 13932
rect 39862 13923 39920 13929
rect 39862 13920 39874 13923
rect 38896 13892 39874 13920
rect 38896 13880 38902 13892
rect 39862 13889 39874 13892
rect 39908 13889 39920 13923
rect 39862 13883 39920 13889
rect 40034 13880 40040 13932
rect 40092 13920 40098 13932
rect 40129 13923 40187 13929
rect 40129 13920 40141 13923
rect 40092 13892 40141 13920
rect 40092 13880 40098 13892
rect 40129 13889 40141 13892
rect 40175 13889 40187 13923
rect 40129 13883 40187 13889
rect 35342 13852 35348 13864
rect 33192 13824 35112 13852
rect 35303 13824 35348 13852
rect 33192 13812 33198 13824
rect 35342 13812 35348 13824
rect 35400 13812 35406 13864
rect 35434 13812 35440 13864
rect 35492 13852 35498 13864
rect 38286 13852 38292 13864
rect 35492 13824 38292 13852
rect 35492 13812 35498 13824
rect 38286 13812 38292 13824
rect 38344 13812 38350 13864
rect 31021 13787 31079 13793
rect 31021 13753 31033 13787
rect 31067 13753 31079 13787
rect 31021 13747 31079 13753
rect 26326 13716 26332 13728
rect 26068 13688 26332 13716
rect 26326 13676 26332 13688
rect 26384 13716 26390 13728
rect 28442 13716 28448 13728
rect 26384 13688 28448 13716
rect 26384 13676 26390 13688
rect 28442 13676 28448 13688
rect 28500 13716 28506 13728
rect 28718 13716 28724 13728
rect 28500 13688 28724 13716
rect 28500 13676 28506 13688
rect 28718 13676 28724 13688
rect 28776 13676 28782 13728
rect 31110 13676 31116 13728
rect 31168 13716 31174 13728
rect 36906 13716 36912 13728
rect 31168 13688 36912 13716
rect 31168 13676 31174 13688
rect 36906 13676 36912 13688
rect 36964 13676 36970 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 10686 13472 10692 13524
rect 10744 13512 10750 13524
rect 15470 13512 15476 13524
rect 10744 13484 15476 13512
rect 10744 13472 10750 13484
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 17862 13512 17868 13524
rect 17823 13484 17868 13512
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 19242 13512 19248 13524
rect 19203 13484 19248 13512
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 22833 13515 22891 13521
rect 22833 13481 22845 13515
rect 22879 13512 22891 13515
rect 22922 13512 22928 13524
rect 22879 13484 22928 13512
rect 22879 13481 22891 13484
rect 22833 13475 22891 13481
rect 22922 13472 22928 13484
rect 22980 13472 22986 13524
rect 25590 13472 25596 13524
rect 25648 13512 25654 13524
rect 26973 13515 27031 13521
rect 26973 13512 26985 13515
rect 25648 13484 26985 13512
rect 25648 13472 25654 13484
rect 26973 13481 26985 13484
rect 27019 13481 27031 13515
rect 26973 13475 27031 13481
rect 28721 13515 28779 13521
rect 28721 13481 28733 13515
rect 28767 13512 28779 13515
rect 29270 13512 29276 13524
rect 28767 13484 29276 13512
rect 28767 13481 28779 13484
rect 28721 13475 28779 13481
rect 29270 13472 29276 13484
rect 29328 13472 29334 13524
rect 29546 13512 29552 13524
rect 29507 13484 29552 13512
rect 29546 13472 29552 13484
rect 29604 13512 29610 13524
rect 30098 13512 30104 13524
rect 29604 13484 30104 13512
rect 29604 13472 29610 13484
rect 30098 13472 30104 13484
rect 30156 13472 30162 13524
rect 32033 13515 32091 13521
rect 32033 13481 32045 13515
rect 32079 13512 32091 13515
rect 32122 13512 32128 13524
rect 32079 13484 32128 13512
rect 32079 13481 32091 13484
rect 32033 13475 32091 13481
rect 32122 13472 32128 13484
rect 32180 13472 32186 13524
rect 36081 13515 36139 13521
rect 36081 13481 36093 13515
rect 36127 13512 36139 13515
rect 36170 13512 36176 13524
rect 36127 13484 36176 13512
rect 36127 13481 36139 13484
rect 36081 13475 36139 13481
rect 36170 13472 36176 13484
rect 36228 13472 36234 13524
rect 38838 13512 38844 13524
rect 38799 13484 38844 13512
rect 38838 13472 38844 13484
rect 38896 13472 38902 13524
rect 12250 13404 12256 13456
rect 12308 13444 12314 13456
rect 16025 13447 16083 13453
rect 16025 13444 16037 13447
rect 12308 13416 16037 13444
rect 12308 13404 12314 13416
rect 16025 13413 16037 13416
rect 16071 13413 16083 13447
rect 16025 13407 16083 13413
rect 14918 13376 14924 13388
rect 14568 13348 14924 13376
rect 8570 13268 8576 13320
rect 8628 13308 8634 13320
rect 9953 13311 10011 13317
rect 9953 13308 9965 13311
rect 8628 13280 9965 13308
rect 8628 13268 8634 13280
rect 9953 13277 9965 13280
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 14568 13317 14596 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 12124 13280 13369 13308
rect 12124 13268 12130 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 14415 13311 14473 13317
rect 14415 13277 14427 13311
rect 14461 13277 14473 13311
rect 14415 13271 14473 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 10220 13243 10278 13249
rect 10220 13209 10232 13243
rect 10266 13240 10278 13243
rect 10502 13240 10508 13252
rect 10266 13212 10508 13240
rect 10266 13209 10278 13212
rect 10220 13203 10278 13209
rect 10502 13200 10508 13212
rect 10560 13200 10566 13252
rect 13173 13243 13231 13249
rect 13173 13209 13185 13243
rect 13219 13240 13231 13243
rect 13262 13240 13268 13252
rect 13219 13212 13268 13240
rect 13219 13209 13231 13212
rect 13173 13203 13231 13209
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13538 13240 13544 13252
rect 13499 13212 13544 13240
rect 13538 13200 13544 13212
rect 13596 13200 13602 13252
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 12342 13172 12348 13184
rect 11379 13144 12348 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 14182 13172 14188 13184
rect 14143 13144 14188 13172
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 14430 13172 14458 13271
rect 14663 13265 14669 13317
rect 14721 13305 14727 13317
rect 14829 13311 14887 13317
rect 14721 13277 14766 13305
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15286 13308 15292 13320
rect 14875 13280 15292 13308
rect 14875 13277 14887 13280
rect 14721 13265 14727 13277
rect 14829 13271 14887 13277
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 16040 13308 16068 13407
rect 22462 13404 22468 13456
rect 22520 13444 22526 13456
rect 24670 13444 24676 13456
rect 22520 13416 24676 13444
rect 22520 13404 22526 13416
rect 24670 13404 24676 13416
rect 24728 13404 24734 13456
rect 24949 13447 25007 13453
rect 24949 13413 24961 13447
rect 24995 13444 25007 13447
rect 26234 13444 26240 13456
rect 24995 13416 26240 13444
rect 24995 13413 25007 13416
rect 24949 13407 25007 13413
rect 26234 13404 26240 13416
rect 26292 13404 26298 13456
rect 26418 13444 26424 13456
rect 26344 13416 26424 13444
rect 21450 13376 21456 13388
rect 21411 13348 21456 13376
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 26344 13376 26372 13416
rect 26418 13404 26424 13416
rect 26476 13404 26482 13456
rect 28258 13404 28264 13456
rect 28316 13444 28322 13456
rect 28316 13416 34744 13444
rect 28316 13404 28322 13416
rect 29914 13376 29920 13388
rect 26344 13348 26464 13376
rect 16577 13311 16635 13317
rect 16577 13308 16589 13311
rect 16040 13280 16589 13308
rect 16577 13277 16589 13280
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13308 19487 13311
rect 20165 13311 20223 13317
rect 20165 13308 20177 13311
rect 19475 13280 20177 13308
rect 19475 13277 19487 13280
rect 19429 13271 19487 13277
rect 20165 13277 20177 13280
rect 20211 13308 20223 13311
rect 20254 13308 20260 13320
rect 20211 13280 20260 13308
rect 20211 13277 20223 13280
rect 20165 13271 20223 13277
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13308 20407 13311
rect 20714 13308 20720 13320
rect 20395 13280 20720 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 21720 13311 21778 13317
rect 21720 13277 21732 13311
rect 21766 13308 21778 13311
rect 25774 13308 25780 13320
rect 21766 13280 25780 13308
rect 21766 13277 21778 13280
rect 21720 13271 21778 13277
rect 25774 13268 25780 13280
rect 25832 13268 25838 13320
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 26145 13311 26203 13317
rect 26145 13277 26157 13311
rect 26191 13277 26203 13311
rect 26145 13271 26203 13277
rect 26065 13256 26096 13271
rect 14918 13200 14924 13252
rect 14976 13240 14982 13252
rect 15194 13240 15200 13252
rect 14976 13212 15200 13240
rect 14976 13200 14982 13212
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 25130 13240 25136 13252
rect 25091 13212 25136 13240
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 25317 13243 25375 13249
rect 25317 13209 25329 13243
rect 25363 13240 25375 13243
rect 25682 13240 25688 13252
rect 25363 13212 25688 13240
rect 25363 13209 25375 13212
rect 25317 13203 25375 13209
rect 25682 13200 25688 13212
rect 25740 13200 25746 13252
rect 25866 13200 25872 13252
rect 25924 13240 25930 13252
rect 26065 13240 26093 13256
rect 25924 13212 26093 13240
rect 25924 13200 25930 13212
rect 15378 13172 15384 13184
rect 14430 13144 15384 13172
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 20530 13172 20536 13184
rect 20491 13144 20536 13172
rect 20530 13132 20536 13144
rect 20588 13132 20594 13184
rect 25774 13172 25780 13184
rect 25735 13144 25780 13172
rect 25774 13132 25780 13144
rect 25832 13132 25838 13184
rect 26160 13172 26188 13271
rect 26234 13268 26240 13320
rect 26292 13317 26298 13320
rect 26436 13317 26464 13348
rect 28184 13348 29920 13376
rect 26292 13308 26300 13317
rect 26433 13311 26491 13317
rect 26292 13280 26337 13308
rect 26292 13271 26300 13280
rect 26433 13277 26445 13311
rect 26479 13277 26491 13311
rect 27249 13311 27307 13317
rect 27249 13296 27261 13311
rect 27295 13296 27307 13311
rect 27341 13311 27399 13317
rect 26433 13271 26491 13277
rect 26292 13268 26298 13271
rect 27246 13244 27252 13296
rect 27304 13244 27310 13296
rect 27341 13277 27353 13311
rect 27387 13277 27399 13311
rect 27341 13271 27399 13277
rect 27154 13172 27160 13184
rect 26160 13144 27160 13172
rect 27154 13132 27160 13144
rect 27212 13172 27218 13184
rect 27356 13172 27384 13271
rect 27430 13268 27436 13320
rect 27488 13305 27494 13320
rect 27617 13311 27675 13317
rect 27488 13277 27530 13305
rect 27617 13277 27629 13311
rect 27663 13308 27675 13311
rect 28074 13308 28080 13320
rect 27663 13280 28080 13308
rect 27663 13277 27675 13280
rect 27488 13268 27494 13277
rect 27617 13271 27675 13277
rect 28074 13268 28080 13280
rect 28132 13268 28138 13320
rect 28184 13302 28212 13348
rect 29914 13336 29920 13348
rect 29972 13336 29978 13388
rect 33045 13379 33103 13385
rect 33045 13345 33057 13379
rect 33091 13376 33103 13379
rect 33134 13376 33140 13388
rect 33091 13348 33140 13376
rect 33091 13345 33103 13348
rect 33045 13339 33103 13345
rect 33134 13336 33140 13348
rect 33192 13336 33198 13388
rect 34716 13376 34744 13416
rect 39022 13404 39028 13456
rect 39080 13444 39086 13456
rect 39853 13447 39911 13453
rect 39853 13444 39865 13447
rect 39080 13416 39865 13444
rect 39080 13404 39086 13416
rect 39853 13413 39865 13416
rect 39899 13413 39911 13447
rect 39853 13407 39911 13413
rect 34716 13348 34836 13376
rect 28240 13305 28298 13311
rect 28240 13302 28252 13305
rect 28184 13274 28252 13302
rect 28240 13271 28252 13274
rect 28286 13271 28298 13305
rect 28240 13265 28298 13271
rect 28350 13268 28356 13320
rect 28408 13308 28414 13320
rect 28534 13317 28540 13320
rect 28491 13311 28540 13317
rect 28408 13280 28453 13308
rect 28408 13268 28414 13280
rect 28491 13277 28503 13311
rect 28537 13277 28540 13311
rect 28491 13271 28540 13277
rect 28534 13268 28540 13271
rect 28592 13268 28598 13320
rect 32766 13308 32772 13320
rect 32727 13280 32772 13308
rect 32766 13268 32772 13280
rect 32824 13268 32830 13320
rect 34698 13308 34704 13320
rect 34659 13280 34704 13308
rect 34698 13268 34704 13280
rect 34756 13268 34762 13320
rect 34808 13308 34836 13348
rect 36538 13336 36544 13388
rect 36596 13376 36602 13388
rect 37090 13376 37096 13388
rect 36596 13348 37096 13376
rect 36596 13336 36602 13348
rect 37090 13336 37096 13348
rect 37148 13376 37154 13388
rect 37148 13348 37504 13376
rect 37148 13336 37154 13348
rect 37476 13317 37504 13348
rect 37369 13311 37427 13317
rect 34808 13280 36676 13308
rect 30098 13200 30104 13252
rect 30156 13240 30162 13252
rect 33502 13240 33508 13252
rect 30156 13212 33508 13240
rect 30156 13200 30162 13212
rect 33502 13200 33508 13212
rect 33560 13240 33566 13252
rect 34422 13240 34428 13252
rect 33560 13212 34428 13240
rect 33560 13200 33566 13212
rect 34422 13200 34428 13212
rect 34480 13200 34486 13252
rect 34790 13200 34796 13252
rect 34848 13240 34854 13252
rect 36648 13249 36676 13280
rect 37369 13277 37381 13311
rect 37415 13277 37427 13311
rect 37369 13271 37427 13277
rect 37461 13311 37519 13317
rect 37461 13277 37473 13311
rect 37507 13277 37519 13311
rect 37461 13271 37519 13277
rect 37553 13311 37611 13317
rect 37553 13277 37565 13311
rect 37599 13308 37611 13311
rect 37642 13308 37648 13320
rect 37599 13280 37648 13308
rect 37599 13277 37611 13280
rect 37553 13271 37611 13277
rect 34946 13243 35004 13249
rect 34946 13240 34958 13243
rect 34848 13212 34958 13240
rect 34848 13200 34854 13212
rect 34946 13209 34958 13212
rect 34992 13209 35004 13243
rect 34946 13203 35004 13209
rect 36633 13243 36691 13249
rect 36633 13209 36645 13243
rect 36679 13240 36691 13243
rect 37384 13240 37412 13271
rect 37642 13268 37648 13280
rect 37700 13268 37706 13320
rect 37734 13268 37740 13320
rect 37792 13308 37798 13320
rect 38194 13308 38200 13320
rect 37792 13280 37837 13308
rect 38155 13280 38200 13308
rect 37792 13268 37798 13280
rect 38194 13268 38200 13280
rect 38252 13268 38258 13320
rect 38378 13308 38384 13320
rect 38339 13280 38384 13308
rect 38378 13268 38384 13280
rect 38436 13268 38442 13320
rect 38473 13311 38531 13317
rect 38473 13277 38485 13311
rect 38519 13277 38531 13311
rect 38473 13271 38531 13277
rect 36679 13212 37492 13240
rect 36679 13209 36691 13212
rect 36633 13203 36691 13209
rect 37090 13172 37096 13184
rect 27212 13144 27384 13172
rect 37051 13144 37096 13172
rect 27212 13132 27218 13144
rect 37090 13132 37096 13144
rect 37148 13132 37154 13184
rect 37464 13172 37492 13212
rect 38286 13200 38292 13252
rect 38344 13240 38350 13252
rect 38488 13240 38516 13271
rect 38562 13268 38568 13320
rect 38620 13308 38626 13320
rect 40037 13311 40095 13317
rect 38620 13280 38665 13308
rect 38620 13268 38626 13280
rect 40037 13277 40049 13311
rect 40083 13308 40095 13311
rect 40218 13308 40224 13320
rect 40083 13280 40224 13308
rect 40083 13277 40095 13280
rect 40037 13271 40095 13277
rect 40218 13268 40224 13280
rect 40276 13268 40282 13320
rect 58158 13308 58164 13320
rect 58119 13280 58164 13308
rect 58158 13268 58164 13280
rect 58216 13268 58222 13320
rect 38344 13212 38516 13240
rect 38344 13200 38350 13212
rect 39114 13172 39120 13184
rect 37464 13144 39120 13172
rect 39114 13132 39120 13144
rect 39172 13132 39178 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 3329 12971 3387 12977
rect 3329 12937 3341 12971
rect 3375 12968 3387 12971
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 3375 12940 4261 12968
rect 3375 12937 3387 12940
rect 3329 12931 3387 12937
rect 4249 12937 4261 12940
rect 4295 12968 4307 12971
rect 4890 12968 4896 12980
rect 4295 12940 4896 12968
rect 4295 12937 4307 12940
rect 4249 12931 4307 12937
rect 4890 12928 4896 12940
rect 4948 12968 4954 12980
rect 5258 12968 5264 12980
rect 4948 12940 5264 12968
rect 4948 12928 4954 12940
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 11790 12968 11796 12980
rect 11751 12940 11796 12968
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 13262 12928 13268 12980
rect 13320 12968 13326 12980
rect 21269 12971 21327 12977
rect 13320 12940 15700 12968
rect 13320 12928 13326 12940
rect 12928 12903 12986 12909
rect 12928 12869 12940 12903
rect 12974 12900 12986 12903
rect 14182 12900 14188 12912
rect 12974 12872 14188 12900
rect 12974 12869 12986 12872
rect 12928 12863 12986 12869
rect 14182 12860 14188 12872
rect 14240 12860 14246 12912
rect 15470 12900 15476 12912
rect 15431 12872 15476 12900
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 15672 12909 15700 12940
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 21726 12968 21732 12980
rect 21315 12940 21732 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 15657 12903 15715 12909
rect 15657 12869 15669 12903
rect 15703 12900 15715 12903
rect 16666 12900 16672 12912
rect 15703 12872 16672 12900
rect 15703 12869 15715 12872
rect 15657 12863 15715 12869
rect 16666 12860 16672 12872
rect 16724 12860 16730 12912
rect 17862 12860 17868 12912
rect 17920 12900 17926 12912
rect 17920 12872 18092 12900
rect 17920 12860 17926 12872
rect 14645 12844 14703 12847
rect 18064 12844 18092 12872
rect 2130 12832 2136 12844
rect 2091 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2363 12804 3004 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2314 12656 2320 12708
rect 2372 12696 2378 12708
rect 2976 12705 3004 12804
rect 7374 12792 7380 12844
rect 7432 12832 7438 12844
rect 7846 12835 7904 12841
rect 7846 12832 7858 12835
rect 7432 12804 7858 12832
rect 7432 12792 7438 12804
rect 7846 12801 7858 12804
rect 7892 12801 7904 12835
rect 7846 12795 7904 12801
rect 8840 12835 8898 12841
rect 8840 12801 8852 12835
rect 8886 12832 8898 12835
rect 9122 12832 9128 12844
rect 8886 12804 9128 12832
rect 8886 12801 8898 12804
rect 8840 12795 8898 12801
rect 9122 12792 9128 12804
rect 9180 12792 9186 12844
rect 14366 12792 14372 12844
rect 14424 12841 14430 12844
rect 14424 12835 14473 12841
rect 14424 12801 14427 12835
rect 14461 12801 14473 12835
rect 14424 12795 14473 12801
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 14424 12792 14430 12795
rect 3418 12764 3424 12776
rect 3379 12736 3424 12764
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 3602 12764 3608 12776
rect 3563 12736 3608 12764
rect 3602 12724 3608 12736
rect 3660 12764 3666 12776
rect 3878 12764 3884 12776
rect 3660 12736 3884 12764
rect 3660 12724 3666 12736
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 8110 12764 8116 12776
rect 8071 12736 8116 12764
rect 8110 12724 8116 12736
rect 8168 12764 8174 12776
rect 8570 12764 8576 12776
rect 8168 12736 8576 12764
rect 8168 12724 8174 12736
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 14090 12764 14096 12776
rect 13219 12736 14096 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 14090 12724 14096 12736
rect 14148 12724 14154 12776
rect 14568 12764 14596 12795
rect 14642 12792 14648 12844
rect 14700 12838 14706 12844
rect 14700 12810 14739 12838
rect 14829 12835 14887 12841
rect 14700 12792 14706 12810
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15286 12832 15292 12844
rect 14875 12804 15292 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 17782 12835 17840 12841
rect 17782 12832 17794 12835
rect 17552 12804 17794 12832
rect 17552 12792 17558 12804
rect 17782 12801 17794 12804
rect 17828 12801 17840 12835
rect 18046 12832 18052 12844
rect 17959 12804 18052 12832
rect 17782 12795 17840 12801
rect 18046 12792 18052 12804
rect 18104 12792 18110 12844
rect 20162 12792 20168 12844
rect 20220 12832 20226 12844
rect 20303 12835 20361 12841
rect 20303 12832 20315 12835
rect 20220 12804 20315 12832
rect 20220 12792 20226 12804
rect 20303 12801 20315 12804
rect 20349 12801 20361 12835
rect 20438 12832 20444 12844
rect 20399 12804 20444 12832
rect 20303 12795 20361 12801
rect 20438 12792 20444 12804
rect 20496 12792 20502 12844
rect 20530 12792 20536 12844
rect 20588 12832 20594 12844
rect 20717 12835 20775 12841
rect 20588 12804 20633 12832
rect 20588 12792 20594 12804
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 21284 12832 21312 12931
rect 21726 12928 21732 12940
rect 21784 12928 21790 12980
rect 24949 12971 25007 12977
rect 24949 12937 24961 12971
rect 24995 12968 25007 12971
rect 25130 12968 25136 12980
rect 24995 12940 25136 12968
rect 24995 12937 25007 12940
rect 24949 12931 25007 12937
rect 25130 12928 25136 12940
rect 25188 12928 25194 12980
rect 27985 12971 28043 12977
rect 27985 12937 27997 12971
rect 28031 12968 28043 12971
rect 28074 12968 28080 12980
rect 28031 12940 28080 12968
rect 28031 12937 28043 12940
rect 27985 12931 28043 12937
rect 28074 12928 28080 12940
rect 28132 12968 28138 12980
rect 28534 12968 28540 12980
rect 28132 12940 28540 12968
rect 28132 12928 28138 12940
rect 28534 12928 28540 12940
rect 28592 12928 28598 12980
rect 31570 12968 31576 12980
rect 31531 12940 31576 12968
rect 31570 12928 31576 12940
rect 31628 12928 31634 12980
rect 32766 12928 32772 12980
rect 32824 12968 32830 12980
rect 33042 12968 33048 12980
rect 32824 12940 33048 12968
rect 32824 12928 32830 12940
rect 33042 12928 33048 12940
rect 33100 12968 33106 12980
rect 33229 12971 33287 12977
rect 33229 12968 33241 12971
rect 33100 12940 33241 12968
rect 33100 12928 33106 12940
rect 33229 12937 33241 12940
rect 33275 12937 33287 12971
rect 37642 12968 37648 12980
rect 37603 12940 37648 12968
rect 33229 12931 33287 12937
rect 37642 12928 37648 12940
rect 37700 12928 37706 12980
rect 25774 12860 25780 12912
rect 25832 12900 25838 12912
rect 26062 12903 26120 12909
rect 26062 12900 26074 12903
rect 25832 12872 26074 12900
rect 25832 12860 25838 12872
rect 26062 12869 26074 12872
rect 26108 12869 26120 12903
rect 26062 12863 26120 12869
rect 28997 12903 29055 12909
rect 28997 12869 29009 12903
rect 29043 12900 29055 12903
rect 31110 12900 31116 12912
rect 29043 12872 31116 12900
rect 29043 12869 29055 12872
rect 28997 12863 29055 12869
rect 26326 12832 26332 12844
rect 20763 12804 21312 12832
rect 26287 12804 26332 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 29748 12841 29776 12872
rect 31110 12860 31116 12872
rect 31168 12860 31174 12912
rect 31297 12903 31355 12909
rect 31297 12869 31309 12903
rect 31343 12900 31355 12903
rect 31846 12900 31852 12912
rect 31343 12872 31852 12900
rect 31343 12869 31355 12872
rect 31297 12863 31355 12869
rect 31846 12860 31852 12872
rect 31904 12860 31910 12912
rect 31938 12860 31944 12912
rect 31996 12900 32002 12912
rect 32306 12900 32312 12912
rect 31996 12872 32312 12900
rect 31996 12860 32002 12872
rect 32306 12860 32312 12872
rect 32364 12900 32370 12912
rect 32364 12872 32536 12900
rect 32364 12860 32370 12872
rect 29733 12835 29791 12841
rect 29733 12801 29745 12835
rect 29779 12801 29791 12835
rect 29733 12795 29791 12801
rect 29825 12835 29883 12841
rect 29825 12801 29837 12835
rect 29871 12801 29883 12835
rect 29825 12795 29883 12801
rect 19153 12767 19211 12773
rect 14568 12736 15056 12764
rect 15028 12708 15056 12736
rect 19153 12733 19165 12767
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 19429 12767 19487 12773
rect 19429 12733 19441 12767
rect 19475 12764 19487 12767
rect 20456 12764 20484 12792
rect 19475 12736 20484 12764
rect 19475 12733 19487 12736
rect 19429 12727 19487 12733
rect 2961 12699 3019 12705
rect 2372 12668 2774 12696
rect 2372 12656 2378 12668
rect 2406 12588 2412 12640
rect 2464 12628 2470 12640
rect 2501 12631 2559 12637
rect 2501 12628 2513 12631
rect 2464 12600 2513 12628
rect 2464 12588 2470 12600
rect 2501 12597 2513 12600
rect 2547 12597 2559 12631
rect 2746 12628 2774 12668
rect 2961 12665 2973 12699
rect 3007 12665 3019 12699
rect 6733 12699 6791 12705
rect 6733 12696 6745 12699
rect 2961 12659 3019 12665
rect 4080 12668 6745 12696
rect 4080 12628 4108 12668
rect 6733 12665 6745 12668
rect 6779 12696 6791 12699
rect 7006 12696 7012 12708
rect 6779 12668 7012 12696
rect 6779 12665 6791 12668
rect 6733 12659 6791 12665
rect 7006 12656 7012 12668
rect 7064 12656 7070 12708
rect 13998 12656 14004 12708
rect 14056 12696 14062 12708
rect 14185 12699 14243 12705
rect 14185 12696 14197 12699
rect 14056 12668 14197 12696
rect 14056 12656 14062 12668
rect 14185 12665 14197 12668
rect 14231 12665 14243 12699
rect 14185 12659 14243 12665
rect 15010 12656 15016 12708
rect 15068 12696 15074 12708
rect 15194 12696 15200 12708
rect 15068 12668 15200 12696
rect 15068 12656 15074 12668
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 16669 12699 16727 12705
rect 16669 12665 16681 12699
rect 16715 12665 16727 12699
rect 16669 12659 16727 12665
rect 2746 12600 4108 12628
rect 9953 12631 10011 12637
rect 2501 12591 2559 12597
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10962 12628 10968 12640
rect 9999 12600 10968 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 10962 12588 10968 12600
rect 11020 12588 11026 12640
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15160 12600 15301 12628
rect 15160 12588 15166 12600
rect 15289 12597 15301 12600
rect 15335 12597 15347 12631
rect 16684 12628 16712 12659
rect 17310 12628 17316 12640
rect 16684 12600 17316 12628
rect 15289 12591 15347 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 17678 12588 17684 12640
rect 17736 12628 17742 12640
rect 19168 12628 19196 12727
rect 29362 12724 29368 12776
rect 29420 12764 29426 12776
rect 29840 12764 29868 12795
rect 29914 12792 29920 12844
rect 29972 12832 29978 12844
rect 30101 12835 30159 12841
rect 29972 12804 30017 12832
rect 29972 12792 29978 12804
rect 30101 12801 30113 12835
rect 30147 12832 30159 12835
rect 30374 12832 30380 12844
rect 30147 12804 30380 12832
rect 30147 12801 30159 12804
rect 30101 12795 30159 12801
rect 30374 12792 30380 12804
rect 30432 12792 30438 12844
rect 30926 12792 30932 12844
rect 30984 12832 30990 12844
rect 31021 12835 31079 12841
rect 31021 12832 31033 12835
rect 30984 12804 31033 12832
rect 30984 12792 30990 12804
rect 31021 12801 31033 12804
rect 31067 12801 31079 12835
rect 31202 12832 31208 12844
rect 31163 12804 31208 12832
rect 31021 12795 31079 12801
rect 31202 12792 31208 12804
rect 31260 12792 31266 12844
rect 31386 12792 31392 12844
rect 31444 12832 31450 12844
rect 31444 12804 31489 12832
rect 31444 12792 31450 12804
rect 32122 12792 32128 12844
rect 32180 12832 32186 12844
rect 32508 12841 32536 12872
rect 37090 12860 37096 12912
rect 37148 12900 37154 12912
rect 39678 12903 39736 12909
rect 39678 12900 39690 12903
rect 37148 12872 39690 12900
rect 37148 12860 37154 12872
rect 39678 12869 39690 12872
rect 39724 12869 39736 12903
rect 39678 12863 39736 12869
rect 32401 12835 32459 12841
rect 32401 12832 32413 12835
rect 32180 12804 32413 12832
rect 32180 12792 32186 12804
rect 32401 12801 32413 12804
rect 32447 12801 32459 12835
rect 32401 12795 32459 12801
rect 32493 12835 32551 12841
rect 32493 12801 32505 12835
rect 32539 12801 32551 12835
rect 32493 12795 32551 12801
rect 32582 12792 32588 12844
rect 32640 12832 32646 12844
rect 32769 12835 32827 12841
rect 32640 12804 32685 12832
rect 32640 12792 32646 12804
rect 32769 12801 32781 12835
rect 32815 12832 32827 12835
rect 32858 12832 32864 12844
rect 32815 12804 32864 12832
rect 32815 12801 32827 12804
rect 32769 12795 32827 12801
rect 29420 12736 29868 12764
rect 29420 12724 29426 12736
rect 30374 12656 30380 12708
rect 30432 12696 30438 12708
rect 32784 12696 32812 12795
rect 32858 12792 32864 12804
rect 32916 12792 32922 12844
rect 35802 12832 35808 12844
rect 35763 12804 35808 12832
rect 35802 12792 35808 12804
rect 35860 12792 35866 12844
rect 36262 12792 36268 12844
rect 36320 12832 36326 12844
rect 36814 12832 36820 12844
rect 36320 12804 36820 12832
rect 36320 12792 36326 12804
rect 36814 12792 36820 12804
rect 36872 12832 36878 12844
rect 37277 12835 37335 12841
rect 37277 12832 37289 12835
rect 36872 12804 37289 12832
rect 36872 12792 36878 12804
rect 37277 12801 37289 12804
rect 37323 12801 37335 12835
rect 37277 12795 37335 12801
rect 37461 12835 37519 12841
rect 37461 12801 37473 12835
rect 37507 12832 37519 12835
rect 37550 12832 37556 12844
rect 37507 12804 37556 12832
rect 37507 12801 37519 12804
rect 37461 12795 37519 12801
rect 37550 12792 37556 12804
rect 37608 12792 37614 12844
rect 39945 12835 40003 12841
rect 39945 12801 39957 12835
rect 39991 12832 40003 12835
rect 40034 12832 40040 12844
rect 39991 12804 40040 12832
rect 39991 12801 40003 12804
rect 39945 12795 40003 12801
rect 40034 12792 40040 12804
rect 40092 12792 40098 12844
rect 35529 12767 35587 12773
rect 35529 12733 35541 12767
rect 35575 12764 35587 12767
rect 35618 12764 35624 12776
rect 35575 12736 35624 12764
rect 35575 12733 35587 12736
rect 35529 12727 35587 12733
rect 35618 12724 35624 12736
rect 35676 12724 35682 12776
rect 30432 12668 32812 12696
rect 37568 12696 37596 12792
rect 38565 12699 38623 12705
rect 38565 12696 38577 12699
rect 37568 12668 38577 12696
rect 30432 12656 30438 12668
rect 38565 12665 38577 12668
rect 38611 12665 38623 12699
rect 38565 12659 38623 12665
rect 20070 12628 20076 12640
rect 17736 12600 19196 12628
rect 20031 12600 20076 12628
rect 17736 12588 17742 12600
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 27065 12631 27123 12637
rect 27065 12597 27077 12631
rect 27111 12628 27123 12631
rect 27246 12628 27252 12640
rect 27111 12600 27252 12628
rect 27111 12597 27123 12600
rect 27065 12591 27123 12597
rect 27246 12588 27252 12600
rect 27304 12588 27310 12640
rect 29454 12628 29460 12640
rect 29415 12600 29460 12628
rect 29454 12588 29460 12600
rect 29512 12588 29518 12640
rect 32125 12631 32183 12637
rect 32125 12597 32137 12631
rect 32171 12628 32183 12631
rect 32582 12628 32588 12640
rect 32171 12600 32588 12628
rect 32171 12597 32183 12600
rect 32125 12591 32183 12597
rect 32582 12588 32588 12600
rect 32640 12588 32646 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 10502 12424 10508 12436
rect 5868 12396 5948 12424
rect 10463 12396 10508 12424
rect 5868 12384 5874 12396
rect 3237 12359 3295 12365
rect 3237 12325 3249 12359
rect 3283 12325 3295 12359
rect 3237 12319 3295 12325
rect 3252 12288 3280 12319
rect 3418 12288 3424 12300
rect 3252 12260 3424 12288
rect 3418 12248 3424 12260
rect 3476 12288 3482 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 3476 12260 5733 12288
rect 3476 12248 3482 12260
rect 5721 12257 5733 12260
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 5920 12232 5948 12396
rect 10502 12384 10508 12396
rect 10560 12384 10566 12436
rect 15470 12424 15476 12436
rect 13924 12396 15056 12424
rect 15431 12396 15476 12424
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 7929 12359 7987 12365
rect 7929 12356 7941 12359
rect 6972 12328 7941 12356
rect 6972 12316 6978 12328
rect 7929 12325 7941 12328
rect 7975 12356 7987 12359
rect 8110 12356 8116 12368
rect 7975 12328 8116 12356
rect 7975 12325 7987 12328
rect 7929 12319 7987 12325
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 9766 12316 9772 12368
rect 9824 12316 9830 12368
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 9784 12288 9812 12316
rect 10137 12291 10195 12297
rect 10137 12288 10149 12291
rect 8536 12260 10149 12288
rect 8536 12248 8542 12260
rect 10137 12257 10149 12260
rect 10183 12257 10195 12291
rect 11057 12291 11115 12297
rect 11057 12288 11069 12291
rect 10137 12251 10195 12257
rect 10244 12260 11069 12288
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 3142 12220 3148 12232
rect 1903 12192 3148 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 5810 12220 5816 12232
rect 5771 12192 5816 12220
rect 5810 12180 5816 12192
rect 5868 12180 5874 12232
rect 5902 12180 5908 12232
rect 5960 12180 5966 12232
rect 5994 12180 6000 12232
rect 6052 12220 6058 12232
rect 6454 12220 6460 12232
rect 6052 12192 6460 12220
rect 6052 12180 6058 12192
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 8386 12180 8392 12232
rect 8444 12220 8450 12232
rect 9398 12220 9404 12232
rect 8444 12192 9404 12220
rect 8444 12180 8450 12192
rect 9398 12180 9404 12192
rect 9456 12220 9462 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9456 12192 9781 12220
rect 9456 12180 9462 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 9769 12183 9827 12189
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12189 10011 12223
rect 9953 12183 10011 12189
rect 2124 12155 2182 12161
rect 2124 12121 2136 12155
rect 2170 12152 2182 12155
rect 2222 12152 2228 12164
rect 2170 12124 2228 12152
rect 2170 12121 2182 12124
rect 2124 12115 2182 12121
rect 2222 12112 2228 12124
rect 2280 12112 2286 12164
rect 5442 12112 5448 12164
rect 5500 12152 5506 12164
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 5500 12124 6653 12152
rect 5500 12112 5506 12124
rect 6641 12121 6653 12124
rect 6687 12121 6699 12155
rect 9968 12152 9996 12183
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10100 12192 10145 12220
rect 10100 12180 10106 12192
rect 10244 12152 10272 12260
rect 11057 12257 11069 12260
rect 11103 12288 11115 12291
rect 13924 12288 13952 12396
rect 15028 12356 15056 12396
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 17494 12424 17500 12436
rect 17455 12396 17500 12424
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 17586 12384 17592 12436
rect 17644 12424 17650 12436
rect 20530 12424 20536 12436
rect 17644 12396 20536 12424
rect 17644 12384 17650 12396
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21177 12427 21235 12433
rect 21177 12424 21189 12427
rect 20772 12396 21189 12424
rect 20772 12384 20778 12396
rect 21177 12393 21189 12396
rect 21223 12393 21235 12427
rect 29914 12424 29920 12436
rect 29875 12396 29920 12424
rect 21177 12387 21235 12393
rect 29914 12384 29920 12396
rect 29972 12384 29978 12436
rect 34422 12384 34428 12436
rect 34480 12424 34486 12436
rect 35894 12424 35900 12436
rect 34480 12396 35900 12424
rect 34480 12384 34486 12396
rect 35894 12384 35900 12396
rect 35952 12384 35958 12436
rect 36354 12424 36360 12436
rect 36315 12396 36360 12424
rect 36354 12384 36360 12396
rect 36412 12424 36418 12436
rect 37182 12424 37188 12436
rect 36412 12396 37188 12424
rect 36412 12384 36418 12396
rect 37182 12384 37188 12396
rect 37240 12384 37246 12436
rect 18414 12356 18420 12368
rect 15028 12328 18420 12356
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 22741 12359 22799 12365
rect 22741 12325 22753 12359
rect 22787 12356 22799 12359
rect 23014 12356 23020 12368
rect 22787 12328 23020 12356
rect 22787 12325 22799 12328
rect 22741 12319 22799 12325
rect 23014 12316 23020 12328
rect 23072 12356 23078 12368
rect 24394 12356 24400 12368
rect 23072 12328 24400 12356
rect 23072 12316 23078 12328
rect 24394 12316 24400 12328
rect 24452 12316 24458 12368
rect 31389 12359 31447 12365
rect 31389 12325 31401 12359
rect 31435 12356 31447 12359
rect 32214 12356 32220 12368
rect 31435 12328 32220 12356
rect 31435 12325 31447 12328
rect 31389 12319 31447 12325
rect 32214 12316 32220 12328
rect 32272 12316 32278 12368
rect 35526 12356 35532 12368
rect 34992 12328 35532 12356
rect 11103 12260 13952 12288
rect 11103 12257 11115 12260
rect 11057 12251 11115 12257
rect 17678 12248 17684 12300
rect 17736 12288 17742 12300
rect 17736 12260 17908 12288
rect 17736 12248 17742 12260
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 11422 12220 11428 12232
rect 10367 12192 11428 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 11790 12180 11796 12232
rect 11848 12220 11854 12232
rect 13173 12223 13231 12229
rect 11848 12192 12434 12220
rect 11848 12180 11854 12192
rect 12250 12152 12256 12164
rect 9968 12124 10272 12152
rect 11072 12124 12256 12152
rect 6641 12115 6699 12121
rect 5353 12087 5411 12093
rect 5353 12053 5365 12087
rect 5399 12084 5411 12087
rect 5718 12084 5724 12096
rect 5399 12056 5724 12084
rect 5399 12053 5411 12056
rect 5353 12047 5411 12053
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6656 12084 6684 12115
rect 11072 12096 11100 12124
rect 12250 12112 12256 12124
rect 12308 12112 12314 12164
rect 12406 12152 12434 12192
rect 13173 12189 13185 12223
rect 13219 12220 13231 12223
rect 13262 12220 13268 12232
rect 13219 12192 13268 12220
rect 13219 12189 13231 12192
rect 13173 12183 13231 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 14090 12220 14096 12232
rect 14051 12192 14096 12220
rect 14090 12180 14096 12192
rect 14148 12180 14154 12232
rect 14734 12220 14740 12232
rect 14200 12192 14740 12220
rect 13357 12155 13415 12161
rect 13357 12152 13369 12155
rect 12406 12124 13369 12152
rect 13357 12121 13369 12124
rect 13403 12121 13415 12155
rect 13357 12115 13415 12121
rect 13541 12155 13599 12161
rect 13541 12121 13553 12155
rect 13587 12152 13599 12155
rect 14200 12152 14228 12192
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 17586 12220 17592 12232
rect 15304 12192 17592 12220
rect 13587 12124 14228 12152
rect 14360 12155 14418 12161
rect 13587 12121 13599 12124
rect 13541 12115 13599 12121
rect 14360 12121 14372 12155
rect 14406 12152 14418 12155
rect 14642 12152 14648 12164
rect 14406 12124 14648 12152
rect 14406 12121 14418 12124
rect 14360 12115 14418 12121
rect 14642 12112 14648 12124
rect 14700 12112 14706 12164
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 6656 12056 8953 12084
rect 8941 12053 8953 12056
rect 8987 12084 8999 12087
rect 11054 12084 11060 12096
rect 8987 12056 11060 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11422 12044 11428 12096
rect 11480 12084 11486 12096
rect 12342 12084 12348 12096
rect 11480 12056 12348 12084
rect 11480 12044 11486 12056
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12986 12044 12992 12096
rect 13044 12084 13050 12096
rect 15304 12084 15332 12192
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17880 12229 17908 12260
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 18104 12260 19809 12288
rect 18104 12248 18110 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 22830 12248 22836 12300
rect 22888 12288 22894 12300
rect 27338 12288 27344 12300
rect 22888 12260 27344 12288
rect 22888 12248 22894 12260
rect 27338 12248 27344 12260
rect 27396 12288 27402 12300
rect 33229 12291 33287 12297
rect 27396 12260 31754 12288
rect 27396 12248 27402 12260
rect 17773 12223 17831 12229
rect 17773 12189 17785 12223
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 16666 12152 16672 12164
rect 16627 12124 16672 12152
rect 16666 12112 16672 12124
rect 16724 12112 16730 12164
rect 16853 12155 16911 12161
rect 16853 12121 16865 12155
rect 16899 12121 16911 12155
rect 17788 12152 17816 12183
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18141 12223 18199 12229
rect 18012 12192 18057 12220
rect 18012 12180 18018 12192
rect 18141 12189 18153 12223
rect 18187 12220 18199 12223
rect 18690 12220 18696 12232
rect 18187 12192 18696 12220
rect 18187 12189 18199 12192
rect 18141 12183 18199 12189
rect 18690 12180 18696 12192
rect 18748 12180 18754 12232
rect 20070 12229 20076 12232
rect 20064 12183 20076 12229
rect 20128 12220 20134 12232
rect 20128 12192 20164 12220
rect 20070 12180 20076 12183
rect 20128 12180 20134 12192
rect 27614 12180 27620 12232
rect 27672 12220 27678 12232
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 27672 12192 29745 12220
rect 27672 12180 27678 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 30834 12220 30840 12232
rect 30795 12192 30840 12220
rect 29733 12183 29791 12189
rect 30834 12180 30840 12192
rect 30892 12180 30898 12232
rect 31205 12223 31263 12229
rect 31205 12189 31217 12223
rect 31251 12220 31263 12223
rect 31386 12220 31392 12232
rect 31251 12192 31392 12220
rect 31251 12189 31263 12192
rect 31205 12183 31263 12189
rect 31386 12180 31392 12192
rect 31444 12180 31450 12232
rect 31726 12220 31754 12260
rect 33229 12257 33241 12291
rect 33275 12288 33287 12291
rect 34698 12288 34704 12300
rect 33275 12260 34704 12288
rect 33275 12257 33287 12260
rect 33229 12251 33287 12257
rect 34698 12248 34704 12260
rect 34756 12248 34762 12300
rect 31726 12192 32536 12220
rect 19337 12155 19395 12161
rect 19337 12152 19349 12155
rect 17788 12124 19349 12152
rect 16853 12115 16911 12121
rect 19337 12121 19349 12124
rect 19383 12152 19395 12155
rect 19426 12152 19432 12164
rect 19383 12124 19432 12152
rect 19383 12121 19395 12124
rect 19337 12115 19395 12121
rect 13044 12056 15332 12084
rect 13044 12044 13050 12056
rect 15838 12044 15844 12096
rect 15896 12084 15902 12096
rect 16482 12084 16488 12096
rect 15896 12056 16488 12084
rect 15896 12044 15902 12056
rect 16482 12044 16488 12056
rect 16540 12084 16546 12096
rect 16868 12084 16896 12115
rect 19426 12112 19432 12124
rect 19484 12112 19490 12164
rect 20530 12112 20536 12164
rect 20588 12152 20594 12164
rect 22005 12155 22063 12161
rect 22005 12152 22017 12155
rect 20588 12124 22017 12152
rect 20588 12112 20594 12124
rect 22005 12121 22017 12124
rect 22051 12152 22063 12155
rect 22557 12155 22615 12161
rect 22557 12152 22569 12155
rect 22051 12124 22569 12152
rect 22051 12121 22063 12124
rect 22005 12115 22063 12121
rect 22557 12121 22569 12124
rect 22603 12152 22615 12155
rect 28810 12152 28816 12164
rect 22603 12124 28816 12152
rect 22603 12121 22615 12124
rect 22557 12115 22615 12121
rect 28810 12112 28816 12124
rect 28868 12112 28874 12164
rect 29549 12155 29607 12161
rect 29549 12121 29561 12155
rect 29595 12152 29607 12155
rect 30466 12152 30472 12164
rect 29595 12124 30472 12152
rect 29595 12121 29607 12124
rect 29549 12115 29607 12121
rect 30466 12112 30472 12124
rect 30524 12152 30530 12164
rect 30742 12152 30748 12164
rect 30524 12124 30748 12152
rect 30524 12112 30530 12124
rect 30742 12112 30748 12124
rect 30800 12112 30806 12164
rect 31021 12155 31079 12161
rect 31021 12121 31033 12155
rect 31067 12121 31079 12155
rect 31021 12115 31079 12121
rect 31113 12155 31171 12161
rect 31113 12121 31125 12155
rect 31159 12152 31171 12155
rect 32030 12152 32036 12164
rect 31159 12124 32036 12152
rect 31159 12121 31171 12124
rect 31113 12115 31171 12121
rect 16540 12056 16896 12084
rect 17037 12087 17095 12093
rect 16540 12044 16546 12056
rect 17037 12053 17049 12087
rect 17083 12084 17095 12087
rect 17954 12084 17960 12096
rect 17083 12056 17960 12084
rect 17083 12053 17095 12056
rect 17037 12047 17095 12053
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 18690 12084 18696 12096
rect 18603 12056 18696 12084
rect 18690 12044 18696 12056
rect 18748 12084 18754 12096
rect 20438 12084 20444 12096
rect 18748 12056 20444 12084
rect 18748 12044 18754 12056
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 25682 12084 25688 12096
rect 25643 12056 25688 12084
rect 25682 12044 25688 12056
rect 25740 12044 25746 12096
rect 31036 12084 31064 12115
rect 32030 12112 32036 12124
rect 32088 12112 32094 12164
rect 31202 12084 31208 12096
rect 31036 12056 31208 12084
rect 31202 12044 31208 12056
rect 31260 12044 31266 12096
rect 31846 12084 31852 12096
rect 31807 12056 31852 12084
rect 31846 12044 31852 12056
rect 31904 12044 31910 12096
rect 32508 12084 32536 12192
rect 32582 12180 32588 12232
rect 32640 12220 32646 12232
rect 34992 12229 35020 12328
rect 35526 12316 35532 12328
rect 35584 12316 35590 12368
rect 35434 12288 35440 12300
rect 35084 12260 35440 12288
rect 35084 12229 35112 12260
rect 35434 12248 35440 12260
rect 35492 12248 35498 12300
rect 32962 12223 33020 12229
rect 32962 12220 32974 12223
rect 32640 12192 32974 12220
rect 32640 12180 32646 12192
rect 32962 12189 32974 12192
rect 33008 12189 33020 12223
rect 32962 12183 33020 12189
rect 34149 12223 34207 12229
rect 34149 12189 34161 12223
rect 34195 12220 34207 12223
rect 34977 12223 35035 12229
rect 34977 12220 34989 12223
rect 34195 12192 34989 12220
rect 34195 12189 34207 12192
rect 34149 12183 34207 12189
rect 34977 12189 34989 12192
rect 35023 12189 35035 12223
rect 34977 12183 35035 12189
rect 35069 12223 35127 12229
rect 35069 12189 35081 12223
rect 35115 12189 35127 12223
rect 35069 12183 35127 12189
rect 35161 12223 35219 12229
rect 35161 12189 35173 12223
rect 35207 12220 35219 12223
rect 35250 12220 35256 12232
rect 35207 12192 35256 12220
rect 35207 12189 35219 12192
rect 35161 12183 35219 12189
rect 35250 12180 35256 12192
rect 35308 12180 35314 12232
rect 35345 12223 35403 12229
rect 35345 12189 35357 12223
rect 35391 12220 35403 12223
rect 35618 12220 35624 12232
rect 35391 12192 35624 12220
rect 35391 12189 35403 12192
rect 35345 12183 35403 12189
rect 35618 12180 35624 12192
rect 35676 12180 35682 12232
rect 34701 12155 34759 12161
rect 34701 12121 34713 12155
rect 34747 12152 34759 12155
rect 34790 12152 34796 12164
rect 34747 12124 34796 12152
rect 34747 12121 34759 12124
rect 34701 12115 34759 12121
rect 34790 12112 34796 12124
rect 34848 12112 34854 12164
rect 34882 12112 34888 12164
rect 34940 12152 34946 12164
rect 36265 12155 36323 12161
rect 36265 12152 36277 12155
rect 34940 12124 36277 12152
rect 34940 12112 34946 12124
rect 36265 12121 36277 12124
rect 36311 12121 36323 12155
rect 36265 12115 36323 12121
rect 38013 12087 38071 12093
rect 38013 12084 38025 12087
rect 32508 12056 38025 12084
rect 38013 12053 38025 12056
rect 38059 12084 38071 12087
rect 38562 12084 38568 12096
rect 38059 12056 38568 12084
rect 38059 12053 38071 12056
rect 38013 12047 38071 12053
rect 38562 12044 38568 12056
rect 38620 12044 38626 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 2222 11880 2228 11892
rect 2183 11852 2228 11880
rect 2222 11840 2228 11852
rect 2280 11840 2286 11892
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 6914 11880 6920 11892
rect 3200 11852 6920 11880
rect 3200 11840 3206 11852
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7193 11883 7251 11889
rect 7193 11849 7205 11883
rect 7239 11880 7251 11883
rect 7374 11880 7380 11892
rect 7239 11852 7380 11880
rect 7239 11849 7251 11852
rect 7193 11843 7251 11849
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 9122 11880 9128 11892
rect 9083 11852 9128 11880
rect 9122 11840 9128 11852
rect 9180 11840 9186 11892
rect 11701 11883 11759 11889
rect 11701 11849 11713 11883
rect 11747 11880 11759 11883
rect 12986 11880 12992 11892
rect 11747 11852 12992 11880
rect 11747 11849 11759 11852
rect 11701 11843 11759 11849
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 14642 11880 14648 11892
rect 14603 11852 14648 11880
rect 14642 11840 14648 11852
rect 14700 11840 14706 11892
rect 15010 11880 15016 11892
rect 15009 11840 15016 11880
rect 15068 11840 15074 11892
rect 16482 11840 16488 11892
rect 16540 11880 16546 11892
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 16540 11852 16681 11880
rect 16540 11840 16546 11852
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 17678 11880 17684 11892
rect 16669 11843 16727 11849
rect 16776 11852 17684 11880
rect 8478 11772 8484 11824
rect 8536 11812 8542 11824
rect 8536 11784 8800 11812
rect 8536 11772 8542 11784
rect 2406 11744 2412 11756
rect 2367 11716 2412 11744
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 3234 11704 3240 11756
rect 3292 11744 3298 11756
rect 3401 11747 3459 11753
rect 3401 11744 3413 11747
rect 3292 11716 3413 11744
rect 3292 11704 3298 11716
rect 3401 11713 3413 11716
rect 3447 11713 3459 11747
rect 3401 11707 3459 11713
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 3142 11676 3148 11688
rect 3103 11648 3148 11676
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 4614 11568 4620 11620
rect 4672 11608 4678 11620
rect 5350 11608 5356 11620
rect 4672 11580 5356 11608
rect 4672 11568 4678 11580
rect 5350 11568 5356 11580
rect 5408 11608 5414 11620
rect 5537 11611 5595 11617
rect 5537 11608 5549 11611
rect 5408 11580 5549 11608
rect 5408 11568 5414 11580
rect 5537 11577 5549 11580
rect 5583 11577 5595 11611
rect 5736 11608 5764 11707
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 6420 11716 6469 11744
rect 6420 11704 6426 11716
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6638 11744 6644 11756
rect 6599 11716 6644 11744
rect 6457 11707 6515 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 7006 11744 7012 11756
rect 6967 11716 7012 11744
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 8386 11744 8392 11756
rect 8347 11716 8392 11744
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 8772 11753 8800 11784
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 8496 11716 8585 11744
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 6052 11648 6745 11676
rect 6052 11636 6058 11648
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7282 11676 7288 11688
rect 6871 11648 7288 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7374 11608 7380 11620
rect 5736 11580 7380 11608
rect 5537 11571 5595 11577
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 8496 11608 8524 11716
rect 8573 11713 8585 11716
rect 8619 11713 8631 11747
rect 8573 11707 8631 11713
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11744 8999 11747
rect 10962 11744 10968 11756
rect 8987 11716 10968 11744
rect 8987 11713 8999 11716
rect 8941 11707 8999 11713
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11514 11744 11520 11756
rect 11475 11716 11520 11744
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 15009 11753 15037 11840
rect 15194 11772 15200 11824
rect 15252 11812 15258 11824
rect 16776 11812 16804 11852
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 19613 11883 19671 11889
rect 19613 11849 19625 11883
rect 19659 11880 19671 11883
rect 20162 11880 20168 11892
rect 19659 11852 20168 11880
rect 19659 11849 19671 11852
rect 19613 11843 19671 11849
rect 20162 11840 20168 11852
rect 20220 11880 20226 11892
rect 22830 11880 22836 11892
rect 20220 11852 22836 11880
rect 20220 11840 20226 11852
rect 22830 11840 22836 11852
rect 22888 11840 22894 11892
rect 23106 11840 23112 11892
rect 23164 11880 23170 11892
rect 24486 11880 24492 11892
rect 23164 11852 24492 11880
rect 23164 11840 23170 11852
rect 24486 11840 24492 11852
rect 24544 11840 24550 11892
rect 27249 11883 27307 11889
rect 27249 11849 27261 11883
rect 27295 11880 27307 11883
rect 27614 11880 27620 11892
rect 27295 11852 27620 11880
rect 27295 11849 27307 11852
rect 27249 11843 27307 11849
rect 27614 11840 27620 11852
rect 27672 11840 27678 11892
rect 28626 11880 28632 11892
rect 27724 11852 28632 11880
rect 15252 11784 16804 11812
rect 15252 11772 15258 11784
rect 17218 11772 17224 11824
rect 17276 11812 17282 11824
rect 17862 11812 17868 11824
rect 17276 11784 17868 11812
rect 17276 11772 17282 11784
rect 17862 11772 17868 11784
rect 17920 11812 17926 11824
rect 17920 11784 18092 11812
rect 17920 11772 17926 11784
rect 14875 11747 14933 11753
rect 14875 11713 14887 11747
rect 14921 11713 14933 11747
rect 14875 11707 14933 11713
rect 14994 11747 15052 11753
rect 14994 11713 15006 11747
rect 15040 11713 15052 11747
rect 14994 11707 15052 11713
rect 15094 11747 15152 11753
rect 15094 11713 15106 11747
rect 15140 11713 15152 11747
rect 15094 11707 15152 11713
rect 8662 11676 8668 11688
rect 8623 11648 8668 11676
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 14734 11676 14740 11688
rect 9723 11648 14740 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 9692 11608 9720 11639
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 8496 11580 9720 11608
rect 4525 11543 4583 11549
rect 4525 11509 4537 11543
rect 4571 11540 4583 11543
rect 5626 11540 5632 11552
rect 4571 11512 5632 11540
rect 4571 11509 4583 11512
rect 4525 11503 4583 11509
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 5994 11500 6000 11552
rect 6052 11540 6058 11552
rect 6362 11540 6368 11552
rect 6052 11512 6368 11540
rect 6052 11500 6058 11512
rect 6362 11500 6368 11512
rect 6420 11540 6426 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 6420 11512 7757 11540
rect 6420 11500 6426 11512
rect 7745 11509 7757 11512
rect 7791 11540 7803 11543
rect 7926 11540 7932 11552
rect 7791 11512 7932 11540
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 14890 11540 14918 11707
rect 15120 11676 15148 11707
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15344 11716 15389 11744
rect 15344 11704 15350 11716
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 18064 11753 18092 11784
rect 20438 11772 20444 11824
rect 20496 11812 20502 11824
rect 25961 11815 26019 11821
rect 25961 11812 25973 11815
rect 20496 11784 25973 11812
rect 20496 11772 20502 11784
rect 25961 11781 25973 11784
rect 26007 11812 26019 11815
rect 27724 11812 27752 11852
rect 28626 11840 28632 11852
rect 28684 11840 28690 11892
rect 31478 11880 31484 11892
rect 31036 11852 31484 11880
rect 26007 11784 27752 11812
rect 28384 11815 28442 11821
rect 26007 11781 26019 11784
rect 25961 11775 26019 11781
rect 28384 11781 28396 11815
rect 28430 11812 28442 11815
rect 29454 11812 29460 11824
rect 28430 11784 29460 11812
rect 28430 11781 28442 11784
rect 28384 11775 28442 11781
rect 29454 11772 29460 11784
rect 29512 11772 29518 11824
rect 17782 11747 17840 11753
rect 17782 11744 17794 11747
rect 17552 11716 17794 11744
rect 17552 11704 17558 11716
rect 17782 11713 17794 11716
rect 17828 11713 17840 11747
rect 17782 11707 17840 11713
rect 18049 11747 18107 11753
rect 18049 11713 18061 11747
rect 18095 11713 18107 11747
rect 18874 11744 18880 11756
rect 18787 11716 18880 11744
rect 18049 11707 18107 11713
rect 18874 11704 18880 11716
rect 18932 11744 18938 11756
rect 19521 11747 19579 11753
rect 19521 11744 19533 11747
rect 18932 11716 19533 11744
rect 18932 11704 18938 11716
rect 19521 11713 19533 11716
rect 19567 11713 19579 11747
rect 22554 11744 22560 11756
rect 22515 11716 22560 11744
rect 19521 11707 19579 11713
rect 22554 11704 22560 11716
rect 22612 11704 22618 11756
rect 22741 11747 22799 11753
rect 22741 11713 22753 11747
rect 22787 11744 22799 11747
rect 23474 11744 23480 11756
rect 22787 11716 23480 11744
rect 22787 11713 22799 11716
rect 22741 11707 22799 11713
rect 23474 11704 23480 11716
rect 23532 11704 23538 11756
rect 24949 11747 25007 11753
rect 24949 11713 24961 11747
rect 24995 11744 25007 11747
rect 25774 11744 25780 11756
rect 24995 11716 25780 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 25774 11704 25780 11716
rect 25832 11704 25838 11756
rect 28629 11747 28687 11753
rect 28629 11713 28641 11747
rect 28675 11744 28687 11747
rect 28718 11744 28724 11756
rect 28675 11716 28724 11744
rect 28675 11713 28687 11716
rect 28629 11707 28687 11713
rect 28718 11704 28724 11716
rect 28776 11704 28782 11756
rect 31036 11753 31064 11852
rect 31478 11840 31484 11852
rect 31536 11840 31542 11892
rect 31573 11883 31631 11889
rect 31573 11849 31585 11883
rect 31619 11880 31631 11883
rect 31754 11880 31760 11892
rect 31619 11852 31760 11880
rect 31619 11849 31631 11852
rect 31573 11843 31631 11849
rect 31754 11840 31760 11852
rect 31812 11840 31818 11892
rect 31294 11812 31300 11824
rect 31255 11784 31300 11812
rect 31294 11772 31300 11784
rect 31352 11772 31358 11824
rect 31021 11747 31079 11753
rect 31021 11713 31033 11747
rect 31067 11713 31079 11747
rect 31202 11744 31208 11756
rect 31163 11716 31208 11744
rect 31021 11707 31079 11713
rect 31202 11704 31208 11716
rect 31260 11704 31266 11756
rect 31386 11744 31392 11756
rect 31347 11716 31392 11744
rect 31386 11704 31392 11716
rect 31444 11704 31450 11756
rect 32766 11744 32772 11756
rect 32679 11716 32772 11744
rect 32766 11704 32772 11716
rect 32824 11744 32830 11756
rect 34882 11744 34888 11756
rect 32824 11716 34888 11744
rect 32824 11704 32830 11716
rect 34882 11704 34888 11716
rect 34940 11704 34946 11756
rect 36078 11744 36084 11756
rect 36039 11716 36084 11744
rect 36078 11704 36084 11716
rect 36136 11704 36142 11756
rect 38286 11704 38292 11756
rect 38344 11744 38350 11756
rect 38473 11747 38531 11753
rect 38473 11744 38485 11747
rect 38344 11716 38485 11744
rect 38344 11704 38350 11716
rect 38473 11713 38485 11716
rect 38519 11713 38531 11747
rect 38473 11707 38531 11713
rect 15194 11676 15200 11688
rect 15120 11648 15200 11676
rect 15194 11636 15200 11648
rect 15252 11636 15258 11688
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 15068 11580 16574 11608
rect 15068 11568 15074 11580
rect 15562 11540 15568 11552
rect 14890 11512 15568 11540
rect 15562 11500 15568 11512
rect 15620 11540 15626 11552
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 15620 11512 15761 11540
rect 15620 11500 15626 11512
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 16546 11540 16574 11580
rect 18322 11540 18328 11552
rect 16546 11512 18328 11540
rect 15749 11503 15807 11509
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 18414 11500 18420 11552
rect 18472 11540 18478 11552
rect 18892 11549 18920 11704
rect 28810 11636 28816 11688
rect 28868 11676 28874 11688
rect 32493 11679 32551 11685
rect 32493 11676 32505 11679
rect 28868 11648 32505 11676
rect 28868 11636 28874 11648
rect 32493 11645 32505 11648
rect 32539 11676 32551 11679
rect 33042 11676 33048 11688
rect 32539 11648 33048 11676
rect 32539 11645 32551 11648
rect 32493 11639 32551 11645
rect 33042 11636 33048 11648
rect 33100 11676 33106 11688
rect 33781 11679 33839 11685
rect 33781 11676 33793 11679
rect 33100 11648 33793 11676
rect 33100 11636 33106 11648
rect 33781 11645 33793 11648
rect 33827 11645 33839 11679
rect 33781 11639 33839 11645
rect 37734 11636 37740 11688
rect 37792 11676 37798 11688
rect 38197 11679 38255 11685
rect 38197 11676 38209 11679
rect 37792 11648 38209 11676
rect 37792 11636 37798 11648
rect 38197 11645 38209 11648
rect 38243 11676 38255 11679
rect 38930 11676 38936 11688
rect 38243 11648 38936 11676
rect 38243 11645 38255 11648
rect 38197 11639 38255 11645
rect 38930 11636 38936 11648
rect 38988 11636 38994 11688
rect 23382 11568 23388 11620
rect 23440 11608 23446 11620
rect 24765 11611 24823 11617
rect 24765 11608 24777 11611
rect 23440 11580 24777 11608
rect 23440 11568 23446 11580
rect 24765 11577 24777 11580
rect 24811 11577 24823 11611
rect 58158 11608 58164 11620
rect 58119 11580 58164 11608
rect 24765 11571 24823 11577
rect 58158 11568 58164 11580
rect 58216 11568 58222 11620
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18472 11512 18889 11540
rect 18472 11500 18478 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 22373 11543 22431 11549
rect 22373 11509 22385 11543
rect 22419 11540 22431 11543
rect 23014 11540 23020 11552
rect 22419 11512 23020 11540
rect 22419 11509 22431 11512
rect 22373 11503 22431 11509
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 35342 11500 35348 11552
rect 35400 11540 35406 11552
rect 36265 11543 36323 11549
rect 36265 11540 36277 11543
rect 35400 11512 36277 11540
rect 35400 11500 35406 11512
rect 36265 11509 36277 11512
rect 36311 11540 36323 11543
rect 37274 11540 37280 11552
rect 36311 11512 37280 11540
rect 36311 11509 36323 11512
rect 36265 11503 36323 11509
rect 37274 11500 37280 11512
rect 37332 11500 37338 11552
rect 39025 11543 39083 11549
rect 39025 11509 39037 11543
rect 39071 11540 39083 11543
rect 39114 11540 39120 11552
rect 39071 11512 39120 11540
rect 39071 11509 39083 11512
rect 39025 11503 39083 11509
rect 39114 11500 39120 11512
rect 39172 11500 39178 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 3234 11336 3240 11348
rect 3195 11308 3240 11336
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 7009 11339 7067 11345
rect 7009 11305 7021 11339
rect 7055 11336 7067 11339
rect 8662 11336 8668 11348
rect 7055 11308 8668 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 14090 11296 14096 11348
rect 14148 11336 14154 11348
rect 17218 11336 17224 11348
rect 14148 11308 17224 11336
rect 14148 11296 14154 11308
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 17494 11336 17500 11348
rect 17455 11308 17500 11336
rect 17494 11296 17500 11308
rect 17552 11296 17558 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 24394 11336 24400 11348
rect 22428 11308 24256 11336
rect 24355 11308 24400 11336
rect 22428 11296 22434 11308
rect 11146 11268 11152 11280
rect 11107 11240 11152 11268
rect 11146 11228 11152 11240
rect 11204 11268 11210 11280
rect 11204 11240 12434 11268
rect 11204 11228 11210 11240
rect 4614 11200 4620 11212
rect 4575 11172 4620 11200
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5626 11200 5632 11212
rect 5587 11172 5632 11200
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11200 5871 11203
rect 5902 11200 5908 11212
rect 5859 11172 5908 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 6144 11172 6377 11200
rect 6144 11160 6150 11172
rect 6365 11169 6377 11172
rect 6411 11169 6423 11203
rect 6365 11163 6423 11169
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 6696 11172 7481 11200
rect 6696 11160 6702 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 12406 11200 12434 11240
rect 15286 11228 15292 11280
rect 15344 11268 15350 11280
rect 15344 11240 18000 11268
rect 15344 11228 15350 11240
rect 16942 11200 16948 11212
rect 12406 11172 16948 11200
rect 7469 11163 7527 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17678 11160 17684 11212
rect 17736 11200 17742 11212
rect 17972 11200 18000 11240
rect 22922 11228 22928 11280
rect 22980 11228 22986 11280
rect 24228 11268 24256 11308
rect 24394 11296 24400 11308
rect 24452 11296 24458 11348
rect 26694 11296 26700 11348
rect 26752 11336 26758 11348
rect 26789 11339 26847 11345
rect 26789 11336 26801 11339
rect 26752 11308 26801 11336
rect 26752 11296 26758 11308
rect 26789 11305 26801 11308
rect 26835 11305 26847 11339
rect 26789 11299 26847 11305
rect 29549 11339 29607 11345
rect 29549 11305 29561 11339
rect 29595 11336 29607 11339
rect 29730 11336 29736 11348
rect 29595 11308 29736 11336
rect 29595 11305 29607 11308
rect 29549 11299 29607 11305
rect 29730 11296 29736 11308
rect 29788 11296 29794 11348
rect 32033 11339 32091 11345
rect 32033 11305 32045 11339
rect 32079 11336 32091 11339
rect 32490 11336 32496 11348
rect 32079 11308 32496 11336
rect 32079 11305 32091 11308
rect 32033 11299 32091 11305
rect 32490 11296 32496 11308
rect 32548 11296 32554 11348
rect 35894 11336 35900 11348
rect 35855 11308 35900 11336
rect 35894 11296 35900 11308
rect 35952 11296 35958 11348
rect 28445 11271 28503 11277
rect 28445 11268 28457 11271
rect 24228 11240 28457 11268
rect 28445 11237 28457 11240
rect 28491 11268 28503 11271
rect 28626 11268 28632 11280
rect 28491 11240 28632 11268
rect 28491 11237 28503 11240
rect 28445 11231 28503 11237
rect 28626 11228 28632 11240
rect 28684 11228 28690 11280
rect 28736 11240 32812 11268
rect 22646 11200 22652 11212
rect 17736 11172 17908 11200
rect 17972 11172 22652 11200
rect 17736 11160 17742 11172
rect 3050 11132 3056 11144
rect 3011 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 5644 11132 5672 11160
rect 6733 11135 6791 11141
rect 6733 11132 6745 11135
rect 5644 11104 6745 11132
rect 4341 11095 4399 11101
rect 6733 11101 6745 11104
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 4356 11064 4384 11095
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 6880 11104 6925 11132
rect 6880 11092 6886 11104
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12492 11104 12537 11132
rect 12492 11092 12498 11104
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 17880 11141 17908 11172
rect 22646 11160 22652 11172
rect 22704 11160 22710 11212
rect 17773 11135 17831 11141
rect 12676 11104 12721 11132
rect 12676 11092 12682 11104
rect 17773 11101 17785 11135
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11101 17923 11135
rect 17865 11095 17923 11101
rect 4614 11064 4620 11076
rect 4356 11036 4620 11064
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 5534 11064 5540 11076
rect 5495 11036 5540 11064
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 5776 11036 6960 11064
rect 5776 11024 5782 11036
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 5169 10999 5227 11005
rect 5169 10996 5181 10999
rect 4304 10968 5181 10996
rect 4304 10956 4310 10968
rect 5169 10965 5181 10968
rect 5215 10965 5227 10999
rect 6932 10996 6960 11036
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 10965 11067 11023 11073
rect 10965 11064 10977 11067
rect 7432 11036 10977 11064
rect 7432 11024 7438 11036
rect 10965 11033 10977 11036
rect 11011 11064 11023 11067
rect 11514 11064 11520 11076
rect 11011 11036 11520 11064
rect 11011 11033 11023 11036
rect 10965 11027 11023 11033
rect 11514 11024 11520 11036
rect 11572 11024 11578 11076
rect 17788 11064 17816 11095
rect 17954 11092 17960 11144
rect 18012 11132 18018 11144
rect 18141 11135 18199 11141
rect 18012 11104 18057 11132
rect 18012 11092 18018 11104
rect 18141 11101 18153 11135
rect 18187 11132 18199 11135
rect 18690 11132 18696 11144
rect 18187 11104 18696 11132
rect 18187 11101 18199 11104
rect 18141 11095 18199 11101
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11132 22155 11135
rect 22830 11132 22836 11144
rect 22143 11104 22836 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 22830 11092 22836 11104
rect 22888 11092 22894 11144
rect 22940 11141 22968 11228
rect 22922 11135 22980 11141
rect 22922 11101 22934 11135
rect 22968 11101 22980 11135
rect 22922 11095 22980 11101
rect 23014 11092 23020 11144
rect 23072 11141 23078 11144
rect 23072 11132 23080 11141
rect 23213 11135 23271 11141
rect 23072 11104 23117 11132
rect 23072 11095 23080 11104
rect 23213 11101 23225 11135
rect 23259 11132 23271 11135
rect 23382 11132 23388 11144
rect 23259 11104 23388 11132
rect 23259 11101 23271 11104
rect 23213 11095 23271 11101
rect 23072 11092 23078 11095
rect 23382 11092 23388 11104
rect 23440 11092 23446 11144
rect 25774 11092 25780 11144
rect 25832 11132 25838 11144
rect 26881 11135 26939 11141
rect 26881 11132 26893 11135
rect 25832 11104 26893 11132
rect 25832 11092 25838 11104
rect 26881 11101 26893 11104
rect 26927 11132 26939 11135
rect 28736 11132 28764 11240
rect 32784 11212 32812 11240
rect 34698 11228 34704 11280
rect 34756 11268 34762 11280
rect 36354 11268 36360 11280
rect 34756 11240 36360 11268
rect 34756 11228 34762 11240
rect 36354 11228 36360 11240
rect 36412 11268 36418 11280
rect 37737 11271 37795 11277
rect 37737 11268 37749 11271
rect 36412 11240 37749 11268
rect 36412 11228 36418 11240
rect 37737 11237 37749 11240
rect 37783 11268 37795 11271
rect 38562 11268 38568 11280
rect 37783 11240 38568 11268
rect 37783 11237 37795 11240
rect 37737 11231 37795 11237
rect 38562 11228 38568 11240
rect 38620 11228 38626 11280
rect 32766 11200 32772 11212
rect 29472 11172 30144 11200
rect 32727 11172 32772 11200
rect 29472 11144 29500 11172
rect 26927 11104 28764 11132
rect 28997 11135 29055 11141
rect 26927 11101 26939 11104
rect 26881 11095 26939 11101
rect 28997 11101 29009 11135
rect 29043 11132 29055 11135
rect 29454 11132 29460 11144
rect 29043 11104 29460 11132
rect 29043 11101 29055 11104
rect 28997 11095 29055 11101
rect 29454 11092 29460 11104
rect 29512 11092 29518 11144
rect 29730 11132 29736 11144
rect 29691 11104 29736 11132
rect 29730 11092 29736 11104
rect 29788 11092 29794 11144
rect 30116 11141 30144 11172
rect 32766 11160 32772 11172
rect 32824 11160 32830 11212
rect 32858 11160 32864 11212
rect 32916 11200 32922 11212
rect 33045 11203 33103 11209
rect 33045 11200 33057 11203
rect 32916 11172 33057 11200
rect 32916 11160 32922 11172
rect 33045 11169 33057 11172
rect 33091 11169 33103 11203
rect 33045 11163 33103 11169
rect 30101 11135 30159 11141
rect 30101 11101 30113 11135
rect 30147 11101 30159 11135
rect 31846 11132 31852 11144
rect 31807 11104 31852 11132
rect 30101 11095 30159 11101
rect 31846 11092 31852 11104
rect 31904 11092 31910 11144
rect 35069 11135 35127 11141
rect 35069 11101 35081 11135
rect 35115 11132 35127 11135
rect 35115 11104 35388 11132
rect 35115 11101 35127 11104
rect 35069 11095 35127 11101
rect 18506 11064 18512 11076
rect 17788 11036 18512 11064
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 28718 11024 28724 11076
rect 28776 11064 28782 11076
rect 29825 11067 29883 11073
rect 29825 11064 29837 11067
rect 28776 11036 29837 11064
rect 28776 11024 28782 11036
rect 29825 11033 29837 11036
rect 29871 11033 29883 11067
rect 29825 11027 29883 11033
rect 29917 11067 29975 11073
rect 29917 11033 29929 11067
rect 29963 11064 29975 11067
rect 30374 11064 30380 11076
rect 29963 11036 30380 11064
rect 29963 11033 29975 11036
rect 29917 11027 29975 11033
rect 30374 11024 30380 11036
rect 30432 11024 30438 11076
rect 30466 11024 30472 11076
rect 30524 11064 30530 11076
rect 31570 11064 31576 11076
rect 30524 11036 31576 11064
rect 30524 11024 30530 11036
rect 31570 11024 31576 11036
rect 31628 11064 31634 11076
rect 31665 11067 31723 11073
rect 31665 11064 31677 11067
rect 31628 11036 31677 11064
rect 31628 11024 31634 11036
rect 31665 11033 31677 11036
rect 31711 11033 31723 11067
rect 35250 11064 35256 11076
rect 35211 11036 35256 11064
rect 31665 11027 31723 11033
rect 35250 11024 35256 11036
rect 35308 11024 35314 11076
rect 35360 11064 35388 11104
rect 35894 11092 35900 11144
rect 35952 11132 35958 11144
rect 36449 11135 36507 11141
rect 36449 11132 36461 11135
rect 35952 11104 36461 11132
rect 35952 11092 35958 11104
rect 36449 11101 36461 11104
rect 36495 11101 36507 11135
rect 36449 11095 36507 11101
rect 37182 11092 37188 11144
rect 37240 11132 37246 11144
rect 38657 11135 38715 11141
rect 38657 11132 38669 11135
rect 37240 11104 38669 11132
rect 37240 11092 37246 11104
rect 38657 11101 38669 11104
rect 38703 11101 38715 11135
rect 38820 11135 38878 11141
rect 38820 11132 38832 11135
rect 38657 11095 38715 11101
rect 38764 11104 38832 11132
rect 35360 11036 35940 11064
rect 35912 11008 35940 11036
rect 37642 11024 37648 11076
rect 37700 11064 37706 11076
rect 38764 11064 38792 11104
rect 38820 11101 38832 11104
rect 38866 11101 38878 11135
rect 38820 11095 38878 11101
rect 38930 11092 38936 11144
rect 38988 11132 38994 11144
rect 39114 11141 39120 11144
rect 39071 11135 39120 11141
rect 38988 11104 39033 11132
rect 38988 11092 38994 11104
rect 39071 11101 39083 11135
rect 39117 11101 39120 11135
rect 39071 11095 39120 11101
rect 39114 11092 39120 11095
rect 39172 11092 39178 11144
rect 37700 11036 38792 11064
rect 37700 11024 37706 11036
rect 7190 10996 7196 11008
rect 6932 10968 7196 10996
rect 5169 10959 5227 10965
rect 7190 10956 7196 10968
rect 7248 10956 7254 11008
rect 11606 10956 11612 11008
rect 11664 10996 11670 11008
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 11664 10968 12265 10996
rect 11664 10956 11670 10968
rect 12253 10965 12265 10968
rect 12299 10965 12311 10999
rect 12253 10959 12311 10965
rect 22278 10956 22284 11008
rect 22336 10996 22342 11008
rect 22557 10999 22615 11005
rect 22557 10996 22569 10999
rect 22336 10968 22569 10996
rect 22336 10956 22342 10968
rect 22557 10965 22569 10968
rect 22603 10965 22615 10999
rect 22557 10959 22615 10965
rect 34885 10999 34943 11005
rect 34885 10965 34897 10999
rect 34931 10996 34943 10999
rect 35434 10996 35440 11008
rect 34931 10968 35440 10996
rect 34931 10965 34943 10968
rect 34885 10959 34943 10965
rect 35434 10956 35440 10968
rect 35492 10956 35498 11008
rect 35894 10956 35900 11008
rect 35952 10956 35958 11008
rect 39298 10996 39304 11008
rect 39259 10968 39304 10996
rect 39298 10956 39304 10968
rect 39356 10956 39362 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 3050 10752 3056 10804
rect 3108 10792 3114 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 3108 10764 4077 10792
rect 3108 10752 3114 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 12345 10795 12403 10801
rect 12345 10761 12357 10795
rect 12391 10792 12403 10795
rect 12434 10792 12440 10804
rect 12391 10764 12440 10792
rect 12391 10761 12403 10764
rect 12345 10755 12403 10761
rect 12434 10752 12440 10764
rect 12492 10752 12498 10804
rect 22373 10795 22431 10801
rect 22373 10761 22385 10795
rect 22419 10792 22431 10795
rect 22462 10792 22468 10804
rect 22419 10764 22468 10792
rect 22419 10761 22431 10764
rect 22373 10755 22431 10761
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 23569 10795 23627 10801
rect 23569 10792 23581 10795
rect 23532 10764 23581 10792
rect 23532 10752 23538 10764
rect 23569 10761 23581 10764
rect 23615 10792 23627 10795
rect 24762 10792 24768 10804
rect 23615 10764 24768 10792
rect 23615 10761 23627 10764
rect 23569 10755 23627 10761
rect 24762 10752 24768 10764
rect 24820 10752 24826 10804
rect 27614 10752 27620 10804
rect 27672 10752 27678 10804
rect 28169 10795 28227 10801
rect 28169 10761 28181 10795
rect 28215 10792 28227 10795
rect 29178 10792 29184 10804
rect 28215 10764 29184 10792
rect 28215 10761 28227 10764
rect 28169 10755 28227 10761
rect 29178 10752 29184 10764
rect 29236 10752 29242 10804
rect 30098 10792 30104 10804
rect 30059 10764 30104 10792
rect 30098 10752 30104 10764
rect 30156 10792 30162 10804
rect 31018 10792 31024 10804
rect 30156 10764 31024 10792
rect 30156 10752 30162 10764
rect 31018 10752 31024 10764
rect 31076 10752 31082 10804
rect 32306 10752 32312 10804
rect 32364 10792 32370 10804
rect 37642 10792 37648 10804
rect 32364 10764 32444 10792
rect 37603 10764 37648 10792
rect 32364 10752 32370 10764
rect 5902 10684 5908 10736
rect 5960 10724 5966 10736
rect 12805 10727 12863 10733
rect 5960 10696 7696 10724
rect 5960 10684 5966 10696
rect 4246 10656 4252 10668
rect 4207 10628 4252 10656
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6641 10659 6699 10665
rect 6641 10656 6653 10659
rect 5868 10628 6653 10656
rect 5868 10616 5874 10628
rect 6641 10625 6653 10628
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 4614 10588 4620 10600
rect 4479 10560 4620 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 6362 10588 6368 10600
rect 6323 10560 6368 10588
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 7668 10597 7696 10696
rect 12805 10693 12817 10727
rect 12851 10724 12863 10727
rect 13170 10724 13176 10736
rect 12851 10696 13176 10724
rect 12851 10693 12863 10696
rect 12805 10687 12863 10693
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 20441 10727 20499 10733
rect 20441 10693 20453 10727
rect 20487 10724 20499 10727
rect 21082 10724 21088 10736
rect 20487 10696 21088 10724
rect 20487 10693 20499 10696
rect 20441 10687 20499 10693
rect 21082 10684 21088 10696
rect 21140 10684 21146 10736
rect 22097 10727 22155 10733
rect 22097 10693 22109 10727
rect 22143 10724 22155 10727
rect 22554 10724 22560 10736
rect 22143 10696 22560 10724
rect 22143 10693 22155 10696
rect 22097 10687 22155 10693
rect 22554 10684 22560 10696
rect 22612 10684 22618 10736
rect 27632 10724 27660 10752
rect 27893 10727 27951 10733
rect 27893 10724 27905 10727
rect 27632 10696 27905 10724
rect 27893 10693 27905 10696
rect 27939 10693 27951 10727
rect 28626 10724 28632 10736
rect 28587 10696 28632 10724
rect 27893 10687 27951 10693
rect 28626 10684 28632 10696
rect 28684 10684 28690 10736
rect 30374 10684 30380 10736
rect 30432 10724 30438 10736
rect 31202 10724 31208 10736
rect 30432 10696 31208 10724
rect 30432 10684 30438 10696
rect 31202 10684 31208 10696
rect 31260 10684 31266 10736
rect 32416 10671 32444 10764
rect 37642 10752 37648 10764
rect 37700 10752 37706 10804
rect 34698 10684 34704 10736
rect 34756 10684 34762 10736
rect 38562 10684 38568 10736
rect 38620 10724 38626 10736
rect 38620 10696 39896 10724
rect 38620 10684 38626 10696
rect 7834 10656 7840 10668
rect 7795 10628 7840 10656
rect 7834 10616 7840 10628
rect 7892 10616 7898 10668
rect 11606 10656 11612 10668
rect 11567 10628 11612 10656
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12710 10656 12716 10668
rect 12623 10628 12716 10656
rect 12710 10616 12716 10628
rect 12768 10656 12774 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 12768 10628 13553 10656
rect 12768 10616 12774 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 18874 10656 18880 10668
rect 17184 10628 18880 10656
rect 17184 10616 17190 10628
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 20070 10656 20076 10668
rect 19751 10628 20076 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 20070 10616 20076 10628
rect 20128 10656 20134 10668
rect 20257 10659 20315 10665
rect 20257 10656 20269 10659
rect 20128 10628 20269 10656
rect 20128 10616 20134 10628
rect 20257 10625 20269 10628
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 21821 10659 21879 10665
rect 21821 10625 21833 10659
rect 21867 10625 21879 10659
rect 22002 10656 22008 10668
rect 21963 10628 22008 10656
rect 21821 10619 21879 10625
rect 7653 10591 7711 10597
rect 7653 10557 7665 10591
rect 7699 10588 7711 10591
rect 9582 10588 9588 10600
rect 7699 10560 9588 10588
rect 7699 10557 7711 10560
rect 7653 10551 7711 10557
rect 9582 10548 9588 10560
rect 9640 10588 9646 10600
rect 12526 10588 12532 10600
rect 9640 10560 12532 10588
rect 9640 10548 9646 10560
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 11793 10523 11851 10529
rect 11793 10489 11805 10523
rect 11839 10520 11851 10523
rect 12544 10520 12572 10548
rect 12912 10520 12940 10551
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 21836 10588 21864 10619
rect 22002 10616 22008 10628
rect 22060 10616 22066 10668
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 23290 10656 23296 10668
rect 22235 10628 23296 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 23290 10616 23296 10628
rect 23348 10616 23354 10668
rect 23753 10659 23811 10665
rect 23753 10625 23765 10659
rect 23799 10656 23811 10659
rect 24026 10656 24032 10668
rect 23799 10628 24032 10656
rect 23799 10625 23811 10628
rect 23753 10619 23811 10625
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 24394 10656 24400 10668
rect 24355 10628 24400 10656
rect 24394 10616 24400 10628
rect 24452 10616 24458 10668
rect 27614 10656 27620 10668
rect 27575 10628 27620 10656
rect 27614 10616 27620 10628
rect 27672 10616 27678 10668
rect 27801 10659 27859 10665
rect 27801 10625 27813 10659
rect 27847 10625 27859 10659
rect 27801 10619 27859 10625
rect 27985 10659 28043 10665
rect 27985 10625 27997 10659
rect 28031 10656 28043 10659
rect 29546 10656 29552 10668
rect 28031 10628 29552 10656
rect 28031 10625 28043 10628
rect 27985 10619 28043 10625
rect 18656 10560 21864 10588
rect 18656 10548 18662 10560
rect 21910 10548 21916 10600
rect 21968 10588 21974 10600
rect 23017 10591 23075 10597
rect 23017 10588 23029 10591
rect 21968 10560 23029 10588
rect 21968 10548 21974 10560
rect 23017 10557 23029 10560
rect 23063 10588 23075 10591
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 23063 10560 23949 10588
rect 23063 10557 23075 10560
rect 23017 10551 23075 10557
rect 23937 10557 23949 10560
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 24673 10591 24731 10597
rect 24673 10557 24685 10591
rect 24719 10588 24731 10591
rect 25222 10588 25228 10600
rect 24719 10560 25228 10588
rect 24719 10557 24731 10560
rect 24673 10551 24731 10557
rect 25222 10548 25228 10560
rect 25280 10548 25286 10600
rect 27816 10588 27844 10619
rect 27890 10588 27896 10600
rect 27816 10560 27896 10588
rect 27890 10548 27896 10560
rect 27948 10548 27954 10600
rect 11839 10492 12434 10520
rect 12544 10492 12940 10520
rect 19061 10523 19119 10529
rect 11839 10489 11851 10492
rect 11793 10483 11851 10489
rect 12406 10464 12434 10492
rect 19061 10489 19073 10523
rect 19107 10520 19119 10523
rect 19107 10492 22094 10520
rect 19107 10489 19119 10492
rect 19061 10483 19119 10489
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10452 8907 10455
rect 9306 10452 9312 10464
rect 8895 10424 9312 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 12406 10424 12440 10464
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 18325 10455 18383 10461
rect 18325 10421 18337 10455
rect 18371 10452 18383 10455
rect 18506 10452 18512 10464
rect 18371 10424 18512 10452
rect 18371 10421 18383 10424
rect 18325 10415 18383 10421
rect 18506 10412 18512 10424
rect 18564 10412 18570 10464
rect 22066 10452 22094 10492
rect 23290 10480 23296 10532
rect 23348 10520 23354 10532
rect 28000 10520 28028 10619
rect 29546 10616 29552 10628
rect 29604 10616 29610 10668
rect 29730 10616 29736 10668
rect 29788 10656 29794 10668
rect 31021 10659 31079 10665
rect 31021 10656 31033 10659
rect 29788 10628 31033 10656
rect 29788 10616 29794 10628
rect 31021 10625 31033 10628
rect 31067 10625 31079 10659
rect 31021 10619 31079 10625
rect 31036 10588 31064 10619
rect 31110 10616 31116 10668
rect 31168 10656 31174 10668
rect 31389 10659 31447 10665
rect 31168 10628 31213 10656
rect 31168 10616 31174 10628
rect 31389 10625 31401 10659
rect 31435 10625 31447 10659
rect 31389 10619 31447 10625
rect 32125 10659 32183 10665
rect 32125 10625 32137 10659
rect 32171 10625 32183 10659
rect 32125 10619 32183 10625
rect 31294 10588 31300 10600
rect 31036 10560 31300 10588
rect 31294 10548 31300 10560
rect 31352 10548 31358 10600
rect 23348 10492 28028 10520
rect 23348 10480 23354 10492
rect 30558 10480 30564 10532
rect 30616 10520 30622 10532
rect 30837 10523 30895 10529
rect 30837 10520 30849 10523
rect 30616 10492 30849 10520
rect 30616 10480 30622 10492
rect 30837 10489 30849 10492
rect 30883 10489 30895 10523
rect 30837 10483 30895 10489
rect 31202 10480 31208 10532
rect 31260 10520 31266 10532
rect 31404 10520 31432 10619
rect 32140 10588 32168 10619
rect 32214 10616 32220 10668
rect 32272 10656 32278 10668
rect 32404 10665 32462 10671
rect 32309 10659 32367 10665
rect 32309 10656 32321 10659
rect 32272 10628 32321 10656
rect 32272 10616 32278 10628
rect 32309 10625 32321 10628
rect 32355 10625 32367 10659
rect 32404 10631 32416 10665
rect 32450 10631 32462 10665
rect 32404 10625 32462 10631
rect 32309 10619 32367 10625
rect 32490 10616 32496 10668
rect 32548 10656 32554 10668
rect 32950 10656 32956 10668
rect 32548 10628 32956 10656
rect 32548 10616 32554 10628
rect 32950 10616 32956 10628
rect 33008 10616 33014 10668
rect 34517 10659 34575 10665
rect 34517 10625 34529 10659
rect 34563 10656 34575 10659
rect 34716 10656 34744 10684
rect 34790 10665 34796 10668
rect 34563 10628 34744 10656
rect 34563 10625 34575 10628
rect 34517 10619 34575 10625
rect 34784 10619 34796 10665
rect 34848 10656 34854 10668
rect 37274 10656 37280 10668
rect 34848 10628 34884 10656
rect 37235 10628 37280 10656
rect 34790 10616 34796 10619
rect 34848 10616 34854 10628
rect 37274 10616 37280 10628
rect 37332 10616 37338 10668
rect 37461 10659 37519 10665
rect 37461 10625 37473 10659
rect 37507 10625 37519 10659
rect 37461 10619 37519 10625
rect 32858 10588 32864 10600
rect 32140 10560 32864 10588
rect 32858 10548 32864 10560
rect 32916 10548 32922 10600
rect 36998 10548 37004 10600
rect 37056 10588 37062 10600
rect 37476 10588 37504 10619
rect 39298 10616 39304 10668
rect 39356 10656 39362 10668
rect 39868 10665 39896 10696
rect 39586 10659 39644 10665
rect 39586 10656 39598 10659
rect 39356 10628 39598 10656
rect 39356 10616 39362 10628
rect 39586 10625 39598 10628
rect 39632 10625 39644 10659
rect 39586 10619 39644 10625
rect 39853 10659 39911 10665
rect 39853 10625 39865 10659
rect 39899 10625 39911 10659
rect 39853 10619 39911 10625
rect 37056 10560 38516 10588
rect 37056 10548 37062 10560
rect 34422 10520 34428 10532
rect 31260 10492 31432 10520
rect 31726 10492 34428 10520
rect 31260 10480 31266 10492
rect 24670 10452 24676 10464
rect 22066 10424 24676 10452
rect 24670 10412 24676 10424
rect 24728 10412 24734 10464
rect 24946 10412 24952 10464
rect 25004 10452 25010 10464
rect 31726 10452 31754 10492
rect 34422 10480 34428 10492
rect 34480 10480 34486 10532
rect 38488 10529 38516 10560
rect 38473 10523 38531 10529
rect 38473 10489 38485 10523
rect 38519 10489 38531 10523
rect 38473 10483 38531 10489
rect 25004 10424 31754 10452
rect 32769 10455 32827 10461
rect 25004 10412 25010 10424
rect 32769 10421 32781 10455
rect 32815 10452 32827 10455
rect 33226 10452 33232 10464
rect 32815 10424 33232 10452
rect 32815 10421 32827 10424
rect 32769 10415 32827 10421
rect 33226 10412 33232 10424
rect 33284 10412 33290 10464
rect 35894 10452 35900 10464
rect 35855 10424 35900 10452
rect 35894 10412 35900 10424
rect 35952 10412 35958 10464
rect 58158 10452 58164 10464
rect 58119 10424 58164 10452
rect 58158 10412 58164 10424
rect 58216 10412 58222 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11054 10248 11060 10260
rect 10919 10220 11060 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 21910 10248 21916 10260
rect 19720 10220 21916 10248
rect 8941 10183 8999 10189
rect 8941 10149 8953 10183
rect 8987 10149 8999 10183
rect 8941 10143 8999 10149
rect 17221 10183 17279 10189
rect 17221 10149 17233 10183
rect 17267 10180 17279 10183
rect 19150 10180 19156 10192
rect 17267 10152 19156 10180
rect 17267 10149 17279 10152
rect 17221 10143 17279 10149
rect 6086 10112 6092 10124
rect 6047 10084 6092 10112
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 6270 10004 6276 10056
rect 6328 10044 6334 10056
rect 6365 10047 6423 10053
rect 6365 10044 6377 10047
rect 6328 10016 6377 10044
rect 6328 10004 6334 10016
rect 6365 10013 6377 10016
rect 6411 10013 6423 10047
rect 7190 10044 7196 10056
rect 7151 10016 7196 10044
rect 6365 10007 6423 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8956 10044 8984 10143
rect 19150 10140 19156 10152
rect 19208 10140 19214 10192
rect 9582 10112 9588 10124
rect 9543 10084 9588 10112
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 12618 10112 12624 10124
rect 12406 10084 12624 10112
rect 12406 10044 12434 10084
rect 12618 10072 12624 10084
rect 12676 10112 12682 10124
rect 13081 10115 13139 10121
rect 13081 10112 13093 10115
rect 12676 10084 13093 10112
rect 12676 10072 12682 10084
rect 13081 10081 13093 10084
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 16485 10115 16543 10121
rect 16485 10081 16497 10115
rect 16531 10112 16543 10115
rect 16574 10112 16580 10124
rect 16531 10084 16580 10112
rect 16531 10081 16543 10084
rect 16485 10075 16543 10081
rect 16574 10072 16580 10084
rect 16632 10112 16638 10124
rect 19720 10112 19748 10220
rect 21910 10208 21916 10220
rect 21968 10208 21974 10260
rect 22189 10251 22247 10257
rect 22189 10217 22201 10251
rect 22235 10248 22247 10251
rect 22554 10248 22560 10260
rect 22235 10220 22560 10248
rect 22235 10217 22247 10220
rect 22189 10211 22247 10217
rect 22554 10208 22560 10220
rect 22612 10208 22618 10260
rect 24670 10208 24676 10260
rect 24728 10248 24734 10260
rect 25041 10251 25099 10257
rect 25041 10248 25053 10251
rect 24728 10220 25053 10248
rect 24728 10208 24734 10220
rect 25041 10217 25053 10220
rect 25087 10217 25099 10251
rect 25041 10211 25099 10217
rect 31941 10251 31999 10257
rect 31941 10217 31953 10251
rect 31987 10248 31999 10251
rect 32214 10248 32220 10260
rect 31987 10220 32220 10248
rect 31987 10217 31999 10220
rect 31941 10211 31999 10217
rect 32214 10208 32220 10220
rect 32272 10208 32278 10260
rect 32490 10248 32496 10260
rect 32451 10220 32496 10248
rect 32490 10208 32496 10220
rect 32548 10208 32554 10260
rect 34701 10251 34759 10257
rect 34701 10217 34713 10251
rect 34747 10248 34759 10251
rect 34790 10248 34796 10260
rect 34747 10220 34796 10248
rect 34747 10217 34759 10220
rect 34701 10211 34759 10217
rect 34790 10208 34796 10220
rect 34848 10208 34854 10260
rect 34974 10248 34980 10260
rect 34900 10220 34980 10248
rect 29362 10180 29368 10192
rect 28460 10152 29368 10180
rect 16632 10084 19748 10112
rect 16632 10072 16638 10084
rect 22922 10072 22928 10124
rect 22980 10112 22986 10124
rect 24489 10115 24547 10121
rect 24489 10112 24501 10115
rect 22980 10084 24501 10112
rect 22980 10072 22986 10084
rect 13262 10044 13268 10056
rect 8067 10016 8984 10044
rect 9048 10016 12434 10044
rect 13223 10016 13268 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 4614 9936 4620 9988
rect 4672 9976 4678 9988
rect 7944 9976 7972 10007
rect 9048 9976 9076 10016
rect 13262 10004 13268 10016
rect 13320 10004 13326 10056
rect 20806 10044 20812 10056
rect 20767 10016 20812 10044
rect 20806 10004 20812 10016
rect 20864 10004 20870 10056
rect 21076 10047 21134 10053
rect 21076 10013 21088 10047
rect 21122 10044 21134 10047
rect 22278 10044 22284 10056
rect 21122 10016 22284 10044
rect 21122 10013 21134 10016
rect 21076 10007 21134 10013
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 23584 10053 23612 10084
rect 24489 10081 24501 10084
rect 24535 10112 24547 10115
rect 27706 10112 27712 10124
rect 24535 10084 27712 10112
rect 24535 10081 24547 10084
rect 24489 10075 24547 10081
rect 27706 10072 27712 10084
rect 27764 10112 27770 10124
rect 28460 10121 28488 10152
rect 29362 10140 29368 10152
rect 29420 10180 29426 10192
rect 32306 10180 32312 10192
rect 29420 10152 32312 10180
rect 29420 10140 29426 10152
rect 32306 10140 32312 10152
rect 32364 10140 32370 10192
rect 34514 10140 34520 10192
rect 34572 10180 34578 10192
rect 34900 10180 34928 10220
rect 34974 10208 34980 10220
rect 35032 10248 35038 10260
rect 35805 10251 35863 10257
rect 35805 10248 35817 10251
rect 35032 10220 35817 10248
rect 35032 10208 35038 10220
rect 35805 10217 35817 10220
rect 35851 10217 35863 10251
rect 35805 10211 35863 10217
rect 37734 10180 37740 10192
rect 34572 10152 34928 10180
rect 35084 10152 37740 10180
rect 34572 10140 34578 10152
rect 28169 10115 28227 10121
rect 28169 10112 28181 10115
rect 27764 10084 28181 10112
rect 27764 10072 27770 10084
rect 28169 10081 28181 10084
rect 28215 10081 28227 10115
rect 28169 10075 28227 10081
rect 28445 10115 28503 10121
rect 28445 10081 28457 10115
rect 28491 10081 28503 10115
rect 28445 10075 28503 10081
rect 28966 10084 29684 10112
rect 23477 10047 23535 10053
rect 23477 10044 23489 10047
rect 22664 10016 23489 10044
rect 12158 9976 12164 9988
rect 4672 9948 9076 9976
rect 12119 9948 12164 9976
rect 4672 9936 4678 9948
rect 12158 9936 12164 9948
rect 12216 9936 12222 9988
rect 16301 9979 16359 9985
rect 16301 9945 16313 9979
rect 16347 9976 16359 9979
rect 16574 9976 16580 9988
rect 16347 9948 16580 9976
rect 16347 9945 16359 9948
rect 16301 9939 16359 9945
rect 16574 9936 16580 9948
rect 16632 9976 16638 9988
rect 17037 9979 17095 9985
rect 17037 9976 17049 9979
rect 16632 9948 17049 9976
rect 16632 9936 16638 9948
rect 17037 9945 17049 9948
rect 17083 9945 17095 9979
rect 17037 9939 17095 9945
rect 19426 9936 19432 9988
rect 19484 9976 19490 9988
rect 22094 9976 22100 9988
rect 19484 9948 22100 9976
rect 19484 9936 19490 9948
rect 22094 9936 22100 9948
rect 22152 9936 22158 9988
rect 2406 9908 2412 9920
rect 2367 9880 2412 9908
rect 2406 9868 2412 9880
rect 2464 9868 2470 9920
rect 7282 9908 7288 9920
rect 7243 9880 7288 9908
rect 7282 9868 7288 9880
rect 7340 9868 7346 9920
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 9122 9908 9128 9920
rect 8251 9880 9128 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9401 9911 9459 9917
rect 9401 9877 9413 9911
rect 9447 9908 9459 9911
rect 9674 9908 9680 9920
rect 9447 9880 9680 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 13354 9868 13360 9920
rect 13412 9908 13418 9920
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13412 9880 13461 9908
rect 13412 9868 13418 9880
rect 13449 9877 13461 9880
rect 13495 9877 13507 9911
rect 13449 9871 13507 9877
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9908 18751 9911
rect 18874 9908 18880 9920
rect 18739 9880 18880 9908
rect 18739 9877 18751 9880
rect 18693 9871 18751 9877
rect 18874 9868 18880 9880
rect 18932 9908 18938 9920
rect 19242 9908 19248 9920
rect 18932 9880 19248 9908
rect 18932 9868 18938 9880
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 19334 9868 19340 9920
rect 19392 9908 19398 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19392 9880 19625 9908
rect 19392 9868 19398 9880
rect 19613 9877 19625 9880
rect 19659 9877 19671 9911
rect 19613 9871 19671 9877
rect 21082 9868 21088 9920
rect 21140 9908 21146 9920
rect 22664 9917 22692 10016
rect 23477 10013 23489 10016
rect 23523 10013 23535 10047
rect 23477 10007 23535 10013
rect 23569 10047 23627 10053
rect 23569 10013 23581 10047
rect 23615 10013 23627 10047
rect 23569 10007 23627 10013
rect 23658 10004 23664 10056
rect 23716 10044 23722 10056
rect 23845 10047 23903 10053
rect 23716 10016 23761 10044
rect 23716 10004 23722 10016
rect 23845 10013 23857 10047
rect 23891 10013 23903 10047
rect 23845 10007 23903 10013
rect 22738 9936 22744 9988
rect 22796 9976 22802 9988
rect 23382 9976 23388 9988
rect 22796 9948 23388 9976
rect 22796 9936 22802 9948
rect 23382 9936 23388 9948
rect 23440 9976 23446 9988
rect 23860 9976 23888 10007
rect 24026 10004 24032 10056
rect 24084 10044 24090 10056
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 24084 10016 24409 10044
rect 24084 10004 24090 10016
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10044 24639 10047
rect 24670 10044 24676 10056
rect 24627 10016 24676 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 26694 10004 26700 10056
rect 26752 10044 26758 10056
rect 28966 10044 28994 10084
rect 29546 10044 29552 10056
rect 26752 10016 28994 10044
rect 29507 10016 29552 10044
rect 26752 10004 26758 10016
rect 29546 10004 29552 10016
rect 29604 10004 29610 10056
rect 29656 10044 29684 10084
rect 29730 10072 29736 10124
rect 29788 10112 29794 10124
rect 29825 10115 29883 10121
rect 29825 10112 29837 10115
rect 29788 10084 29837 10112
rect 29788 10072 29794 10084
rect 29825 10081 29837 10084
rect 29871 10081 29883 10115
rect 29825 10075 29883 10081
rect 34057 10047 34115 10053
rect 34057 10044 34069 10047
rect 29656 10016 34069 10044
rect 34057 10013 34069 10016
rect 34103 10013 34115 10047
rect 34974 10044 34980 10056
rect 34935 10016 34980 10044
rect 34057 10007 34115 10013
rect 27338 9976 27344 9988
rect 23440 9948 23888 9976
rect 27299 9948 27344 9976
rect 23440 9936 23446 9948
rect 27338 9936 27344 9948
rect 27396 9936 27402 9988
rect 27525 9979 27583 9985
rect 27525 9945 27537 9979
rect 27571 9976 27583 9979
rect 31110 9976 31116 9988
rect 27571 9948 31116 9976
rect 27571 9945 27583 9948
rect 27525 9939 27583 9945
rect 31110 9936 31116 9948
rect 31168 9936 31174 9988
rect 31570 9976 31576 9988
rect 31531 9948 31576 9976
rect 31570 9936 31576 9948
rect 31628 9936 31634 9988
rect 31757 9979 31815 9985
rect 31757 9945 31769 9979
rect 31803 9976 31815 9979
rect 32122 9976 32128 9988
rect 31803 9948 32128 9976
rect 31803 9945 31815 9948
rect 31757 9939 31815 9945
rect 32122 9936 32128 9948
rect 32180 9936 32186 9988
rect 22649 9911 22707 9917
rect 22649 9908 22661 9911
rect 21140 9880 22661 9908
rect 21140 9868 21146 9880
rect 22649 9877 22661 9880
rect 22695 9877 22707 9911
rect 23198 9908 23204 9920
rect 23159 9880 23204 9908
rect 22649 9871 22707 9877
rect 23198 9868 23204 9880
rect 23256 9868 23262 9920
rect 27709 9911 27767 9917
rect 27709 9877 27721 9911
rect 27755 9908 27767 9911
rect 28534 9908 28540 9920
rect 27755 9880 28540 9908
rect 27755 9877 27767 9880
rect 27709 9871 27767 9877
rect 28534 9868 28540 9880
rect 28592 9868 28598 9920
rect 34072 9908 34100 10007
rect 34974 10004 34980 10016
rect 35032 10004 35038 10056
rect 35084 10053 35112 10152
rect 37734 10140 37740 10152
rect 37792 10140 37798 10192
rect 35434 10112 35440 10124
rect 35268 10084 35440 10112
rect 35069 10047 35127 10053
rect 35069 10013 35081 10047
rect 35115 10013 35127 10047
rect 35069 10007 35127 10013
rect 35182 10047 35240 10053
rect 35182 10013 35194 10047
rect 35228 10044 35240 10047
rect 35268 10044 35296 10084
rect 35434 10072 35440 10084
rect 35492 10072 35498 10124
rect 38010 10112 38016 10124
rect 36648 10084 38016 10112
rect 35228 10016 35296 10044
rect 35228 10013 35240 10016
rect 35182 10007 35240 10013
rect 35342 10004 35348 10056
rect 35400 10044 35406 10056
rect 36648 10053 36676 10084
rect 38010 10072 38016 10084
rect 38068 10072 38074 10124
rect 36633 10047 36691 10053
rect 35400 10016 35445 10044
rect 35400 10004 35406 10016
rect 36633 10013 36645 10047
rect 36679 10013 36691 10047
rect 36814 10044 36820 10056
rect 36775 10016 36820 10044
rect 36633 10007 36691 10013
rect 36814 10004 36820 10016
rect 36872 10004 36878 10056
rect 37274 10004 37280 10056
rect 37332 10044 37338 10056
rect 37332 10016 38240 10044
rect 37332 10004 37338 10016
rect 36832 9976 36860 10004
rect 38212 9985 38240 10016
rect 38013 9979 38071 9985
rect 38013 9976 38025 9979
rect 35912 9948 36860 9976
rect 37108 9948 38025 9976
rect 35250 9908 35256 9920
rect 34072 9880 35256 9908
rect 35250 9868 35256 9880
rect 35308 9868 35314 9920
rect 35342 9868 35348 9920
rect 35400 9908 35406 9920
rect 35912 9908 35940 9948
rect 35400 9880 35940 9908
rect 35400 9868 35406 9880
rect 36262 9868 36268 9920
rect 36320 9908 36326 9920
rect 36449 9911 36507 9917
rect 36449 9908 36461 9911
rect 36320 9880 36461 9908
rect 36320 9868 36326 9880
rect 36449 9877 36461 9880
rect 36495 9877 36507 9911
rect 36449 9871 36507 9877
rect 36538 9868 36544 9920
rect 36596 9908 36602 9920
rect 37108 9908 37136 9948
rect 38013 9945 38025 9948
rect 38059 9945 38071 9979
rect 38013 9939 38071 9945
rect 38197 9979 38255 9985
rect 38197 9945 38209 9979
rect 38243 9976 38255 9979
rect 38378 9976 38384 9988
rect 38243 9948 38384 9976
rect 38243 9945 38255 9948
rect 38197 9939 38255 9945
rect 37274 9908 37280 9920
rect 36596 9880 37136 9908
rect 37235 9880 37280 9908
rect 36596 9868 36602 9880
rect 37274 9868 37280 9880
rect 37332 9868 37338 9920
rect 37458 9868 37464 9920
rect 37516 9908 37522 9920
rect 37829 9911 37887 9917
rect 37829 9908 37841 9911
rect 37516 9880 37841 9908
rect 37516 9868 37522 9880
rect 37829 9877 37841 9880
rect 37875 9877 37887 9911
rect 38028 9908 38056 9939
rect 38378 9936 38384 9948
rect 38436 9936 38442 9988
rect 39942 9908 39948 9920
rect 38028 9880 39948 9908
rect 37829 9871 37887 9877
rect 39942 9868 39948 9880
rect 40000 9868 40006 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 9674 9704 9680 9716
rect 9635 9676 9680 9704
rect 9674 9664 9680 9676
rect 9732 9704 9738 9716
rect 11701 9707 11759 9713
rect 9732 9676 10456 9704
rect 9732 9664 9738 9676
rect 2406 9645 2412 9648
rect 2400 9636 2412 9645
rect 2367 9608 2412 9636
rect 2400 9599 2412 9608
rect 2406 9596 2412 9599
rect 2464 9596 2470 9648
rect 7834 9636 7840 9648
rect 5552 9608 7840 9636
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9568 4399 9571
rect 5258 9568 5264 9580
rect 4387 9540 5264 9568
rect 4387 9537 4399 9540
rect 4341 9531 4399 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 2130 9500 2136 9512
rect 2091 9472 2136 9500
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9469 4491 9503
rect 4433 9463 4491 9469
rect 3513 9435 3571 9441
rect 3513 9401 3525 9435
rect 3559 9432 3571 9435
rect 4448 9432 4476 9463
rect 4614 9460 4620 9512
rect 4672 9500 4678 9512
rect 5552 9500 5580 9608
rect 7834 9596 7840 9608
rect 7892 9596 7898 9648
rect 7926 9596 7932 9648
rect 7984 9636 7990 9648
rect 7984 9608 9352 9636
rect 7984 9596 7990 9608
rect 6362 9528 6368 9580
rect 6420 9568 6426 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6420 9540 6561 9568
rect 6420 9528 6426 9540
rect 6549 9537 6561 9540
rect 6595 9568 6607 9571
rect 7006 9568 7012 9580
rect 6595 9540 7012 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8297 9571 8355 9577
rect 8297 9568 8309 9571
rect 8260 9540 8309 9568
rect 8260 9528 8266 9540
rect 8297 9537 8309 9540
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 8564 9571 8622 9577
rect 8564 9537 8576 9571
rect 8610 9568 8622 9571
rect 8938 9568 8944 9580
rect 8610 9540 8944 9568
rect 8610 9537 8622 9540
rect 8564 9531 8622 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 4672 9472 5580 9500
rect 4672 9460 4678 9472
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6822 9500 6828 9512
rect 5684 9472 6828 9500
rect 5684 9460 5690 9472
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 5534 9432 5540 9444
rect 3559 9404 5540 9432
rect 3559 9401 3571 9404
rect 3513 9395 3571 9401
rect 5534 9392 5540 9404
rect 5592 9392 5598 9444
rect 9324 9432 9352 9608
rect 10042 9596 10048 9648
rect 10100 9636 10106 9648
rect 10137 9639 10195 9645
rect 10137 9636 10149 9639
rect 10100 9608 10149 9636
rect 10100 9596 10106 9608
rect 10137 9605 10149 9608
rect 10183 9605 10195 9639
rect 10137 9599 10195 9605
rect 10428 9577 10456 9676
rect 11701 9673 11713 9707
rect 11747 9704 11759 9707
rect 12158 9704 12164 9716
rect 11747 9676 12164 9704
rect 11747 9673 11759 9676
rect 11701 9667 11759 9673
rect 12158 9664 12164 9676
rect 12216 9704 12222 9716
rect 22370 9704 22376 9716
rect 12216 9676 22376 9704
rect 12216 9664 12222 9676
rect 22370 9664 22376 9676
rect 22428 9664 22434 9716
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 24489 9707 24547 9713
rect 24489 9704 24501 9707
rect 23716 9676 24501 9704
rect 23716 9664 23722 9676
rect 24489 9673 24501 9676
rect 24535 9673 24547 9707
rect 24489 9667 24547 9673
rect 28074 9664 28080 9716
rect 28132 9704 28138 9716
rect 34698 9704 34704 9716
rect 28132 9676 34468 9704
rect 28132 9664 28138 9676
rect 13446 9636 13452 9648
rect 12176 9608 13452 9636
rect 12176 9577 12204 9608
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 18138 9636 18144 9648
rect 14476 9608 18144 9636
rect 12434 9577 12440 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12428 9531 12440 9577
rect 12492 9568 12498 9580
rect 12492 9540 12528 9568
rect 12434 9528 12440 9531
rect 12492 9528 12498 9540
rect 10318 9500 10324 9512
rect 10279 9472 10324 9500
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10778 9500 10784 9512
rect 10739 9472 10784 9500
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 14476 9432 14504 9608
rect 18138 9596 18144 9608
rect 18196 9596 18202 9648
rect 19153 9639 19211 9645
rect 19153 9605 19165 9639
rect 19199 9636 19211 9639
rect 20162 9636 20168 9648
rect 19199 9608 20168 9636
rect 19199 9605 19211 9608
rect 19153 9599 19211 9605
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 14608 9540 15209 9568
rect 14608 9528 14614 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 15197 9531 15255 9537
rect 17972 9540 18337 9568
rect 17972 9512 18000 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9500 17371 9503
rect 17954 9500 17960 9512
rect 17359 9472 17960 9500
rect 17359 9469 17371 9472
rect 17313 9463 17371 9469
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 19168 9432 19196 9599
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 25590 9636 25596 9648
rect 22664 9608 25596 9636
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19797 9571 19855 9577
rect 19797 9568 19809 9571
rect 19392 9540 19809 9568
rect 19392 9528 19398 9540
rect 19797 9537 19809 9540
rect 19843 9537 19855 9571
rect 19978 9568 19984 9580
rect 19939 9540 19984 9568
rect 19797 9531 19855 9537
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 22664 9577 22692 9608
rect 25590 9596 25596 9608
rect 25648 9596 25654 9648
rect 31570 9636 31576 9648
rect 27908 9608 31576 9636
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 22916 9571 22974 9577
rect 22916 9537 22928 9571
rect 22962 9568 22974 9571
rect 23198 9568 23204 9580
rect 22962 9540 23204 9568
rect 22962 9537 22974 9540
rect 22916 9531 22974 9537
rect 23198 9528 23204 9540
rect 23256 9528 23262 9580
rect 24673 9571 24731 9577
rect 24673 9568 24685 9571
rect 24044 9540 24685 9568
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9500 19947 9503
rect 20438 9500 20444 9512
rect 19935 9472 20444 9500
rect 19935 9469 19947 9472
rect 19889 9463 19947 9469
rect 20438 9460 20444 9472
rect 20496 9460 20502 9512
rect 20717 9503 20775 9509
rect 20717 9469 20729 9503
rect 20763 9500 20775 9503
rect 20763 9472 22094 9500
rect 20763 9469 20775 9472
rect 20717 9463 20775 9469
rect 9324 9404 11560 9432
rect 3970 9364 3976 9376
rect 3931 9336 3976 9364
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 5258 9364 5264 9376
rect 5219 9336 5264 9364
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 11532 9364 11560 9404
rect 13096 9404 14504 9432
rect 18248 9404 19196 9432
rect 19337 9435 19395 9441
rect 13096 9364 13124 9404
rect 11532 9336 13124 9364
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 13541 9367 13599 9373
rect 13541 9364 13553 9367
rect 13228 9336 13553 9364
rect 13228 9324 13234 9336
rect 13541 9333 13553 9336
rect 13587 9333 13599 9367
rect 14550 9364 14556 9376
rect 14511 9336 14556 9364
rect 13541 9327 13599 9333
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15378 9364 15384 9376
rect 15335 9336 15384 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15378 9324 15384 9336
rect 15436 9364 15442 9376
rect 16850 9364 16856 9376
rect 15436 9336 16856 9364
rect 15436 9324 15442 9336
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 17865 9367 17923 9373
rect 17865 9333 17877 9367
rect 17911 9364 17923 9367
rect 18248 9364 18276 9404
rect 19337 9401 19349 9435
rect 19383 9432 19395 9435
rect 19426 9432 19432 9444
rect 19383 9404 19432 9432
rect 19383 9401 19395 9404
rect 19337 9395 19395 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 18506 9364 18512 9376
rect 17911 9336 18276 9364
rect 18467 9336 18512 9364
rect 17911 9333 17923 9336
rect 17865 9327 17923 9333
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 22066 9364 22094 9472
rect 24044 9376 24072 9540
rect 24673 9537 24685 9540
rect 24719 9537 24731 9571
rect 24673 9531 24731 9537
rect 24762 9528 24768 9580
rect 24820 9568 24826 9580
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24820 9540 24869 9568
rect 24820 9528 24826 9540
rect 24857 9537 24869 9540
rect 24903 9537 24915 9571
rect 25314 9568 25320 9580
rect 25275 9540 25320 9568
rect 24857 9531 24915 9537
rect 24872 9500 24900 9531
rect 25314 9528 25320 9540
rect 25372 9528 25378 9580
rect 25498 9568 25504 9580
rect 25459 9540 25504 9568
rect 25498 9528 25504 9540
rect 25556 9528 25562 9580
rect 27908 9577 27936 9608
rect 31570 9596 31576 9608
rect 31628 9596 31634 9648
rect 33226 9596 33232 9648
rect 33284 9645 33290 9648
rect 33284 9636 33296 9645
rect 33284 9608 33329 9636
rect 33284 9599 33296 9608
rect 33284 9596 33290 9599
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9568 27215 9571
rect 27617 9571 27675 9577
rect 27617 9568 27629 9571
rect 27203 9540 27629 9568
rect 27203 9537 27215 9540
rect 27157 9531 27215 9537
rect 27617 9537 27629 9540
rect 27663 9537 27675 9571
rect 27617 9531 27675 9537
rect 27893 9571 27951 9577
rect 27893 9537 27905 9571
rect 27939 9537 27951 9571
rect 27893 9531 27951 9537
rect 29825 9571 29883 9577
rect 29825 9537 29837 9571
rect 29871 9568 29883 9571
rect 30374 9568 30380 9580
rect 29871 9540 30380 9568
rect 29871 9537 29883 9540
rect 29825 9531 29883 9537
rect 27172 9500 27200 9531
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 31726 9540 34376 9568
rect 24872 9472 27200 9500
rect 27982 9460 27988 9512
rect 28040 9500 28046 9512
rect 28902 9500 28908 9512
rect 28040 9472 28908 9500
rect 28040 9460 28046 9472
rect 28902 9460 28908 9472
rect 28960 9500 28966 9512
rect 29549 9503 29607 9509
rect 29549 9500 29561 9503
rect 28960 9472 29561 9500
rect 28960 9460 28966 9472
rect 29549 9469 29561 9472
rect 29595 9469 29607 9503
rect 29549 9463 29607 9469
rect 25314 9392 25320 9444
rect 25372 9432 25378 9444
rect 25372 9404 26188 9432
rect 25372 9392 25378 9404
rect 26160 9376 26188 9404
rect 27798 9392 27804 9444
rect 27856 9432 27862 9444
rect 31726 9432 31754 9540
rect 33505 9503 33563 9509
rect 33505 9469 33517 9503
rect 33551 9469 33563 9503
rect 33505 9463 33563 9469
rect 27856 9404 31754 9432
rect 27856 9392 27862 9404
rect 23290 9364 23296 9376
rect 22066 9336 23296 9364
rect 23290 9324 23296 9336
rect 23348 9324 23354 9376
rect 24026 9364 24032 9376
rect 23987 9336 24032 9364
rect 24026 9324 24032 9336
rect 24084 9324 24090 9376
rect 25406 9324 25412 9376
rect 25464 9364 25470 9376
rect 25685 9367 25743 9373
rect 25685 9364 25697 9367
rect 25464 9336 25697 9364
rect 25464 9324 25470 9336
rect 25685 9333 25697 9336
rect 25731 9333 25743 9367
rect 25685 9327 25743 9333
rect 26142 9324 26148 9376
rect 26200 9364 26206 9376
rect 26973 9367 27031 9373
rect 26973 9364 26985 9367
rect 26200 9336 26985 9364
rect 26200 9324 26206 9336
rect 26973 9333 26985 9336
rect 27019 9364 27031 9367
rect 27338 9364 27344 9376
rect 27019 9336 27344 9364
rect 27019 9333 27031 9336
rect 26973 9327 27031 9333
rect 27338 9324 27344 9336
rect 27396 9324 27402 9376
rect 32122 9364 32128 9376
rect 32083 9336 32128 9364
rect 32122 9324 32128 9336
rect 32180 9324 32186 9376
rect 32766 9324 32772 9376
rect 32824 9364 32830 9376
rect 33520 9364 33548 9463
rect 34348 9441 34376 9540
rect 34333 9435 34391 9441
rect 34333 9401 34345 9435
rect 34379 9401 34391 9435
rect 34440 9432 34468 9676
rect 34532 9676 34704 9704
rect 34532 9577 34560 9676
rect 34698 9664 34704 9676
rect 34756 9664 34762 9716
rect 36630 9704 36636 9716
rect 36372 9676 36636 9704
rect 34609 9639 34667 9645
rect 34609 9605 34621 9639
rect 34655 9636 34667 9639
rect 35894 9636 35900 9648
rect 34655 9608 35900 9636
rect 34655 9605 34667 9608
rect 34609 9599 34667 9605
rect 35894 9596 35900 9608
rect 35952 9596 35958 9648
rect 35986 9596 35992 9648
rect 36044 9636 36050 9648
rect 36372 9636 36400 9676
rect 36630 9664 36636 9676
rect 36688 9664 36694 9716
rect 37274 9664 37280 9716
rect 37332 9704 37338 9716
rect 39942 9704 39948 9716
rect 37332 9676 38025 9704
rect 39903 9676 39948 9704
rect 37332 9664 37338 9676
rect 36044 9608 36400 9636
rect 36044 9596 36050 9608
rect 34517 9571 34575 9577
rect 34517 9537 34529 9571
rect 34563 9537 34575 9571
rect 34698 9568 34704 9580
rect 34659 9540 34704 9568
rect 34517 9531 34575 9537
rect 34532 9500 34560 9531
rect 34698 9528 34704 9540
rect 34756 9528 34762 9580
rect 34790 9528 34796 9580
rect 34848 9568 34854 9580
rect 34885 9571 34943 9577
rect 34885 9568 34897 9571
rect 34848 9540 34897 9568
rect 34848 9528 34854 9540
rect 34885 9537 34897 9540
rect 34931 9537 34943 9571
rect 34885 9531 34943 9537
rect 36081 9571 36139 9577
rect 36081 9537 36093 9571
rect 36127 9537 36139 9571
rect 36262 9568 36268 9580
rect 36223 9540 36268 9568
rect 36081 9531 36139 9537
rect 35434 9500 35440 9512
rect 34532 9472 35440 9500
rect 35434 9460 35440 9472
rect 35492 9460 35498 9512
rect 35618 9460 35624 9512
rect 35676 9500 35682 9512
rect 36096 9500 36124 9531
rect 36262 9528 36268 9540
rect 36320 9528 36326 9580
rect 36372 9577 36400 9608
rect 36357 9571 36415 9577
rect 36357 9537 36369 9571
rect 36403 9537 36415 9571
rect 36357 9531 36415 9537
rect 36449 9571 36507 9577
rect 36449 9537 36461 9571
rect 36495 9537 36507 9571
rect 36449 9531 36507 9537
rect 36464 9500 36492 9531
rect 37182 9528 37188 9580
rect 37240 9568 37246 9580
rect 37624 9577 37682 9583
rect 37449 9571 37507 9577
rect 37624 9574 37636 9577
rect 37449 9568 37461 9571
rect 37240 9540 37461 9568
rect 37240 9528 37246 9540
rect 37449 9537 37461 9540
rect 37495 9537 37507 9571
rect 37449 9531 37507 9537
rect 37568 9546 37636 9574
rect 37274 9500 37280 9512
rect 35676 9472 36124 9500
rect 36372 9472 37280 9500
rect 35676 9460 35682 9472
rect 35529 9435 35587 9441
rect 35529 9432 35541 9435
rect 34440 9404 35541 9432
rect 34333 9395 34391 9401
rect 35529 9401 35541 9404
rect 35575 9432 35587 9435
rect 36372 9432 36400 9472
rect 37274 9460 37280 9472
rect 37332 9460 37338 9512
rect 35575 9404 36400 9432
rect 35575 9401 35587 9404
rect 35529 9395 35587 9401
rect 37458 9392 37464 9444
rect 37516 9432 37522 9444
rect 37568 9432 37596 9546
rect 37624 9543 37636 9546
rect 37670 9543 37682 9577
rect 37624 9537 37682 9543
rect 37721 9531 37727 9583
rect 37779 9574 37785 9583
rect 37779 9546 37821 9574
rect 37875 9571 37933 9577
rect 37779 9531 37785 9546
rect 37875 9537 37887 9571
rect 37921 9568 37933 9571
rect 37997 9568 38025 9676
rect 39942 9664 39948 9676
rect 40000 9664 40006 9716
rect 38105 9639 38163 9645
rect 38105 9605 38117 9639
rect 38151 9636 38163 9639
rect 38810 9639 38868 9645
rect 38810 9636 38822 9639
rect 38151 9608 38822 9636
rect 38151 9605 38163 9608
rect 38105 9599 38163 9605
rect 38810 9605 38822 9608
rect 38856 9605 38868 9639
rect 38810 9599 38868 9605
rect 38562 9568 38568 9580
rect 37921 9540 38025 9568
rect 38523 9540 38568 9568
rect 37921 9537 37933 9540
rect 37875 9531 37933 9537
rect 38562 9528 38568 9540
rect 38620 9528 38626 9580
rect 37516 9404 37596 9432
rect 37516 9392 37522 9404
rect 32824 9336 33548 9364
rect 32824 9324 32830 9336
rect 36630 9324 36636 9376
rect 36688 9364 36694 9376
rect 36725 9367 36783 9373
rect 36725 9364 36737 9367
rect 36688 9336 36737 9364
rect 36688 9324 36694 9336
rect 36725 9333 36737 9336
rect 36771 9333 36783 9367
rect 36725 9327 36783 9333
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 2685 9163 2743 9169
rect 2685 9160 2697 9163
rect 2648 9132 2697 9160
rect 2648 9120 2654 9132
rect 2685 9129 2697 9132
rect 2731 9129 2743 9163
rect 8938 9160 8944 9172
rect 8899 9132 8944 9160
rect 2685 9123 2743 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 12805 9163 12863 9169
rect 10060 9132 12664 9160
rect 3878 9052 3884 9104
rect 3936 9092 3942 9104
rect 4157 9095 4215 9101
rect 4157 9092 4169 9095
rect 3936 9064 4169 9092
rect 3936 9052 3942 9064
rect 4157 9061 4169 9064
rect 4203 9061 4215 9095
rect 4157 9055 4215 9061
rect 3970 9024 3976 9036
rect 2884 8996 3976 9024
rect 2884 8965 2912 8996
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 4706 9024 4712 9036
rect 4264 8996 4712 9024
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 4264 8956 4292 8996
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 6822 8984 6828 9036
rect 6880 9024 6886 9036
rect 10060 9033 10088 9132
rect 12526 9092 12532 9104
rect 10336 9064 10916 9092
rect 10336 9036 10364 9064
rect 10045 9027 10103 9033
rect 6880 8996 9260 9024
rect 6880 8984 6886 8996
rect 3099 8928 4292 8956
rect 4341 8959 4399 8965
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 4614 8956 4620 8968
rect 4387 8928 4620 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6365 8959 6423 8965
rect 6365 8956 6377 8959
rect 6328 8928 6377 8956
rect 6328 8916 6334 8928
rect 6365 8925 6377 8928
rect 6411 8925 6423 8959
rect 6365 8919 6423 8925
rect 6641 8959 6699 8965
rect 6641 8925 6653 8959
rect 6687 8956 6699 8959
rect 7190 8956 7196 8968
rect 6687 8928 7196 8956
rect 6687 8925 6699 8928
rect 6641 8919 6699 8925
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 6656 8888 6684 8919
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 7432 8928 7665 8956
rect 7432 8916 7438 8928
rect 7653 8925 7665 8928
rect 7699 8925 7711 8959
rect 9122 8956 9128 8968
rect 9083 8928 9128 8956
rect 7653 8919 7711 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9232 8956 9260 8996
rect 10045 8993 10057 9027
rect 10091 8993 10103 9027
rect 10318 9024 10324 9036
rect 10045 8987 10103 8993
rect 10152 8996 10324 9024
rect 10152 8965 10180 8996
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10778 9024 10784 9036
rect 10739 8996 10784 9024
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 9232 8928 10149 8956
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10796 8956 10824 8984
rect 10137 8919 10195 8925
rect 10244 8928 10824 8956
rect 10888 8956 10916 9064
rect 12268 9064 12532 9092
rect 12268 9033 12296 9064
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 9024 11207 9027
rect 12253 9027 12311 9033
rect 11195 8996 11836 9024
rect 11195 8993 11207 8996
rect 11149 8987 11207 8993
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 10888 8928 11253 8956
rect 5776 8860 6684 8888
rect 5776 8848 5782 8860
rect 6730 8848 6736 8900
rect 6788 8888 6794 8900
rect 9677 8891 9735 8897
rect 9677 8888 9689 8891
rect 6788 8860 9689 8888
rect 6788 8848 6794 8860
rect 9677 8857 9689 8860
rect 9723 8888 9735 8891
rect 10244 8888 10272 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11808 8956 11836 8996
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 12636 9024 12664 9132
rect 12805 9129 12817 9163
rect 12851 9160 12863 9163
rect 13262 9160 13268 9172
rect 12851 9132 13268 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 15562 9120 15568 9172
rect 15620 9160 15626 9172
rect 18598 9160 18604 9172
rect 15620 9132 18460 9160
rect 18559 9132 18604 9160
rect 15620 9120 15626 9132
rect 18432 9092 18460 9132
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 23198 9160 23204 9172
rect 18708 9132 23204 9160
rect 18708 9092 18736 9132
rect 23198 9120 23204 9132
rect 23256 9120 23262 9172
rect 23477 9163 23535 9169
rect 23477 9129 23489 9163
rect 23523 9160 23535 9163
rect 24118 9160 24124 9172
rect 23523 9132 24124 9160
rect 23523 9129 23535 9132
rect 23477 9123 23535 9129
rect 24118 9120 24124 9132
rect 24176 9120 24182 9172
rect 25314 9120 25320 9172
rect 25372 9160 25378 9172
rect 28258 9160 28264 9172
rect 25372 9132 28264 9160
rect 25372 9120 25378 9132
rect 28258 9120 28264 9132
rect 28316 9160 28322 9172
rect 28626 9160 28632 9172
rect 28316 9132 28632 9160
rect 28316 9120 28322 9132
rect 28626 9120 28632 9132
rect 28684 9160 28690 9172
rect 28905 9163 28963 9169
rect 28905 9160 28917 9163
rect 28684 9132 28917 9160
rect 28684 9120 28690 9132
rect 28905 9129 28917 9132
rect 28951 9129 28963 9163
rect 28905 9123 28963 9129
rect 31110 9120 31116 9172
rect 31168 9160 31174 9172
rect 31205 9163 31263 9169
rect 31205 9160 31217 9163
rect 31168 9132 31217 9160
rect 31168 9120 31174 9132
rect 31205 9129 31217 9132
rect 31251 9129 31263 9163
rect 31205 9123 31263 9129
rect 37737 9163 37795 9169
rect 37737 9129 37749 9163
rect 37783 9160 37795 9163
rect 38010 9160 38016 9172
rect 37783 9132 38016 9160
rect 37783 9129 37795 9132
rect 37737 9123 37795 9129
rect 38010 9120 38016 9132
rect 38068 9120 38074 9172
rect 23934 9092 23940 9104
rect 18432 9064 18736 9092
rect 22066 9064 23940 9092
rect 12802 9024 12808 9036
rect 12391 8996 12808 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12802 8984 12808 8996
rect 12860 8984 12866 9036
rect 17218 9024 17224 9036
rect 17179 8996 17224 9024
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 19889 9027 19947 9033
rect 19889 9024 19901 9027
rect 18248 8996 19901 9024
rect 13170 8956 13176 8968
rect 11808 8928 13176 8956
rect 11241 8919 11299 8925
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 13354 8956 13360 8968
rect 13315 8928 13360 8956
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 14918 8956 14924 8968
rect 13504 8928 14924 8956
rect 13504 8916 13510 8928
rect 14918 8916 14924 8928
rect 14976 8956 14982 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 14976 8928 15393 8956
rect 14976 8916 14982 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 18248 8956 18276 8996
rect 19889 8993 19901 8996
rect 19935 9024 19947 9027
rect 19978 9024 19984 9036
rect 19935 8996 19984 9024
rect 19935 8993 19947 8996
rect 19889 8987 19947 8993
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 20438 8984 20444 9036
rect 20496 9024 20502 9036
rect 20809 9027 20867 9033
rect 20809 9024 20821 9027
rect 20496 8996 20821 9024
rect 20496 8984 20502 8996
rect 20809 8993 20821 8996
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 21085 9027 21143 9033
rect 21085 8993 21097 9027
rect 21131 9024 21143 9027
rect 22066 9024 22094 9064
rect 23934 9052 23940 9064
rect 23992 9052 23998 9104
rect 25038 9052 25044 9104
rect 25096 9092 25102 9104
rect 25498 9092 25504 9104
rect 25096 9064 25504 9092
rect 25096 9052 25102 9064
rect 25498 9052 25504 9064
rect 25556 9052 25562 9104
rect 24026 9024 24032 9036
rect 21131 8996 22094 9024
rect 23216 8996 24032 9024
rect 21131 8993 21143 8996
rect 21085 8987 21143 8993
rect 19242 8956 19248 8968
rect 15381 8919 15439 8925
rect 16592 8928 18276 8956
rect 19203 8928 19248 8956
rect 9723 8860 10272 8888
rect 10321 8891 10379 8897
rect 9723 8857 9735 8860
rect 9677 8851 9735 8857
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 11974 8888 11980 8900
rect 10367 8860 11980 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 11974 8848 11980 8860
rect 12032 8848 12038 8900
rect 12066 8848 12072 8900
rect 12124 8888 12130 8900
rect 12124 8860 15424 8888
rect 12124 8848 12130 8860
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 5040 8792 5181 8820
rect 5040 8780 5046 8792
rect 5169 8789 5181 8792
rect 5215 8789 5227 8823
rect 5169 8783 5227 8789
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 6972 8792 7849 8820
rect 6972 8780 6978 8792
rect 7837 8789 7849 8792
rect 7883 8820 7895 8823
rect 11146 8820 11152 8832
rect 7883 8792 11152 8820
rect 7883 8789 7895 8792
rect 7837 8783 7895 8789
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 11296 8792 11437 8820
rect 11296 8780 11302 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 12437 8823 12495 8829
rect 12437 8789 12449 8823
rect 12483 8820 12495 8823
rect 12526 8820 12532 8832
rect 12483 8792 12532 8820
rect 12483 8789 12495 8792
rect 12437 8783 12495 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 13538 8820 13544 8832
rect 13499 8792 13544 8820
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 15396 8820 15424 8860
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 15626 8891 15684 8897
rect 15626 8888 15638 8891
rect 15528 8860 15638 8888
rect 15528 8848 15534 8860
rect 15626 8857 15638 8860
rect 15672 8857 15684 8891
rect 15626 8851 15684 8857
rect 16592 8820 16620 8928
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 19426 8956 19432 8968
rect 19387 8928 19432 8956
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 21266 8916 21272 8968
rect 21324 8956 21330 8968
rect 23216 8965 23244 8996
rect 24026 8984 24032 8996
rect 24084 8984 24090 9036
rect 25590 9024 25596 9036
rect 25551 8996 25596 9024
rect 25590 8984 25596 8996
rect 25648 8984 25654 9036
rect 27617 9027 27675 9033
rect 27617 8993 27629 9027
rect 27663 9024 27675 9027
rect 27706 9024 27712 9036
rect 27663 8996 27712 9024
rect 27663 8993 27675 8996
rect 27617 8987 27675 8993
rect 27706 8984 27712 8996
rect 27764 8984 27770 9036
rect 36354 9024 36360 9036
rect 36315 8996 36360 9024
rect 36354 8984 36360 8996
rect 36412 8984 36418 9036
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 21324 8928 22937 8956
rect 21324 8916 21330 8928
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23201 8959 23259 8965
rect 23201 8925 23213 8959
rect 23247 8925 23259 8959
rect 23201 8919 23259 8925
rect 23290 8916 23296 8968
rect 23348 8956 23354 8968
rect 27798 8956 27804 8968
rect 23348 8928 23393 8956
rect 25792 8928 27804 8956
rect 23348 8916 23354 8928
rect 17488 8891 17546 8897
rect 17488 8857 17500 8891
rect 17534 8888 17546 8891
rect 18046 8888 18052 8900
rect 17534 8860 18052 8888
rect 17534 8857 17546 8860
rect 17488 8851 17546 8857
rect 18046 8848 18052 8860
rect 18104 8848 18110 8900
rect 18506 8848 18512 8900
rect 18564 8888 18570 8900
rect 18564 8860 20024 8888
rect 18564 8848 18570 8860
rect 16758 8820 16764 8832
rect 15396 8792 16620 8820
rect 16719 8792 16764 8820
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 16850 8780 16856 8832
rect 16908 8820 16914 8832
rect 19150 8820 19156 8832
rect 16908 8792 19156 8820
rect 16908 8780 16914 8792
rect 19150 8780 19156 8792
rect 19208 8780 19214 8832
rect 19334 8820 19340 8832
rect 19295 8792 19340 8820
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 19996 8820 20024 8860
rect 21174 8848 21180 8900
rect 21232 8888 21238 8900
rect 22002 8888 22008 8900
rect 21232 8860 22008 8888
rect 21232 8848 21238 8860
rect 22002 8848 22008 8860
rect 22060 8888 22066 8900
rect 23109 8891 23167 8897
rect 23109 8888 23121 8891
rect 22060 8860 23121 8888
rect 22060 8848 22066 8860
rect 23109 8857 23121 8860
rect 23155 8888 23167 8891
rect 25792 8888 25820 8928
rect 27798 8916 27804 8928
rect 27856 8916 27862 8968
rect 27893 8959 27951 8965
rect 27893 8925 27905 8959
rect 27939 8956 27951 8959
rect 27982 8956 27988 8968
rect 27939 8928 27988 8956
rect 27939 8925 27951 8928
rect 27893 8919 27951 8925
rect 27982 8916 27988 8928
rect 28040 8916 28046 8968
rect 29822 8956 29828 8968
rect 29783 8928 29828 8956
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 36630 8965 36636 8968
rect 36624 8956 36636 8965
rect 36591 8928 36636 8956
rect 36624 8919 36636 8928
rect 36630 8916 36636 8919
rect 36688 8916 36694 8968
rect 58158 8956 58164 8968
rect 58119 8928 58164 8956
rect 58158 8916 58164 8928
rect 58216 8916 58222 8968
rect 25866 8897 25872 8900
rect 23155 8860 25820 8888
rect 23155 8857 23167 8860
rect 23109 8851 23167 8857
rect 25860 8851 25872 8897
rect 25924 8888 25930 8900
rect 25924 8860 25960 8888
rect 25866 8848 25872 8851
rect 25924 8848 25930 8860
rect 28994 8848 29000 8900
rect 29052 8888 29058 8900
rect 30070 8891 30128 8897
rect 30070 8888 30082 8891
rect 29052 8860 30082 8888
rect 29052 8848 29058 8860
rect 30070 8857 30082 8860
rect 30116 8857 30128 8891
rect 30070 8851 30128 8857
rect 25314 8820 25320 8832
rect 19996 8792 25320 8820
rect 25314 8780 25320 8792
rect 25372 8780 25378 8832
rect 25498 8780 25504 8832
rect 25556 8820 25562 8832
rect 26973 8823 27031 8829
rect 26973 8820 26985 8823
rect 25556 8792 26985 8820
rect 25556 8780 25562 8792
rect 26973 8789 26985 8792
rect 27019 8789 27031 8823
rect 26973 8783 27031 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 6178 8616 6184 8628
rect 4632 8588 6184 8616
rect 3786 8508 3792 8560
rect 3844 8548 3850 8560
rect 4632 8557 4660 8588
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 11701 8619 11759 8625
rect 11701 8616 11713 8619
rect 7892 8588 11713 8616
rect 7892 8576 7898 8588
rect 11701 8585 11713 8588
rect 11747 8585 11759 8619
rect 11701 8579 11759 8585
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 12860 8588 13553 8616
rect 12860 8576 12866 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 15010 8616 15016 8628
rect 13541 8579 13599 8585
rect 13740 8588 15016 8616
rect 4617 8551 4675 8557
rect 4617 8548 4629 8551
rect 3844 8520 4629 8548
rect 3844 8508 3850 8520
rect 4617 8517 4629 8520
rect 4663 8517 4675 8551
rect 4617 8511 4675 8517
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 5215 8520 6684 8548
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 5534 8480 5540 8492
rect 3191 8452 3372 8480
rect 5495 8452 5540 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3234 8412 3240 8424
rect 3195 8384 3240 8412
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 1762 8304 1768 8356
rect 1820 8344 1826 8356
rect 1949 8347 2007 8353
rect 1949 8344 1961 8347
rect 1820 8316 1961 8344
rect 1820 8304 1826 8316
rect 1949 8313 1961 8316
rect 1995 8313 2007 8347
rect 3344 8344 3372 8452
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 6656 8489 6684 8520
rect 7190 8508 7196 8560
rect 7248 8548 7254 8560
rect 7466 8548 7472 8560
rect 7248 8520 7472 8548
rect 7248 8508 7254 8520
rect 7466 8508 7472 8520
rect 7524 8548 7530 8560
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 7524 8520 8217 8548
rect 7524 8508 7530 8520
rect 8205 8517 8217 8520
rect 8251 8517 8263 8551
rect 13740 8548 13768 8588
rect 15010 8576 15016 8588
rect 15068 8616 15074 8628
rect 15562 8616 15568 8628
rect 15068 8588 15424 8616
rect 15523 8588 15568 8616
rect 15068 8576 15074 8588
rect 8205 8511 8263 8517
rect 8312 8520 13768 8548
rect 6641 8483 6699 8489
rect 5684 8452 5729 8480
rect 5684 8440 5690 8452
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 6730 8480 6736 8492
rect 6687 8452 6736 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 8312 8480 8340 8520
rect 7484 8452 8340 8480
rect 10965 8483 11023 8489
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8412 3479 8415
rect 4614 8412 4620 8424
rect 3467 8384 4620 8412
rect 3467 8381 3479 8384
rect 3421 8375 3479 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 5408 8384 6224 8412
rect 5408 8372 5414 8384
rect 3970 8344 3976 8356
rect 3344 8316 3976 8344
rect 1949 8307 2007 8313
rect 3970 8304 3976 8316
rect 4028 8304 4034 8356
rect 6196 8344 6224 8384
rect 6270 8372 6276 8424
rect 6328 8412 6334 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6328 8384 6377 8412
rect 6328 8372 6334 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 7484 8344 7512 8452
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11790 8480 11796 8492
rect 11011 8452 11796 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11790 8440 11796 8452
rect 11848 8480 11854 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11848 8452 11897 8480
rect 11848 8440 11854 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 12406 8452 13492 8480
rect 7558 8372 7564 8424
rect 7616 8412 7622 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 7616 8384 11529 8412
rect 7616 8372 7622 8384
rect 11517 8381 11529 8384
rect 11563 8412 11575 8415
rect 12406 8412 12434 8452
rect 12526 8412 12532 8424
rect 11563 8384 12434 8412
rect 12487 8384 12532 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 13464 8412 13492 8452
rect 13538 8440 13544 8492
rect 13596 8480 13602 8492
rect 15396 8489 15424 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 18046 8616 18052 8628
rect 18007 8588 18052 8616
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 18690 8616 18696 8628
rect 18196 8588 18696 8616
rect 18196 8576 18202 8588
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 23017 8619 23075 8625
rect 23017 8585 23029 8619
rect 23063 8616 23075 8619
rect 23106 8616 23112 8628
rect 23063 8588 23112 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 23106 8576 23112 8588
rect 23164 8576 23170 8628
rect 24670 8576 24676 8628
rect 24728 8616 24734 8628
rect 25866 8616 25872 8628
rect 24728 8588 25636 8616
rect 25827 8588 25872 8616
rect 24728 8576 24734 8588
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 22741 8551 22799 8557
rect 16816 8520 22094 8548
rect 16816 8508 16822 8520
rect 14654 8483 14712 8489
rect 14654 8480 14666 8483
rect 13596 8452 14666 8480
rect 13596 8440 13602 8452
rect 14654 8449 14666 8452
rect 14700 8449 14712 8483
rect 14654 8443 14712 8449
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8449 17187 8483
rect 18322 8480 18328 8492
rect 18283 8452 18328 8480
rect 17129 8443 17187 8449
rect 13906 8412 13912 8424
rect 13464 8384 13912 8412
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 14918 8412 14924 8424
rect 14879 8384 14924 8412
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 15102 8372 15108 8424
rect 15160 8412 15166 8424
rect 16574 8412 16580 8424
rect 15160 8384 16580 8412
rect 15160 8372 15166 8384
rect 16574 8372 16580 8384
rect 16632 8412 16638 8424
rect 17144 8412 17172 8443
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 16632 8384 17172 8412
rect 18432 8412 18460 8443
rect 18506 8440 18512 8492
rect 18564 8480 18570 8492
rect 18564 8452 18609 8480
rect 18564 8440 18570 8452
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 19705 8483 19763 8489
rect 18748 8452 18793 8480
rect 18748 8440 18754 8452
rect 19705 8449 19717 8483
rect 19751 8480 19763 8483
rect 21174 8480 21180 8492
rect 19751 8452 21180 8480
rect 19751 8449 19763 8452
rect 19705 8443 19763 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 22066 8480 22094 8520
rect 22741 8517 22753 8551
rect 22787 8548 22799 8551
rect 25038 8548 25044 8560
rect 22787 8520 25044 8548
rect 22787 8517 22799 8520
rect 22741 8511 22799 8517
rect 25038 8508 25044 8520
rect 25096 8508 25102 8560
rect 25608 8548 25636 8588
rect 25866 8576 25872 8588
rect 25924 8576 25930 8628
rect 27890 8616 27896 8628
rect 25976 8588 27896 8616
rect 25682 8548 25688 8560
rect 25595 8520 25688 8548
rect 22465 8483 22523 8489
rect 22465 8480 22477 8483
rect 22066 8452 22477 8480
rect 22465 8449 22477 8452
rect 22511 8449 22523 8483
rect 22465 8443 22523 8449
rect 22554 8440 22560 8492
rect 22612 8480 22618 8492
rect 22649 8483 22707 8489
rect 22649 8480 22661 8483
rect 22612 8452 22661 8480
rect 22612 8440 22618 8452
rect 22649 8449 22661 8452
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8480 22891 8483
rect 23474 8480 23480 8492
rect 22879 8452 23480 8480
rect 22879 8449 22891 8452
rect 22833 8443 22891 8449
rect 23474 8440 23480 8452
rect 23532 8480 23538 8492
rect 23934 8480 23940 8492
rect 23532 8452 23940 8480
rect 23532 8440 23538 8452
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 25222 8480 25228 8492
rect 25183 8452 25228 8480
rect 25222 8440 25228 8452
rect 25280 8440 25286 8492
rect 25406 8480 25412 8492
rect 25367 8452 25412 8480
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 25608 8489 25636 8520
rect 25682 8508 25688 8520
rect 25740 8548 25746 8560
rect 25976 8548 26004 8588
rect 27890 8576 27896 8588
rect 27948 8576 27954 8628
rect 28626 8576 28632 8628
rect 28684 8616 28690 8628
rect 28994 8616 29000 8628
rect 28684 8588 28764 8616
rect 28955 8588 29000 8616
rect 28684 8576 28690 8588
rect 25740 8520 26004 8548
rect 25740 8508 25746 8520
rect 27154 8508 27160 8560
rect 27212 8548 27218 8560
rect 27212 8520 27936 8548
rect 27212 8508 27218 8520
rect 25501 8483 25559 8489
rect 25501 8449 25513 8483
rect 25547 8449 25559 8483
rect 25501 8443 25559 8449
rect 25593 8483 25651 8489
rect 25593 8449 25605 8483
rect 25639 8449 25651 8483
rect 25593 8443 25651 8449
rect 19334 8412 19340 8424
rect 18432 8384 19340 8412
rect 16632 8372 16638 8384
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 19518 8412 19524 8424
rect 19475 8384 19524 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 19518 8372 19524 8384
rect 19576 8372 19582 8424
rect 20714 8412 20720 8424
rect 20675 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 23198 8372 23204 8424
rect 23256 8412 23262 8424
rect 24762 8412 24768 8424
rect 23256 8384 24768 8412
rect 23256 8372 23262 8384
rect 24762 8372 24768 8384
rect 24820 8412 24826 8424
rect 25516 8412 25544 8443
rect 27430 8440 27436 8492
rect 27488 8480 27494 8492
rect 27525 8483 27583 8489
rect 27525 8480 27537 8483
rect 27488 8452 27537 8480
rect 27488 8440 27494 8452
rect 27525 8449 27537 8452
rect 27571 8449 27583 8483
rect 27525 8443 27583 8449
rect 27617 8483 27675 8489
rect 27617 8449 27629 8483
rect 27663 8449 27675 8483
rect 27617 8443 27675 8449
rect 27709 8483 27767 8489
rect 27709 8449 27721 8483
rect 27755 8480 27767 8483
rect 27798 8480 27804 8492
rect 27755 8452 27804 8480
rect 27755 8449 27767 8452
rect 27709 8443 27767 8449
rect 27632 8412 27660 8443
rect 27798 8440 27804 8452
rect 27856 8440 27862 8492
rect 27908 8489 27936 8520
rect 27893 8483 27951 8489
rect 27893 8449 27905 8483
rect 27939 8480 27951 8483
rect 28353 8483 28411 8489
rect 28353 8480 28365 8483
rect 27939 8452 28365 8480
rect 27939 8449 27951 8452
rect 27893 8443 27951 8449
rect 28353 8449 28365 8452
rect 28399 8449 28411 8483
rect 28534 8480 28540 8492
rect 28495 8452 28540 8480
rect 28353 8443 28411 8449
rect 28534 8440 28540 8452
rect 28592 8440 28598 8492
rect 28736 8489 28764 8588
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 30006 8616 30012 8628
rect 29967 8588 30012 8616
rect 30006 8576 30012 8588
rect 30064 8576 30070 8628
rect 28902 8508 28908 8560
rect 28960 8548 28966 8560
rect 29641 8551 29699 8557
rect 29641 8548 29653 8551
rect 28960 8520 29653 8548
rect 28960 8508 28966 8520
rect 29641 8517 29653 8520
rect 29687 8517 29699 8551
rect 29641 8511 29699 8517
rect 29733 8551 29791 8557
rect 29733 8517 29745 8551
rect 29779 8548 29791 8551
rect 32122 8548 32128 8560
rect 29779 8520 32128 8548
rect 29779 8517 29791 8520
rect 29733 8511 29791 8517
rect 32122 8508 32128 8520
rect 32180 8508 32186 8560
rect 35986 8548 35992 8560
rect 34624 8520 35992 8548
rect 28629 8483 28687 8489
rect 28629 8449 28641 8483
rect 28675 8449 28687 8483
rect 28629 8443 28687 8449
rect 28721 8483 28779 8489
rect 28721 8449 28733 8483
rect 28767 8449 28779 8483
rect 28721 8443 28779 8449
rect 27982 8412 27988 8424
rect 24820 8384 27988 8412
rect 24820 8372 24826 8384
rect 27982 8372 27988 8384
rect 28040 8412 28046 8424
rect 28644 8412 28672 8443
rect 28810 8440 28816 8492
rect 28868 8480 28874 8492
rect 29457 8483 29515 8489
rect 29457 8480 29469 8483
rect 28868 8452 29469 8480
rect 28868 8440 28874 8452
rect 29457 8449 29469 8452
rect 29503 8449 29515 8483
rect 29457 8443 29515 8449
rect 29546 8440 29552 8492
rect 29604 8480 29610 8492
rect 29825 8483 29883 8489
rect 29825 8480 29837 8483
rect 29604 8452 29837 8480
rect 29604 8440 29610 8452
rect 29825 8449 29837 8452
rect 29871 8449 29883 8483
rect 34514 8480 34520 8492
rect 29825 8443 29883 8449
rect 33704 8452 34520 8480
rect 28040 8384 28672 8412
rect 28040 8372 28046 8384
rect 8386 8344 8392 8356
rect 5644 8316 5948 8344
rect 6196 8316 7512 8344
rect 8347 8316 8392 8344
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 2832 8248 2877 8276
rect 2832 8236 2838 8248
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 5644 8276 5672 8316
rect 5810 8276 5816 8288
rect 4120 8248 5672 8276
rect 5771 8248 5816 8276
rect 4120 8236 4126 8248
rect 5810 8236 5816 8248
rect 5868 8236 5874 8288
rect 5920 8276 5948 8316
rect 8386 8304 8392 8316
rect 8444 8304 8450 8356
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 10410 8344 10416 8356
rect 10367 8316 10416 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 6914 8276 6920 8288
rect 5920 8248 6920 8276
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 9214 8236 9220 8288
rect 9272 8276 9278 8288
rect 10336 8276 10364 8307
rect 10410 8304 10416 8316
rect 10468 8344 10474 8356
rect 17313 8347 17371 8353
rect 10468 8316 11008 8344
rect 10468 8304 10474 8316
rect 9272 8248 10364 8276
rect 10980 8276 11008 8316
rect 17313 8313 17325 8347
rect 17359 8344 17371 8347
rect 18782 8344 18788 8356
rect 17359 8316 18788 8344
rect 17359 8313 17371 8316
rect 17313 8307 17371 8313
rect 18782 8304 18788 8316
rect 18840 8304 18846 8356
rect 19150 8304 19156 8356
rect 19208 8344 19214 8356
rect 24670 8344 24676 8356
rect 19208 8316 24676 8344
rect 19208 8304 19214 8316
rect 24670 8304 24676 8316
rect 24728 8304 24734 8356
rect 25222 8304 25228 8356
rect 25280 8344 25286 8356
rect 27154 8344 27160 8356
rect 25280 8316 27160 8344
rect 25280 8304 25286 8316
rect 27154 8304 27160 8316
rect 27212 8304 27218 8356
rect 27249 8347 27307 8353
rect 27249 8313 27261 8347
rect 27295 8344 27307 8347
rect 27706 8344 27712 8356
rect 27295 8316 27712 8344
rect 27295 8313 27307 8316
rect 27249 8307 27307 8313
rect 27706 8304 27712 8316
rect 27764 8304 27770 8356
rect 27890 8304 27896 8356
rect 27948 8344 27954 8356
rect 33704 8353 33732 8452
rect 34514 8440 34520 8452
rect 34572 8440 34578 8492
rect 34624 8489 34652 8520
rect 35986 8508 35992 8520
rect 36044 8508 36050 8560
rect 34609 8483 34667 8489
rect 34609 8449 34621 8483
rect 34655 8449 34667 8483
rect 34609 8443 34667 8449
rect 34698 8440 34704 8492
rect 34756 8480 34762 8492
rect 34885 8483 34943 8489
rect 34756 8452 34801 8480
rect 34756 8440 34762 8452
rect 34885 8449 34897 8483
rect 34931 8480 34943 8483
rect 35618 8480 35624 8492
rect 34931 8452 35624 8480
rect 34931 8449 34943 8452
rect 34885 8443 34943 8449
rect 35618 8440 35624 8452
rect 35676 8440 35682 8492
rect 33689 8347 33747 8353
rect 33689 8344 33701 8347
rect 27948 8316 33701 8344
rect 27948 8304 27954 8316
rect 33689 8313 33701 8316
rect 33735 8313 33747 8347
rect 33689 8307 33747 8313
rect 11885 8279 11943 8285
rect 11885 8276 11897 8279
rect 10980 8248 11897 8276
rect 9272 8236 9278 8248
rect 11885 8245 11897 8248
rect 11931 8245 11943 8279
rect 11885 8239 11943 8245
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 12434 8276 12440 8288
rect 12032 8248 12440 8276
rect 12032 8236 12038 8248
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 22002 8276 22008 8288
rect 15620 8248 22008 8276
rect 15620 8236 15626 8248
rect 22002 8236 22008 8248
rect 22060 8236 22066 8288
rect 22094 8236 22100 8288
rect 22152 8276 22158 8288
rect 26329 8279 26387 8285
rect 26329 8276 26341 8279
rect 22152 8248 26341 8276
rect 22152 8236 22158 8248
rect 26329 8245 26341 8248
rect 26375 8276 26387 8279
rect 27430 8276 27436 8288
rect 26375 8248 27436 8276
rect 26375 8245 26387 8248
rect 26329 8239 26387 8245
rect 27430 8236 27436 8248
rect 27488 8276 27494 8288
rect 28074 8276 28080 8288
rect 27488 8248 28080 8276
rect 27488 8236 27494 8248
rect 28074 8236 28080 8248
rect 28132 8236 28138 8288
rect 34238 8276 34244 8288
rect 34199 8248 34244 8276
rect 34238 8236 34244 8248
rect 34296 8236 34302 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 3881 8075 3939 8081
rect 3881 8072 3893 8075
rect 2424 8044 3893 8072
rect 1578 7896 1584 7948
rect 1636 7936 1642 7948
rect 2424 7945 2452 8044
rect 3881 8041 3893 8044
rect 3927 8072 3939 8075
rect 4062 8072 4068 8084
rect 3927 8044 4068 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 9950 8072 9956 8084
rect 5592 8044 9956 8072
rect 5592 8032 5598 8044
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 13262 8072 13268 8084
rect 10796 8044 12756 8072
rect 13223 8044 13268 8072
rect 6454 8004 6460 8016
rect 3160 7976 6460 8004
rect 2409 7939 2467 7945
rect 2409 7936 2421 7939
rect 1636 7908 2421 7936
rect 1636 7896 1642 7908
rect 2409 7905 2421 7908
rect 2455 7905 2467 7939
rect 2409 7899 2467 7905
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2774 7868 2780 7880
rect 2639 7840 2780 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 1949 7803 2007 7809
rect 1949 7769 1961 7803
rect 1995 7800 2007 7803
rect 2866 7800 2872 7812
rect 1995 7772 2872 7800
rect 1995 7769 2007 7772
rect 1949 7763 2007 7769
rect 2866 7760 2872 7772
rect 2924 7800 2930 7812
rect 3160 7800 3188 7976
rect 6454 7964 6460 7976
rect 6512 7964 6518 8016
rect 3326 7896 3332 7948
rect 3384 7936 3390 7948
rect 5353 7939 5411 7945
rect 5353 7936 5365 7939
rect 3384 7908 5365 7936
rect 3384 7896 3390 7908
rect 5353 7905 5365 7908
rect 5399 7905 5411 7939
rect 5810 7936 5816 7948
rect 5771 7908 5816 7936
rect 5353 7899 5411 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7936 6607 7939
rect 6730 7936 6736 7948
rect 6595 7908 6736 7936
rect 6595 7905 6607 7908
rect 6549 7899 6607 7905
rect 6730 7896 6736 7908
rect 6788 7896 6794 7948
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5537 7871 5595 7877
rect 5537 7868 5549 7871
rect 4764 7840 5549 7868
rect 4764 7828 4770 7840
rect 5537 7837 5549 7840
rect 5583 7837 5595 7871
rect 5718 7868 5724 7880
rect 5679 7840 5724 7868
rect 5537 7831 5595 7837
rect 5718 7828 5724 7840
rect 5776 7828 5782 7880
rect 5902 7868 5908 7880
rect 5863 7840 5908 7868
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6086 7868 6092 7880
rect 6047 7840 6092 7868
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 2924 7772 3188 7800
rect 2924 7760 2930 7772
rect 3234 7760 3240 7812
rect 3292 7800 3298 7812
rect 3970 7800 3976 7812
rect 3292 7772 3976 7800
rect 3292 7760 3298 7772
rect 3970 7760 3976 7772
rect 4028 7800 4034 7812
rect 6932 7800 6960 7831
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 7064 7840 7109 7868
rect 7064 7828 7070 7840
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 10796 7877 10824 8044
rect 11606 8004 11612 8016
rect 10980 7976 11612 8004
rect 10980 7877 11008 7976
rect 11606 7964 11612 7976
rect 11664 7964 11670 8016
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 11204 7908 12357 7936
rect 11204 7896 11210 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 12434 7896 12440 7948
rect 12492 7936 12498 7948
rect 12492 7908 12537 7936
rect 12492 7896 12498 7908
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 9548 7840 10793 7868
rect 9548 7828 9554 7840
rect 10781 7837 10793 7840
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 10965 7871 11023 7877
rect 10965 7837 10977 7871
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11057 7871 11115 7877
rect 11057 7837 11069 7871
rect 11103 7837 11115 7871
rect 11057 7831 11115 7837
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 8297 7803 8355 7809
rect 8297 7800 8309 7803
rect 4028 7772 6960 7800
rect 7024 7772 8309 7800
rect 4028 7760 4034 7772
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 4433 7735 4491 7741
rect 2832 7704 2877 7732
rect 2832 7692 2838 7704
rect 4433 7701 4445 7735
rect 4479 7732 4491 7735
rect 5810 7732 5816 7744
rect 4479 7704 5816 7732
rect 4479 7701 4491 7704
rect 4433 7695 4491 7701
rect 5810 7692 5816 7704
rect 5868 7692 5874 7744
rect 6178 7692 6184 7744
rect 6236 7732 6242 7744
rect 7024 7732 7052 7772
rect 8297 7769 8309 7772
rect 8343 7769 8355 7803
rect 8297 7763 8355 7769
rect 8386 7760 8392 7812
rect 8444 7800 8450 7812
rect 11072 7800 11100 7831
rect 11238 7800 11244 7812
rect 8444 7772 9674 7800
rect 11072 7772 11244 7800
rect 8444 7760 8450 7772
rect 7190 7732 7196 7744
rect 6236 7704 7052 7732
rect 7151 7704 7196 7732
rect 6236 7692 6242 7704
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 7742 7732 7748 7744
rect 7703 7704 7748 7732
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8536 7704 8953 7732
rect 8536 7692 8542 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 9646 7732 9674 7772
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 11348 7800 11376 7831
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12161 7871 12219 7877
rect 12161 7868 12173 7871
rect 12032 7840 12173 7868
rect 12032 7828 12038 7840
rect 12161 7837 12173 7840
rect 12207 7837 12219 7871
rect 12526 7868 12532 7880
rect 12487 7840 12532 7868
rect 12161 7831 12219 7837
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 12728 7877 12756 8044
rect 13262 8032 13268 8044
rect 13320 8032 13326 8084
rect 15010 8032 15016 8084
rect 15068 8072 15074 8084
rect 16025 8075 16083 8081
rect 16025 8072 16037 8075
rect 15068 8044 16037 8072
rect 15068 8032 15074 8044
rect 16025 8041 16037 8044
rect 16071 8041 16083 8075
rect 16025 8035 16083 8041
rect 17865 8075 17923 8081
rect 17865 8041 17877 8075
rect 17911 8072 17923 8075
rect 18138 8072 18144 8084
rect 17911 8044 18144 8072
rect 17911 8041 17923 8044
rect 17865 8035 17923 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18325 8075 18383 8081
rect 18325 8041 18337 8075
rect 18371 8072 18383 8075
rect 18506 8072 18512 8084
rect 18371 8044 18512 8072
rect 18371 8041 18383 8044
rect 18325 8035 18383 8041
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 22925 8075 22983 8081
rect 22925 8041 22937 8075
rect 22971 8072 22983 8075
rect 23566 8072 23572 8084
rect 22971 8044 23572 8072
rect 22971 8041 22983 8044
rect 22925 8035 22983 8041
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 28718 8032 28724 8084
rect 28776 8072 28782 8084
rect 28813 8075 28871 8081
rect 28813 8072 28825 8075
rect 28776 8044 28825 8072
rect 28776 8032 28782 8044
rect 28813 8041 28825 8044
rect 28859 8041 28871 8075
rect 34698 8072 34704 8084
rect 34659 8044 34704 8072
rect 28813 8035 28871 8041
rect 34698 8032 34704 8044
rect 34756 8032 34762 8084
rect 14553 8007 14611 8013
rect 14553 7973 14565 8007
rect 14599 8004 14611 8007
rect 19242 8004 19248 8016
rect 14599 7976 19248 8004
rect 14599 7973 14611 7976
rect 14553 7967 14611 7973
rect 19242 7964 19248 7976
rect 19300 7964 19306 8016
rect 34149 8007 34207 8013
rect 34149 7973 34161 8007
rect 34195 8004 34207 8007
rect 34790 8004 34796 8016
rect 34195 7976 34796 8004
rect 34195 7973 34207 7976
rect 34149 7967 34207 7973
rect 34790 7964 34796 7976
rect 34848 7964 34854 8016
rect 37366 7964 37372 8016
rect 37424 7964 37430 8016
rect 17126 7896 17132 7948
rect 17184 7936 17190 7948
rect 32766 7936 32772 7948
rect 17184 7908 22094 7936
rect 32727 7908 32772 7936
rect 17184 7896 17190 7908
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 13964 7840 14749 7868
rect 13964 7828 13970 7840
rect 14737 7837 14749 7840
rect 14783 7868 14795 7871
rect 15102 7868 15108 7880
rect 14783 7840 15108 7868
rect 14783 7837 14795 7840
rect 14737 7831 14795 7837
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 15286 7868 15292 7880
rect 15247 7840 15292 7868
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7868 18567 7871
rect 18598 7868 18604 7880
rect 18555 7840 18604 7868
rect 18555 7837 18567 7840
rect 18509 7831 18567 7837
rect 18598 7828 18604 7840
rect 18656 7828 18662 7880
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 19521 7871 19579 7877
rect 19521 7837 19533 7871
rect 19567 7868 19579 7871
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19567 7840 20085 7868
rect 19567 7837 19579 7840
rect 19521 7831 19579 7837
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 22066 7868 22094 7908
rect 32766 7896 32772 7908
rect 32824 7896 32830 7948
rect 22373 7871 22431 7877
rect 22373 7868 22385 7871
rect 22066 7840 22385 7868
rect 20073 7831 20131 7837
rect 22373 7837 22385 7840
rect 22419 7837 22431 7871
rect 22554 7868 22560 7880
rect 22515 7840 22560 7868
rect 22373 7831 22431 7837
rect 12618 7800 12624 7812
rect 11348 7772 12624 7800
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 18322 7800 18328 7812
rect 17236 7772 18328 7800
rect 17236 7744 17264 7772
rect 18322 7760 18328 7772
rect 18380 7760 18386 7812
rect 18693 7803 18751 7809
rect 18693 7769 18705 7803
rect 18739 7769 18751 7803
rect 18693 7763 18751 7769
rect 11146 7732 11152 7744
rect 9646 7704 11152 7732
rect 8941 7695 8999 7701
rect 11146 7692 11152 7704
rect 11204 7692 11210 7744
rect 11514 7732 11520 7744
rect 11475 7704 11520 7732
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 11977 7735 12035 7741
rect 11977 7701 11989 7735
rect 12023 7732 12035 7735
rect 12802 7732 12808 7744
rect 12023 7704 12808 7732
rect 12023 7701 12035 7704
rect 11977 7695 12035 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 14424 7704 15485 7732
rect 14424 7692 14430 7704
rect 15473 7701 15485 7704
rect 15519 7732 15531 7735
rect 15562 7732 15568 7744
rect 15519 7704 15568 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 17218 7732 17224 7744
rect 17179 7704 17224 7732
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 18708 7732 18736 7763
rect 18782 7760 18788 7812
rect 18840 7800 18846 7812
rect 19536 7800 19564 7831
rect 22554 7828 22560 7840
rect 22612 7828 22618 7880
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7868 22799 7871
rect 23474 7868 23480 7880
rect 22787 7840 23480 7868
rect 22787 7837 22799 7840
rect 22741 7831 22799 7837
rect 23474 7828 23480 7840
rect 23532 7828 23538 7880
rect 27062 7828 27068 7880
rect 27120 7868 27126 7880
rect 27433 7871 27491 7877
rect 27433 7868 27445 7871
rect 27120 7840 27445 7868
rect 27120 7828 27126 7840
rect 27433 7837 27445 7840
rect 27479 7868 27491 7871
rect 29822 7868 29828 7880
rect 27479 7840 29828 7868
rect 27479 7837 27491 7840
rect 27433 7831 27491 7837
rect 29822 7828 29828 7840
rect 29880 7828 29886 7880
rect 33036 7871 33094 7877
rect 33036 7837 33048 7871
rect 33082 7868 33094 7871
rect 34238 7868 34244 7880
rect 33082 7840 34244 7868
rect 33082 7837 33094 7840
rect 33036 7831 33094 7837
rect 34238 7828 34244 7840
rect 34296 7828 34302 7880
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 34885 7871 34943 7877
rect 34885 7868 34897 7871
rect 34848 7840 34897 7868
rect 34848 7828 34854 7840
rect 34885 7837 34897 7840
rect 34931 7837 34943 7871
rect 34885 7831 34943 7837
rect 35069 7871 35127 7877
rect 35069 7837 35081 7871
rect 35115 7868 35127 7871
rect 35342 7868 35348 7880
rect 35115 7840 35348 7868
rect 35115 7837 35127 7840
rect 35069 7831 35127 7837
rect 35342 7828 35348 7840
rect 35400 7868 35406 7880
rect 35526 7868 35532 7880
rect 35400 7840 35532 7868
rect 35400 7828 35406 7840
rect 35526 7828 35532 7840
rect 35584 7828 35590 7880
rect 37182 7868 37188 7880
rect 37143 7840 37188 7868
rect 37182 7828 37188 7840
rect 37240 7828 37246 7880
rect 37384 7877 37412 7964
rect 37734 7936 37740 7948
rect 37476 7908 37740 7936
rect 37476 7877 37504 7908
rect 37734 7896 37740 7908
rect 37792 7896 37798 7948
rect 37348 7871 37412 7877
rect 37348 7837 37360 7871
rect 37394 7840 37412 7871
rect 37461 7871 37519 7877
rect 37394 7837 37406 7840
rect 37348 7831 37406 7837
rect 37461 7837 37473 7871
rect 37507 7837 37519 7871
rect 37461 7831 37519 7837
rect 37599 7871 37657 7877
rect 37599 7837 37611 7871
rect 37645 7868 37657 7871
rect 58158 7868 58164 7880
rect 37645 7840 37767 7868
rect 58119 7840 58164 7868
rect 37645 7837 37657 7840
rect 37599 7831 37657 7837
rect 18840 7772 19564 7800
rect 22649 7803 22707 7809
rect 18840 7760 18846 7772
rect 22649 7769 22661 7803
rect 22695 7800 22707 7803
rect 24946 7800 24952 7812
rect 22695 7772 24952 7800
rect 22695 7769 22707 7772
rect 22649 7763 22707 7769
rect 24946 7760 24952 7772
rect 25004 7800 25010 7812
rect 25682 7800 25688 7812
rect 25004 7772 25688 7800
rect 25004 7760 25010 7772
rect 25682 7760 25688 7772
rect 25740 7760 25746 7812
rect 27706 7809 27712 7812
rect 27700 7800 27712 7809
rect 27667 7772 27712 7800
rect 27700 7763 27712 7772
rect 27706 7760 27712 7763
rect 27764 7760 27770 7812
rect 36725 7803 36783 7809
rect 36725 7800 36737 7803
rect 35866 7772 36737 7800
rect 19242 7732 19248 7744
rect 18708 7704 19248 7732
rect 19242 7692 19248 7704
rect 19300 7692 19306 7744
rect 23290 7692 23296 7744
rect 23348 7732 23354 7744
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 23348 7704 23489 7732
rect 23348 7692 23354 7704
rect 23477 7701 23489 7704
rect 23523 7732 23535 7735
rect 25958 7732 25964 7744
rect 23523 7704 25964 7732
rect 23523 7701 23535 7704
rect 23477 7695 23535 7701
rect 25958 7692 25964 7704
rect 26016 7732 26022 7744
rect 33778 7732 33784 7744
rect 26016 7704 33784 7732
rect 26016 7692 26022 7704
rect 33778 7692 33784 7704
rect 33836 7732 33842 7744
rect 35866 7732 35894 7772
rect 36725 7769 36737 7772
rect 36771 7800 36783 7803
rect 37739 7800 37767 7840
rect 58158 7828 58164 7840
rect 58216 7828 58222 7880
rect 36771 7772 37767 7800
rect 36771 7769 36783 7772
rect 36725 7763 36783 7769
rect 37826 7732 37832 7744
rect 33836 7704 35894 7732
rect 37787 7704 37832 7732
rect 33836 7692 33842 7704
rect 37826 7692 37832 7704
rect 37884 7692 37890 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 3789 7531 3847 7537
rect 3789 7497 3801 7531
rect 3835 7528 3847 7531
rect 3970 7528 3976 7540
rect 3835 7500 3976 7528
rect 3835 7497 3847 7500
rect 3789 7491 3847 7497
rect 3970 7488 3976 7500
rect 4028 7488 4034 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 7926 7528 7932 7540
rect 5859 7500 7932 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 12158 7528 12164 7540
rect 11112 7500 12164 7528
rect 11112 7488 11118 7500
rect 12158 7488 12164 7500
rect 12216 7488 12222 7540
rect 19426 7528 19432 7540
rect 12406 7500 13768 7528
rect 5902 7420 5908 7472
rect 5960 7460 5966 7472
rect 6457 7463 6515 7469
rect 6457 7460 6469 7463
rect 5960 7432 6469 7460
rect 5960 7420 5966 7432
rect 6457 7429 6469 7432
rect 6503 7460 6515 7463
rect 11606 7460 11612 7472
rect 6503 7432 8432 7460
rect 11567 7432 11612 7460
rect 6503 7429 6515 7432
rect 6457 7423 6515 7429
rect 2130 7352 2136 7404
rect 2188 7392 2194 7404
rect 2682 7401 2688 7404
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 2188 7364 2421 7392
rect 2188 7352 2194 7364
rect 2409 7361 2421 7364
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2676 7355 2688 7401
rect 2740 7392 2746 7404
rect 2740 7364 2776 7392
rect 2682 7352 2688 7355
rect 2740 7352 2746 7364
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 8306 7395 8364 7401
rect 8306 7392 8318 7395
rect 7892 7364 8318 7392
rect 7892 7352 7898 7364
rect 8306 7361 8318 7364
rect 8352 7361 8364 7395
rect 8404 7392 8432 7432
rect 11606 7420 11612 7432
rect 11664 7420 11670 7472
rect 12406 7460 12434 7500
rect 11716 7432 12434 7460
rect 12713 7463 12771 7469
rect 11716 7392 11744 7432
rect 12713 7429 12725 7463
rect 12759 7429 12771 7463
rect 12713 7423 12771 7429
rect 12728 7392 12756 7423
rect 8404 7364 11744 7392
rect 12406 7364 12756 7392
rect 8306 7355 8364 7361
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7324 8631 7327
rect 11238 7324 11244 7336
rect 8619 7296 11244 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 11238 7284 11244 7296
rect 11296 7284 11302 7336
rect 12158 7216 12164 7268
rect 12216 7256 12222 7268
rect 12406 7256 12434 7364
rect 12216 7228 12434 7256
rect 12728 7256 12756 7364
rect 13740 7324 13768 7500
rect 19168 7500 19432 7528
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7392 14522 7404
rect 14918 7392 14924 7404
rect 14516 7364 14924 7392
rect 14516 7352 14522 7364
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 16758 7352 16764 7404
rect 16816 7392 16822 7404
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 16816 7364 16865 7392
rect 16816 7352 16822 7364
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 17034 7392 17040 7404
rect 16995 7364 17040 7392
rect 16853 7355 16911 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 19168 7401 19196 7500
rect 19426 7488 19432 7500
rect 19484 7528 19490 7540
rect 21266 7528 21272 7540
rect 19484 7500 21036 7528
rect 21227 7500 21272 7528
rect 19484 7488 19490 7500
rect 20806 7460 20812 7472
rect 19904 7432 20812 7460
rect 19904 7401 19932 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 21008 7460 21036 7500
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 22554 7528 22560 7540
rect 22388 7500 22560 7528
rect 22388 7469 22416 7500
rect 22554 7488 22560 7500
rect 22612 7488 22618 7540
rect 22741 7531 22799 7537
rect 22741 7497 22753 7531
rect 22787 7528 22799 7531
rect 24578 7528 24584 7540
rect 22787 7500 24584 7528
rect 22787 7497 22799 7500
rect 22741 7491 22799 7497
rect 24578 7488 24584 7500
rect 24636 7488 24642 7540
rect 24762 7488 24768 7540
rect 24820 7488 24826 7540
rect 27798 7488 27804 7540
rect 27856 7528 27862 7540
rect 28353 7531 28411 7537
rect 28353 7528 28365 7531
rect 27856 7500 28365 7528
rect 27856 7488 27862 7500
rect 28353 7497 28365 7500
rect 28399 7497 28411 7531
rect 34422 7528 34428 7540
rect 34383 7500 34428 7528
rect 28353 7491 28411 7497
rect 34422 7488 34428 7500
rect 34480 7488 34486 7540
rect 34790 7488 34796 7540
rect 34848 7528 34854 7540
rect 35802 7528 35808 7540
rect 34848 7500 35808 7528
rect 34848 7488 34854 7500
rect 35802 7488 35808 7500
rect 35860 7488 35866 7540
rect 37366 7488 37372 7540
rect 37424 7528 37430 7540
rect 38749 7531 38807 7537
rect 38749 7528 38761 7531
rect 37424 7500 38761 7528
rect 37424 7488 37430 7500
rect 38749 7497 38761 7500
rect 38795 7497 38807 7531
rect 38749 7491 38807 7497
rect 22373 7463 22431 7469
rect 22373 7460 22385 7463
rect 21008 7432 22385 7460
rect 22373 7429 22385 7432
rect 22419 7429 22431 7463
rect 22373 7423 22431 7429
rect 23290 7420 23296 7472
rect 23348 7460 23354 7472
rect 24780 7460 24808 7488
rect 23348 7432 23520 7460
rect 23348 7420 23354 7432
rect 19153 7395 19211 7401
rect 19153 7361 19165 7395
rect 19199 7361 19211 7395
rect 19153 7355 19211 7361
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 19978 7352 19984 7404
rect 20036 7392 20042 7404
rect 20145 7395 20203 7401
rect 20145 7392 20157 7395
rect 20036 7364 20157 7392
rect 20036 7352 20042 7364
rect 20145 7361 20157 7364
rect 20191 7361 20203 7395
rect 20145 7355 20203 7361
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 22189 7395 22247 7401
rect 22189 7392 22201 7395
rect 20772 7364 22201 7392
rect 20772 7352 20778 7364
rect 22189 7361 22201 7364
rect 22235 7361 22247 7395
rect 22189 7355 22247 7361
rect 22465 7395 22523 7401
rect 22465 7361 22477 7395
rect 22511 7361 22523 7395
rect 22465 7355 22523 7361
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7392 22615 7395
rect 23382 7392 23388 7404
rect 22603 7364 23388 7392
rect 22603 7361 22615 7364
rect 22557 7355 22615 7361
rect 17402 7324 17408 7336
rect 13740 7296 17408 7324
rect 17402 7284 17408 7296
rect 17460 7284 17466 7336
rect 19426 7324 19432 7336
rect 19387 7296 19432 7324
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 18046 7256 18052 7268
rect 12728 7228 18052 7256
rect 12216 7216 12222 7228
rect 18046 7216 18052 7228
rect 18104 7216 18110 7268
rect 22480 7256 22508 7355
rect 23382 7352 23388 7364
rect 23440 7352 23446 7404
rect 23492 7401 23520 7432
rect 24688 7432 24808 7460
rect 24688 7404 24716 7432
rect 24854 7420 24860 7472
rect 24912 7460 24918 7472
rect 25501 7463 25559 7469
rect 25501 7460 25513 7463
rect 24912 7432 25513 7460
rect 24912 7420 24918 7432
rect 25501 7429 25513 7432
rect 25547 7429 25559 7463
rect 25682 7460 25688 7472
rect 25643 7432 25688 7460
rect 25501 7423 25559 7429
rect 25682 7420 25688 7432
rect 25740 7420 25746 7472
rect 26786 7420 26792 7472
rect 26844 7460 26850 7472
rect 27065 7463 27123 7469
rect 27065 7460 27077 7463
rect 26844 7432 27077 7460
rect 26844 7420 26850 7432
rect 27065 7429 27077 7432
rect 27111 7460 27123 7463
rect 31018 7460 31024 7472
rect 27111 7432 31024 7460
rect 27111 7429 27123 7432
rect 27065 7423 27123 7429
rect 31018 7420 31024 7432
rect 31076 7460 31082 7472
rect 31481 7463 31539 7469
rect 31481 7460 31493 7463
rect 31076 7432 31493 7460
rect 31076 7420 31082 7432
rect 31481 7429 31493 7432
rect 31527 7460 31539 7463
rect 34054 7460 34060 7472
rect 31527 7432 34060 7460
rect 31527 7429 31539 7432
rect 31481 7423 31539 7429
rect 34054 7420 34060 7432
rect 34112 7420 34118 7472
rect 35434 7460 35440 7472
rect 34624 7432 35440 7460
rect 23477 7395 23535 7401
rect 23477 7361 23489 7395
rect 23523 7361 23535 7395
rect 23477 7355 23535 7361
rect 23566 7395 23624 7401
rect 23566 7361 23578 7395
rect 23612 7361 23624 7395
rect 23566 7355 23624 7361
rect 23198 7284 23204 7336
rect 23256 7324 23262 7336
rect 23584 7324 23612 7355
rect 23658 7352 23664 7404
rect 23716 7392 23722 7404
rect 23845 7395 23903 7401
rect 23716 7364 23761 7392
rect 23716 7352 23722 7364
rect 23845 7361 23857 7395
rect 23891 7392 23903 7395
rect 24394 7392 24400 7404
rect 23891 7364 24400 7392
rect 23891 7361 23903 7364
rect 23845 7355 23903 7361
rect 24394 7352 24400 7364
rect 24452 7352 24458 7404
rect 24486 7352 24492 7404
rect 24544 7401 24550 7404
rect 24544 7395 24593 7401
rect 24544 7361 24547 7395
rect 24581 7361 24593 7395
rect 24544 7355 24593 7361
rect 24670 7398 24728 7404
rect 24670 7364 24682 7398
rect 24716 7364 24728 7398
rect 24670 7358 24728 7364
rect 24544 7352 24550 7355
rect 24762 7352 24768 7404
rect 24820 7401 24826 7404
rect 24820 7392 24828 7401
rect 24949 7395 25007 7401
rect 24820 7364 24865 7392
rect 24820 7355 24828 7364
rect 24949 7361 24961 7395
rect 24995 7392 25007 7395
rect 25222 7392 25228 7404
rect 24995 7364 25228 7392
rect 24995 7361 25007 7364
rect 24949 7355 25007 7361
rect 24820 7352 24826 7355
rect 23256 7296 23612 7324
rect 23256 7284 23262 7296
rect 23474 7256 23480 7268
rect 22480 7228 23480 7256
rect 23474 7216 23480 7228
rect 23532 7216 23538 7268
rect 23658 7216 23664 7268
rect 23716 7256 23722 7268
rect 24854 7256 24860 7268
rect 23716 7228 24860 7256
rect 23716 7216 23722 7228
rect 24854 7216 24860 7228
rect 24912 7216 24918 7268
rect 1946 7188 1952 7200
rect 1907 7160 1952 7188
rect 1946 7148 1952 7160
rect 2004 7148 2010 7200
rect 4798 7188 4804 7200
rect 4759 7160 4804 7188
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 7193 7191 7251 7197
rect 7193 7157 7205 7191
rect 7239 7188 7251 7191
rect 7650 7188 7656 7200
rect 7239 7160 7656 7188
rect 7239 7157 7251 7160
rect 7193 7151 7251 7157
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 9398 7188 9404 7200
rect 9359 7160 9404 7188
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9582 7148 9588 7200
rect 9640 7188 9646 7200
rect 9861 7191 9919 7197
rect 9861 7188 9873 7191
rect 9640 7160 9873 7188
rect 9640 7148 9646 7160
rect 9861 7157 9873 7160
rect 9907 7157 9919 7191
rect 9861 7151 9919 7157
rect 14642 7148 14648 7200
rect 14700 7188 14706 7200
rect 15105 7191 15163 7197
rect 15105 7188 15117 7191
rect 14700 7160 15117 7188
rect 14700 7148 14706 7160
rect 15105 7157 15117 7160
rect 15151 7188 15163 7191
rect 15286 7188 15292 7200
rect 15151 7160 15292 7188
rect 15151 7157 15163 7160
rect 15105 7151 15163 7157
rect 15286 7148 15292 7160
rect 15344 7148 15350 7200
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 15896 7160 16681 7188
rect 15896 7148 15902 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 23201 7191 23259 7197
rect 23201 7157 23213 7191
rect 23247 7188 23259 7191
rect 23566 7188 23572 7200
rect 23247 7160 23572 7188
rect 23247 7157 23259 7160
rect 23201 7151 23259 7157
rect 23566 7148 23572 7160
rect 23624 7148 23630 7200
rect 24210 7148 24216 7200
rect 24268 7188 24274 7200
rect 24305 7191 24363 7197
rect 24305 7188 24317 7191
rect 24268 7160 24317 7188
rect 24268 7148 24274 7160
rect 24305 7157 24317 7160
rect 24351 7157 24363 7191
rect 24305 7151 24363 7157
rect 24394 7148 24400 7200
rect 24452 7188 24458 7200
rect 24964 7188 24992 7355
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 25866 7392 25872 7404
rect 25827 7364 25872 7392
rect 25866 7352 25872 7364
rect 25924 7392 25930 7404
rect 26142 7392 26148 7404
rect 25924 7364 26148 7392
rect 25924 7352 25930 7364
rect 26142 7352 26148 7364
rect 26200 7392 26206 7404
rect 27985 7395 28043 7401
rect 27985 7392 27997 7395
rect 26200 7364 27997 7392
rect 26200 7352 26206 7364
rect 27985 7361 27997 7364
rect 28031 7361 28043 7395
rect 27985 7355 28043 7361
rect 28169 7395 28227 7401
rect 28169 7361 28181 7395
rect 28215 7392 28227 7395
rect 28718 7392 28724 7404
rect 28215 7364 28724 7392
rect 28215 7361 28227 7364
rect 28169 7355 28227 7361
rect 28718 7352 28724 7364
rect 28776 7352 28782 7404
rect 34624 7401 34652 7432
rect 35434 7420 35440 7432
rect 35492 7420 35498 7472
rect 35713 7463 35771 7469
rect 35713 7429 35725 7463
rect 35759 7460 35771 7463
rect 37182 7460 37188 7472
rect 35759 7432 37188 7460
rect 35759 7429 35771 7432
rect 35713 7423 35771 7429
rect 37182 7420 37188 7432
rect 37240 7420 37246 7472
rect 34609 7395 34667 7401
rect 34609 7361 34621 7395
rect 34655 7361 34667 7395
rect 34609 7355 34667 7361
rect 34701 7395 34759 7401
rect 34701 7361 34713 7395
rect 34747 7361 34759 7395
rect 34701 7355 34759 7361
rect 34716 7324 34744 7355
rect 34790 7352 34796 7404
rect 34848 7392 34854 7404
rect 34977 7395 35035 7401
rect 34848 7364 34893 7392
rect 34848 7352 34854 7364
rect 34977 7361 34989 7395
rect 35023 7392 35035 7395
rect 35342 7392 35348 7404
rect 35023 7364 35348 7392
rect 35023 7361 35035 7364
rect 34977 7355 35035 7361
rect 35342 7352 35348 7364
rect 35400 7352 35406 7404
rect 35452 7392 35480 7420
rect 35621 7395 35679 7401
rect 35621 7392 35633 7395
rect 35452 7364 35633 7392
rect 35621 7361 35633 7364
rect 35667 7361 35679 7395
rect 35802 7392 35808 7404
rect 35763 7364 35808 7392
rect 35621 7355 35679 7361
rect 35802 7352 35808 7364
rect 35860 7352 35866 7404
rect 35986 7392 35992 7404
rect 35947 7364 35992 7392
rect 35986 7352 35992 7364
rect 36044 7352 36050 7404
rect 36078 7352 36084 7404
rect 36136 7392 36142 7404
rect 36722 7392 36728 7404
rect 36136 7364 36728 7392
rect 36136 7352 36142 7364
rect 36722 7352 36728 7364
rect 36780 7352 36786 7404
rect 37090 7352 37096 7404
rect 37148 7392 37154 7404
rect 37458 7401 37464 7404
rect 37277 7395 37335 7401
rect 37277 7392 37289 7395
rect 37148 7364 37289 7392
rect 37148 7352 37154 7364
rect 37277 7361 37289 7364
rect 37323 7361 37335 7395
rect 37456 7392 37464 7401
rect 37419 7364 37464 7392
rect 37277 7355 37335 7361
rect 37456 7355 37464 7364
rect 37458 7352 37464 7355
rect 37516 7352 37522 7404
rect 37572 7395 37630 7401
rect 37572 7361 37584 7395
rect 37618 7361 37630 7395
rect 37572 7355 37630 7361
rect 37691 7395 37749 7401
rect 37691 7361 37703 7395
rect 37737 7392 37749 7395
rect 37918 7392 37924 7404
rect 37737 7364 37924 7392
rect 37737 7361 37749 7364
rect 37691 7355 37749 7361
rect 37587 7324 37615 7355
rect 37918 7352 37924 7364
rect 37976 7352 37982 7404
rect 38378 7392 38384 7404
rect 38339 7364 38384 7392
rect 38378 7352 38384 7364
rect 38436 7352 38442 7404
rect 38565 7395 38623 7401
rect 38565 7361 38577 7395
rect 38611 7361 38623 7395
rect 38565 7355 38623 7361
rect 38580 7324 38608 7355
rect 39114 7324 39120 7336
rect 34716 7296 35894 7324
rect 37587 7296 37780 7324
rect 25130 7216 25136 7268
rect 25188 7256 25194 7268
rect 35437 7259 35495 7265
rect 35437 7256 35449 7259
rect 25188 7228 35449 7256
rect 25188 7216 25194 7228
rect 35437 7225 35449 7228
rect 35483 7225 35495 7259
rect 35437 7219 35495 7225
rect 24452 7160 24992 7188
rect 29733 7191 29791 7197
rect 24452 7148 24458 7160
rect 29733 7157 29745 7191
rect 29779 7188 29791 7191
rect 29822 7188 29828 7200
rect 29779 7160 29828 7188
rect 29779 7157 29791 7160
rect 29733 7151 29791 7157
rect 29822 7148 29828 7160
rect 29880 7188 29886 7200
rect 30190 7188 30196 7200
rect 29880 7160 30196 7188
rect 29880 7148 29886 7160
rect 30190 7148 30196 7160
rect 30248 7148 30254 7200
rect 35866 7188 35894 7296
rect 37752 7268 37780 7296
rect 37844 7296 39120 7324
rect 37734 7216 37740 7268
rect 37792 7216 37798 7268
rect 37844 7188 37872 7296
rect 39114 7284 39120 7296
rect 39172 7284 39178 7336
rect 35866 7160 37872 7188
rect 37921 7191 37979 7197
rect 37921 7157 37933 7191
rect 37967 7188 37979 7191
rect 38010 7188 38016 7200
rect 37967 7160 38016 7188
rect 37967 7157 37979 7160
rect 37921 7151 37979 7157
rect 38010 7148 38016 7160
rect 38068 7148 38074 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 1578 6984 1584 6996
rect 1539 6956 1584 6984
rect 1578 6944 1584 6956
rect 1636 6944 1642 6996
rect 2593 6987 2651 6993
rect 2593 6953 2605 6987
rect 2639 6984 2651 6987
rect 2682 6984 2688 6996
rect 2639 6956 2688 6984
rect 2639 6953 2651 6956
rect 2593 6947 2651 6953
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 20806 6944 20812 6996
rect 20864 6984 20870 6996
rect 20901 6987 20959 6993
rect 20901 6984 20913 6987
rect 20864 6956 20913 6984
rect 20864 6944 20870 6956
rect 20901 6953 20913 6956
rect 20947 6953 20959 6987
rect 20901 6947 20959 6953
rect 22002 6944 22008 6996
rect 22060 6984 22066 6996
rect 24486 6984 24492 6996
rect 22060 6956 24492 6984
rect 22060 6944 22066 6956
rect 24486 6944 24492 6956
rect 24544 6984 24550 6996
rect 27246 6984 27252 6996
rect 24544 6956 27252 6984
rect 24544 6944 24550 6956
rect 27246 6944 27252 6956
rect 27304 6984 27310 6996
rect 36078 6984 36084 6996
rect 27304 6956 36084 6984
rect 27304 6944 27310 6956
rect 36078 6944 36084 6956
rect 36136 6944 36142 6996
rect 9490 6916 9496 6928
rect 7116 6888 9496 6916
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 6086 6848 6092 6860
rect 2464 6820 6092 6848
rect 2464 6808 2470 6820
rect 6086 6808 6092 6820
rect 6144 6808 6150 6860
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 5353 6783 5411 6789
rect 2832 6752 2877 6780
rect 2832 6740 2838 6752
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 6104 6780 6132 6808
rect 7116 6789 7144 6888
rect 9490 6876 9496 6888
rect 9548 6916 9554 6928
rect 9548 6888 9904 6916
rect 9548 6876 9554 6888
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 7377 6851 7435 6857
rect 7377 6848 7389 6851
rect 7248 6820 7389 6848
rect 7248 6808 7254 6820
rect 7377 6817 7389 6820
rect 7423 6817 7435 6851
rect 7377 6811 7435 6817
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7834 6848 7840 6860
rect 7524 6820 7569 6848
rect 7795 6820 7840 6848
rect 7524 6808 7530 6820
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 8018 6808 8024 6860
rect 8076 6848 8082 6860
rect 9876 6857 9904 6888
rect 14918 6876 14924 6928
rect 14976 6916 14982 6928
rect 14976 6888 15792 6916
rect 14976 6876 14982 6888
rect 9861 6851 9919 6857
rect 8076 6820 9076 6848
rect 8076 6808 8082 6820
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 5399 6752 6040 6780
rect 6104 6752 7113 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 6012 6712 6040 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6749 7343 6783
rect 7650 6780 7656 6792
rect 7563 6752 7656 6780
rect 7285 6743 7343 6749
rect 7190 6712 7196 6724
rect 6012 6684 7196 6712
rect 7190 6672 7196 6684
rect 7248 6672 7254 6724
rect 7300 6712 7328 6743
rect 7650 6740 7656 6752
rect 7708 6780 7714 6792
rect 8202 6780 8208 6792
rect 7708 6752 8208 6780
rect 7708 6740 7714 6752
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 7300 6684 8248 6712
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 3050 6644 3056 6656
rect 2179 6616 3056 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3970 6644 3976 6656
rect 3931 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6644 4583 6647
rect 4614 6644 4620 6656
rect 4571 6616 4620 6644
rect 4571 6613 4583 6616
rect 4525 6607 4583 6613
rect 4614 6604 4620 6616
rect 4672 6644 4678 6656
rect 5442 6644 5448 6656
rect 4672 6616 5448 6644
rect 4672 6604 4678 6616
rect 5442 6604 5448 6616
rect 5500 6604 5506 6656
rect 5994 6644 6000 6656
rect 5955 6616 6000 6644
rect 5994 6604 6000 6616
rect 6052 6604 6058 6656
rect 6546 6644 6552 6656
rect 6507 6616 6552 6644
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 8220 6644 8248 6684
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 8941 6715 8999 6721
rect 8941 6712 8953 6715
rect 8720 6684 8953 6712
rect 8720 6672 8726 6684
rect 8941 6681 8953 6684
rect 8987 6681 8999 6715
rect 8941 6675 8999 6681
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 8220 6616 8401 6644
rect 8389 6613 8401 6616
rect 8435 6644 8447 6647
rect 8846 6644 8852 6656
rect 8435 6616 8852 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9048 6644 9076 6820
rect 9861 6817 9873 6851
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 15381 6851 15439 6857
rect 15381 6817 15393 6851
rect 15427 6848 15439 6851
rect 15470 6848 15476 6860
rect 15427 6820 15476 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9585 6783 9643 6789
rect 9585 6780 9597 6783
rect 9548 6752 9597 6780
rect 9548 6740 9554 6752
rect 9585 6749 9597 6752
rect 9631 6749 9643 6783
rect 11238 6780 11244 6792
rect 11151 6752 11244 6780
rect 9585 6743 9643 6749
rect 11238 6740 11244 6752
rect 11296 6780 11302 6792
rect 13078 6780 13084 6792
rect 11296 6752 13084 6780
rect 11296 6740 11302 6752
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 15764 6789 15792 6888
rect 34054 6848 34060 6860
rect 34015 6820 34060 6848
rect 34054 6808 34060 6820
rect 34112 6848 34118 6860
rect 34112 6820 36952 6848
rect 34112 6808 34118 6820
rect 15611 6783 15669 6789
rect 15611 6780 15623 6783
rect 14844 6752 15623 6780
rect 11514 6721 11520 6724
rect 11508 6712 11520 6721
rect 11475 6684 11520 6712
rect 11508 6675 11520 6684
rect 11514 6672 11520 6675
rect 11572 6672 11578 6724
rect 14550 6712 14556 6724
rect 12452 6684 14556 6712
rect 12452 6644 12480 6684
rect 14550 6672 14556 6684
rect 14608 6712 14614 6724
rect 14844 6721 14872 6752
rect 15611 6749 15623 6752
rect 15657 6749 15669 6783
rect 15611 6743 15669 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15838 6740 15844 6792
rect 15896 6780 15902 6792
rect 16025 6783 16083 6789
rect 15896 6752 15941 6780
rect 15896 6740 15902 6752
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 17126 6780 17132 6792
rect 16025 6743 16083 6749
rect 16684 6752 17132 6780
rect 14829 6715 14887 6721
rect 14829 6712 14841 6715
rect 14608 6684 14841 6712
rect 14608 6672 14614 6684
rect 14829 6681 14841 6684
rect 14875 6681 14887 6715
rect 14829 6675 14887 6681
rect 15286 6672 15292 6724
rect 15344 6712 15350 6724
rect 16040 6712 16068 6743
rect 16684 6724 16712 6752
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 18693 6783 18751 6789
rect 18693 6749 18705 6783
rect 18739 6780 18751 6783
rect 19242 6780 19248 6792
rect 18739 6752 19248 6780
rect 18739 6749 18751 6752
rect 18693 6743 18751 6749
rect 19242 6740 19248 6752
rect 19300 6780 19306 6792
rect 22186 6780 22192 6792
rect 19300 6752 22192 6780
rect 19300 6740 19306 6752
rect 22186 6740 22192 6752
rect 22244 6780 22250 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 22244 6752 22477 6780
rect 22244 6740 22250 6752
rect 22465 6749 22477 6752
rect 22511 6749 22523 6783
rect 22465 6743 22523 6749
rect 22741 6783 22799 6789
rect 22741 6749 22753 6783
rect 22787 6749 22799 6783
rect 26786 6780 26792 6792
rect 26747 6752 26792 6780
rect 22741 6743 22799 6749
rect 16666 6712 16672 6724
rect 15344 6684 16068 6712
rect 16579 6684 16672 6712
rect 15344 6672 15350 6684
rect 16666 6672 16672 6684
rect 16724 6672 16730 6724
rect 16853 6715 16911 6721
rect 16853 6681 16865 6715
rect 16899 6681 16911 6715
rect 18046 6712 18052 6724
rect 17959 6684 18052 6712
rect 16853 6675 16911 6681
rect 12618 6644 12624 6656
rect 9048 6616 12480 6644
rect 12579 6616 12624 6644
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 15102 6604 15108 6656
rect 15160 6644 15166 6656
rect 16485 6647 16543 6653
rect 16485 6644 16497 6647
rect 15160 6616 16497 6644
rect 15160 6604 15166 6616
rect 16485 6613 16497 6616
rect 16531 6613 16543 6647
rect 16868 6644 16896 6675
rect 18046 6672 18052 6684
rect 18104 6712 18110 6724
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 18104 6684 19625 6712
rect 18104 6672 18110 6684
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 22756 6712 22784 6743
rect 26786 6740 26792 6752
rect 26844 6740 26850 6792
rect 27893 6783 27951 6789
rect 27893 6749 27905 6783
rect 27939 6780 27951 6783
rect 28810 6780 28816 6792
rect 27939 6752 28816 6780
rect 27939 6749 27951 6752
rect 27893 6743 27951 6749
rect 28810 6740 28816 6752
rect 28868 6740 28874 6792
rect 30190 6780 30196 6792
rect 30151 6752 30196 6780
rect 30190 6740 30196 6752
rect 30248 6740 30254 6792
rect 32766 6740 32772 6792
rect 32824 6780 32830 6792
rect 36924 6789 36952 6820
rect 35161 6783 35219 6789
rect 35161 6780 35173 6783
rect 32824 6752 35173 6780
rect 32824 6740 32830 6752
rect 35161 6749 35173 6752
rect 35207 6749 35219 6783
rect 35161 6743 35219 6749
rect 36909 6783 36967 6789
rect 36909 6749 36921 6783
rect 36955 6749 36967 6783
rect 37921 6783 37979 6789
rect 37921 6780 37933 6783
rect 36909 6743 36967 6749
rect 37292 6752 37933 6780
rect 28077 6715 28135 6721
rect 28077 6712 28089 6715
rect 22756 6684 28089 6712
rect 19613 6675 19671 6681
rect 28077 6681 28089 6684
rect 28123 6712 28135 6715
rect 29270 6712 29276 6724
rect 28123 6684 29276 6712
rect 28123 6681 28135 6684
rect 28077 6675 28135 6681
rect 29270 6672 29276 6684
rect 29328 6672 29334 6724
rect 30460 6715 30518 6721
rect 30460 6681 30472 6715
rect 30506 6712 30518 6715
rect 30742 6712 30748 6724
rect 30506 6684 30748 6712
rect 30506 6681 30518 6684
rect 30460 6675 30518 6681
rect 30742 6672 30748 6684
rect 30800 6672 30806 6724
rect 35176 6712 35204 6743
rect 37292 6724 37320 6752
rect 37921 6749 37933 6752
rect 37967 6749 37979 6783
rect 37921 6743 37979 6749
rect 38010 6740 38016 6792
rect 38068 6780 38074 6792
rect 38177 6783 38235 6789
rect 38177 6780 38189 6783
rect 38068 6752 38189 6780
rect 38068 6740 38074 6752
rect 38177 6749 38189 6752
rect 38223 6749 38235 6783
rect 38177 6743 38235 6749
rect 37274 6712 37280 6724
rect 35176 6684 37280 6712
rect 37274 6672 37280 6684
rect 37332 6672 37338 6724
rect 17034 6644 17040 6656
rect 16868 6616 17040 6644
rect 16485 6607 16543 6613
rect 17034 6604 17040 6616
rect 17092 6644 17098 6656
rect 17862 6644 17868 6656
rect 17092 6616 17868 6644
rect 17092 6604 17098 6616
rect 17862 6604 17868 6616
rect 17920 6644 17926 6656
rect 18509 6647 18567 6653
rect 18509 6644 18521 6647
rect 17920 6616 18521 6644
rect 17920 6604 17926 6616
rect 18509 6613 18521 6616
rect 18555 6613 18567 6647
rect 18509 6607 18567 6613
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 20438 6644 20444 6656
rect 18748 6616 20444 6644
rect 18748 6604 18754 6616
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 25501 6647 25559 6653
rect 25501 6613 25513 6647
rect 25547 6644 25559 6647
rect 25590 6644 25596 6656
rect 25547 6616 25596 6644
rect 25547 6613 25559 6616
rect 25501 6607 25559 6613
rect 25590 6604 25596 6616
rect 25648 6604 25654 6656
rect 27430 6604 27436 6656
rect 27488 6644 27494 6656
rect 27709 6647 27767 6653
rect 27709 6644 27721 6647
rect 27488 6616 27721 6644
rect 27488 6604 27494 6616
rect 27709 6613 27721 6616
rect 27755 6613 27767 6647
rect 27709 6607 27767 6613
rect 29178 6604 29184 6656
rect 29236 6644 29242 6656
rect 30558 6644 30564 6656
rect 29236 6616 30564 6644
rect 29236 6604 29242 6616
rect 30558 6604 30564 6616
rect 30616 6604 30622 6656
rect 31478 6604 31484 6656
rect 31536 6644 31542 6656
rect 31573 6647 31631 6653
rect 31573 6644 31585 6647
rect 31536 6616 31585 6644
rect 31536 6604 31542 6616
rect 31573 6613 31585 6616
rect 31619 6613 31631 6647
rect 31573 6607 31631 6613
rect 37182 6604 37188 6656
rect 37240 6644 37246 6656
rect 39301 6647 39359 6653
rect 39301 6644 39313 6647
rect 37240 6616 39313 6644
rect 37240 6604 37246 6616
rect 39301 6613 39313 6616
rect 39347 6613 39359 6647
rect 39301 6607 39359 6613
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 3513 6443 3571 6449
rect 3513 6409 3525 6443
rect 3559 6440 3571 6443
rect 4433 6443 4491 6449
rect 4433 6440 4445 6443
rect 3559 6412 4445 6440
rect 3559 6409 3571 6412
rect 3513 6403 3571 6409
rect 4433 6409 4445 6412
rect 4479 6440 4491 6443
rect 4890 6440 4896 6452
rect 4479 6412 4896 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4890 6400 4896 6412
rect 4948 6440 4954 6452
rect 8018 6440 8024 6452
rect 4948 6412 8024 6440
rect 4948 6400 4954 6412
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6409 8355 6443
rect 8297 6403 8355 6409
rect 1857 6375 1915 6381
rect 1857 6341 1869 6375
rect 1903 6372 1915 6375
rect 4062 6372 4068 6384
rect 1903 6344 4068 6372
rect 1903 6341 1915 6344
rect 1857 6335 1915 6341
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 7282 6372 7288 6384
rect 5460 6344 7288 6372
rect 2406 6304 2412 6316
rect 2367 6276 2412 6304
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6304 2559 6307
rect 2547 6276 2774 6304
rect 2547 6273 2559 6276
rect 2501 6267 2559 6273
rect 2746 6168 2774 6276
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5460 6313 5488 6344
rect 7282 6332 7288 6344
rect 7340 6332 7346 6384
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 7892 6344 8156 6372
rect 7892 6332 7898 6344
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 5224 6276 5273 6304
rect 5224 6264 5230 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 5718 6304 5724 6316
rect 5675 6276 5724 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 5994 6304 6000 6316
rect 5859 6276 6000 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 3602 6236 3608 6248
rect 3563 6208 3608 6236
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3789 6239 3847 6245
rect 3789 6205 3801 6239
rect 3835 6236 3847 6239
rect 3878 6236 3884 6248
rect 3835 6208 3884 6236
rect 3835 6205 3847 6208
rect 3789 6199 3847 6205
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 5534 6236 5540 6248
rect 5495 6208 5540 6236
rect 5534 6196 5540 6208
rect 5592 6196 5598 6248
rect 6380 6236 6408 6267
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6549 6307 6607 6313
rect 6549 6304 6561 6307
rect 6512 6276 6561 6304
rect 6512 6264 6518 6276
rect 6549 6273 6561 6276
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 8018 6304 8024 6316
rect 7515 6276 8024 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8128 6313 8156 6344
rect 8312 6316 8340 6403
rect 15194 6400 15200 6452
rect 15252 6400 15258 6452
rect 15562 6400 15568 6452
rect 15620 6440 15626 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 15620 6412 16681 6440
rect 15620 6400 15626 6412
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 16669 6403 16727 6409
rect 19797 6443 19855 6449
rect 19797 6409 19809 6443
rect 19843 6440 19855 6443
rect 19978 6440 19984 6452
rect 19843 6412 19984 6440
rect 19843 6409 19855 6412
rect 19797 6403 19855 6409
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 24673 6443 24731 6449
rect 24673 6409 24685 6443
rect 24719 6440 24731 6443
rect 24946 6440 24952 6452
rect 24719 6412 24952 6440
rect 24719 6409 24731 6412
rect 24673 6403 24731 6409
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 28445 6443 28503 6449
rect 28445 6409 28457 6443
rect 28491 6440 28503 6443
rect 28810 6440 28816 6452
rect 28491 6412 28816 6440
rect 28491 6409 28503 6412
rect 28445 6403 28503 6409
rect 28810 6400 28816 6412
rect 28868 6400 28874 6452
rect 30742 6440 30748 6452
rect 30703 6412 30748 6440
rect 30742 6400 30748 6412
rect 30800 6400 30806 6452
rect 33778 6440 33784 6452
rect 33739 6412 33784 6440
rect 33778 6400 33784 6412
rect 33836 6400 33842 6452
rect 35894 6400 35900 6452
rect 35952 6400 35958 6452
rect 39114 6440 39120 6452
rect 39075 6412 39120 6440
rect 39114 6400 39120 6412
rect 39172 6400 39178 6452
rect 12802 6332 12808 6384
rect 12860 6381 12866 6384
rect 12860 6372 12872 6381
rect 15212 6372 15240 6400
rect 17037 6375 17095 6381
rect 12860 6344 12905 6372
rect 15212 6344 15332 6372
rect 12860 6335 12872 6344
rect 12860 6332 12866 6335
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8754 6304 8760 6316
rect 8715 6276 8760 6304
rect 8754 6264 8760 6276
rect 8812 6264 8818 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 8904 6276 13032 6304
rect 8904 6264 8910 6276
rect 7558 6236 7564 6248
rect 5644 6208 7564 6236
rect 5644 6180 5672 6208
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 8036 6236 8064 6264
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 8036 6208 9413 6236
rect 9401 6205 9413 6208
rect 9447 6205 9459 6239
rect 13004 6236 13032 6276
rect 13078 6264 13084 6316
rect 13136 6304 13142 6316
rect 14458 6304 14464 6316
rect 13136 6276 14464 6304
rect 13136 6264 13142 6276
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 15194 6304 15200 6316
rect 15155 6276 15200 6304
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15304 6304 15332 6344
rect 17037 6341 17049 6375
rect 17083 6372 17095 6375
rect 17862 6372 17868 6384
rect 17083 6344 17868 6372
rect 17083 6341 17095 6344
rect 17037 6335 17095 6341
rect 17862 6332 17868 6344
rect 17920 6332 17926 6384
rect 20714 6372 20720 6384
rect 18616 6344 20720 6372
rect 15360 6307 15418 6313
rect 15360 6304 15372 6307
rect 15304 6276 15372 6304
rect 15360 6273 15372 6276
rect 15406 6273 15418 6307
rect 15360 6267 15418 6273
rect 15476 6307 15534 6313
rect 15476 6273 15488 6307
rect 15522 6273 15534 6307
rect 15476 6267 15534 6273
rect 15565 6307 15623 6313
rect 15565 6273 15577 6307
rect 15611 6304 15623 6307
rect 15654 6304 15660 6316
rect 15611 6276 15660 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 13004 6208 13124 6236
rect 9401 6199 9459 6205
rect 3145 6171 3203 6177
rect 3145 6168 3157 6171
rect 2746 6140 3157 6168
rect 3145 6137 3157 6140
rect 3191 6137 3203 6171
rect 3145 6131 3203 6137
rect 3510 6128 3516 6180
rect 3568 6168 3574 6180
rect 3568 6140 5580 6168
rect 3568 6128 3574 6140
rect 2685 6103 2743 6109
rect 2685 6069 2697 6103
rect 2731 6100 2743 6103
rect 2866 6100 2872 6112
rect 2731 6072 2872 6100
rect 2731 6069 2743 6072
rect 2685 6063 2743 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 5074 6100 5080 6112
rect 5035 6072 5080 6100
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5552 6100 5580 6140
rect 5626 6128 5632 6180
rect 5684 6128 5690 6180
rect 7653 6171 7711 6177
rect 6196 6140 6960 6168
rect 6196 6100 6224 6140
rect 6362 6100 6368 6112
rect 5552 6072 6224 6100
rect 6323 6072 6368 6100
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6932 6100 6960 6140
rect 7653 6137 7665 6171
rect 7699 6168 7711 6171
rect 8386 6168 8392 6180
rect 7699 6140 8392 6168
rect 7699 6137 7711 6140
rect 7653 6131 7711 6137
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 13096 6168 13124 6208
rect 14918 6196 14924 6248
rect 14976 6236 14982 6248
rect 15488 6236 15516 6267
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6304 16911 6307
rect 18616 6304 18644 6344
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 21266 6332 21272 6384
rect 21324 6372 21330 6384
rect 22005 6375 22063 6381
rect 22005 6372 22017 6375
rect 21324 6344 22017 6372
rect 21324 6332 21330 6344
rect 22005 6341 22017 6344
rect 22051 6341 22063 6375
rect 22186 6372 22192 6384
rect 22147 6344 22192 6372
rect 22005 6335 22063 6341
rect 22186 6332 22192 6344
rect 22244 6332 22250 6384
rect 24854 6372 24860 6384
rect 23308 6344 24860 6372
rect 20070 6304 20076 6316
rect 16899 6276 18644 6304
rect 20031 6276 20076 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17052 6248 17080 6276
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6273 20315 6307
rect 20438 6304 20444 6316
rect 20399 6276 20444 6304
rect 20257 6267 20315 6273
rect 14976 6208 15516 6236
rect 14976 6196 14982 6208
rect 17034 6196 17040 6248
rect 17092 6196 17098 6248
rect 19058 6236 19064 6248
rect 19019 6208 19064 6236
rect 19058 6196 19064 6208
rect 19116 6196 19122 6248
rect 19334 6236 19340 6248
rect 19247 6208 19340 6236
rect 19334 6196 19340 6208
rect 19392 6236 19398 6248
rect 20180 6236 20208 6267
rect 19392 6208 20208 6236
rect 20272 6236 20300 6267
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 23308 6313 23336 6344
rect 24854 6332 24860 6344
rect 24912 6372 24918 6384
rect 25590 6372 25596 6384
rect 24912 6344 25596 6372
rect 24912 6332 24918 6344
rect 25590 6332 25596 6344
rect 25648 6332 25654 6384
rect 29270 6372 29276 6384
rect 29231 6344 29276 6372
rect 29270 6332 29276 6344
rect 29328 6332 29334 6384
rect 29457 6375 29515 6381
rect 29457 6341 29469 6375
rect 29503 6372 29515 6375
rect 31478 6372 31484 6384
rect 29503 6344 31484 6372
rect 29503 6341 29515 6344
rect 29457 6335 29515 6341
rect 31478 6332 31484 6344
rect 31536 6332 31542 6384
rect 23566 6313 23572 6316
rect 23293 6307 23351 6313
rect 23293 6273 23305 6307
rect 23339 6273 23351 6307
rect 23560 6304 23572 6313
rect 23527 6276 23572 6304
rect 23293 6267 23351 6273
rect 23560 6267 23572 6276
rect 23566 6264 23572 6267
rect 23624 6264 23630 6316
rect 27062 6304 27068 6316
rect 27023 6276 27068 6304
rect 27062 6264 27068 6276
rect 27120 6264 27126 6316
rect 27154 6264 27160 6316
rect 27212 6304 27218 6316
rect 27321 6307 27379 6313
rect 27321 6304 27333 6307
rect 27212 6276 27333 6304
rect 27212 6264 27218 6276
rect 27321 6273 27333 6276
rect 27367 6273 27379 6307
rect 27321 6267 27379 6273
rect 30006 6264 30012 6316
rect 30064 6304 30070 6316
rect 30101 6307 30159 6313
rect 30101 6304 30113 6307
rect 30064 6276 30113 6304
rect 30064 6264 30070 6276
rect 30101 6273 30113 6276
rect 30147 6273 30159 6307
rect 30101 6267 30159 6273
rect 30285 6307 30343 6313
rect 30285 6273 30297 6307
rect 30331 6273 30343 6307
rect 30285 6267 30343 6273
rect 30377 6307 30435 6313
rect 30377 6273 30389 6307
rect 30423 6273 30435 6307
rect 30377 6267 30435 6273
rect 30469 6307 30527 6313
rect 30469 6273 30481 6307
rect 30515 6304 30527 6307
rect 30558 6304 30564 6316
rect 30515 6276 30564 6304
rect 30515 6273 30527 6276
rect 30469 6267 30527 6273
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 20272 6208 21833 6236
rect 19392 6196 19398 6208
rect 18966 6168 18972 6180
rect 8864 6140 12204 6168
rect 13096 6140 18972 6168
rect 8864 6100 8892 6140
rect 6932 6072 8892 6100
rect 8941 6103 8999 6109
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 9306 6100 9312 6112
rect 8987 6072 9312 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 10318 6100 10324 6112
rect 10183 6072 10324 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10597 6103 10655 6109
rect 10597 6100 10609 6103
rect 10560 6072 10609 6100
rect 10560 6060 10566 6072
rect 10597 6069 10609 6072
rect 10643 6069 10655 6103
rect 10597 6063 10655 6069
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11664 6072 11713 6100
rect 11664 6060 11670 6072
rect 11701 6069 11713 6072
rect 11747 6100 11759 6103
rect 11974 6100 11980 6112
rect 11747 6072 11980 6100
rect 11747 6069 11759 6072
rect 11701 6063 11759 6069
rect 11974 6060 11980 6072
rect 12032 6060 12038 6112
rect 12176 6100 12204 6140
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 20180 6168 20208 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 25593 6239 25651 6245
rect 25593 6205 25605 6239
rect 25639 6205 25651 6239
rect 25593 6199 25651 6205
rect 25869 6239 25927 6245
rect 25869 6205 25881 6239
rect 25915 6236 25927 6239
rect 26970 6236 26976 6248
rect 25915 6208 26976 6236
rect 25915 6205 25927 6208
rect 25869 6199 25927 6205
rect 25608 6168 25636 6199
rect 26970 6196 26976 6208
rect 27028 6196 27034 6248
rect 29641 6239 29699 6245
rect 29641 6205 29653 6239
rect 29687 6236 29699 6239
rect 30300 6236 30328 6267
rect 29687 6208 30328 6236
rect 30392 6236 30420 6267
rect 30558 6264 30564 6276
rect 30616 6304 30622 6316
rect 31205 6307 31263 6313
rect 31205 6304 31217 6307
rect 30616 6276 31217 6304
rect 30616 6264 30622 6276
rect 31205 6273 31217 6276
rect 31251 6273 31263 6307
rect 33796 6304 33824 6400
rect 35912 6372 35940 6400
rect 34716 6344 36032 6372
rect 34716 6313 34744 6344
rect 34609 6307 34667 6313
rect 34609 6304 34621 6307
rect 33796 6276 34621 6304
rect 31205 6267 31263 6273
rect 34609 6273 34621 6276
rect 34655 6273 34667 6307
rect 34609 6267 34667 6273
rect 34701 6307 34759 6313
rect 34701 6273 34713 6307
rect 34747 6273 34759 6307
rect 34701 6267 34759 6273
rect 34790 6264 34796 6316
rect 34848 6304 34854 6316
rect 34977 6307 35035 6313
rect 34848 6276 34893 6304
rect 34848 6264 34854 6276
rect 34977 6273 34989 6307
rect 35023 6304 35035 6307
rect 35618 6304 35624 6316
rect 35023 6276 35624 6304
rect 35023 6273 35035 6276
rect 34977 6267 35035 6273
rect 35618 6264 35624 6276
rect 35676 6304 35682 6316
rect 35713 6307 35771 6313
rect 35713 6304 35725 6307
rect 35676 6276 35725 6304
rect 35676 6264 35682 6276
rect 35713 6273 35725 6276
rect 35759 6273 35771 6307
rect 35894 6304 35900 6316
rect 35855 6276 35900 6304
rect 35713 6267 35771 6273
rect 35894 6264 35900 6276
rect 35952 6264 35958 6316
rect 36004 6313 36032 6344
rect 37826 6332 37832 6384
rect 37884 6372 37890 6384
rect 37982 6375 38040 6381
rect 37982 6372 37994 6375
rect 37884 6344 37994 6372
rect 37884 6332 37890 6344
rect 37982 6341 37994 6344
rect 38028 6341 38040 6375
rect 37982 6335 38040 6341
rect 35989 6307 36047 6313
rect 35989 6273 36001 6307
rect 36035 6273 36047 6307
rect 35989 6267 36047 6273
rect 36078 6264 36084 6316
rect 36136 6304 36142 6316
rect 36136 6276 36181 6304
rect 36136 6264 36142 6276
rect 37274 6264 37280 6316
rect 37332 6304 37338 6316
rect 37737 6307 37795 6313
rect 37737 6304 37749 6307
rect 37332 6276 37749 6304
rect 37332 6264 37338 6276
rect 37737 6273 37749 6276
rect 37783 6273 37795 6307
rect 37737 6267 37795 6273
rect 30392 6208 30512 6236
rect 29687 6205 29699 6208
rect 29641 6199 29699 6205
rect 30484 6180 30512 6208
rect 20180 6140 22094 6168
rect 14642 6100 14648 6112
rect 12176 6072 14648 6100
rect 14642 6060 14648 6072
rect 14700 6100 14706 6112
rect 15654 6100 15660 6112
rect 14700 6072 15660 6100
rect 14700 6060 14706 6072
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 15746 6060 15752 6112
rect 15804 6100 15810 6112
rect 15841 6103 15899 6109
rect 15841 6100 15853 6103
rect 15804 6072 15853 6100
rect 15804 6060 15810 6072
rect 15841 6069 15853 6072
rect 15887 6069 15899 6103
rect 15841 6063 15899 6069
rect 20070 6060 20076 6112
rect 20128 6100 20134 6112
rect 20901 6103 20959 6109
rect 20901 6100 20913 6103
rect 20128 6072 20913 6100
rect 20128 6060 20134 6072
rect 20901 6069 20913 6072
rect 20947 6069 20959 6103
rect 22066 6100 22094 6140
rect 24228 6140 25636 6168
rect 24228 6100 24256 6140
rect 30466 6128 30472 6180
rect 30524 6128 30530 6180
rect 58158 6168 58164 6180
rect 58119 6140 58164 6168
rect 58158 6128 58164 6140
rect 58216 6128 58222 6180
rect 34330 6100 34336 6112
rect 22066 6072 24256 6100
rect 34291 6072 34336 6100
rect 20901 6063 20959 6069
rect 34330 6060 34336 6072
rect 34388 6060 34394 6112
rect 36357 6103 36415 6109
rect 36357 6069 36369 6103
rect 36403 6100 36415 6103
rect 36998 6100 37004 6112
rect 36403 6072 37004 6100
rect 36403 6069 36415 6072
rect 36357 6063 36415 6069
rect 36998 6060 37004 6072
rect 37056 6060 37062 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 2130 5896 2136 5908
rect 1872 5868 2136 5896
rect 1872 5769 1900 5868
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 5718 5896 5724 5908
rect 5679 5868 5724 5896
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 6730 5896 6736 5908
rect 6691 5868 6736 5896
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 7616 5868 9352 5896
rect 7616 5856 7622 5868
rect 3237 5831 3295 5837
rect 3237 5797 3249 5831
rect 3283 5797 3295 5831
rect 3237 5791 3295 5797
rect 6825 5831 6883 5837
rect 6825 5797 6837 5831
rect 6871 5828 6883 5831
rect 8018 5828 8024 5840
rect 6871 5800 8024 5828
rect 6871 5797 6883 5800
rect 6825 5791 6883 5797
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5729 1915 5763
rect 3252 5760 3280 5791
rect 8018 5788 8024 5800
rect 8076 5828 8082 5840
rect 8205 5831 8263 5837
rect 8205 5828 8217 5831
rect 8076 5800 8217 5828
rect 8076 5788 8082 5800
rect 8205 5797 8217 5800
rect 8251 5797 8263 5831
rect 9324 5828 9352 5868
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 11882 5896 11888 5908
rect 9824 5868 11888 5896
rect 9824 5856 9830 5868
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 12406 5868 12817 5896
rect 10137 5831 10195 5837
rect 10137 5828 10149 5831
rect 9324 5800 10149 5828
rect 8205 5791 8263 5797
rect 10137 5797 10149 5800
rect 10183 5828 10195 5831
rect 10410 5828 10416 5840
rect 10183 5800 10416 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 10505 5831 10563 5837
rect 10505 5797 10517 5831
rect 10551 5828 10563 5831
rect 11790 5828 11796 5840
rect 10551 5800 11796 5828
rect 10551 5797 10563 5800
rect 10505 5791 10563 5797
rect 11790 5788 11796 5800
rect 11848 5828 11854 5840
rect 12406 5828 12434 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 13357 5899 13415 5905
rect 13357 5865 13369 5899
rect 13403 5896 13415 5899
rect 17034 5896 17040 5908
rect 13403 5868 16896 5896
rect 16995 5868 17040 5896
rect 13403 5865 13415 5868
rect 13357 5859 13415 5865
rect 11848 5800 12434 5828
rect 11848 5788 11854 5800
rect 3602 5760 3608 5772
rect 3252 5732 3608 5760
rect 1857 5723 1915 5729
rect 3602 5720 3608 5732
rect 3660 5760 3666 5772
rect 5445 5763 5503 5769
rect 5445 5760 5457 5763
rect 3660 5732 5457 5760
rect 3660 5720 3666 5732
rect 5445 5729 5457 5732
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 10229 5763 10287 5769
rect 10229 5760 10241 5763
rect 6512 5732 10241 5760
rect 6512 5720 6518 5732
rect 10229 5729 10241 5732
rect 10275 5760 10287 5763
rect 10594 5760 10600 5772
rect 10275 5732 10600 5760
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 12820 5760 12848 5859
rect 14918 5788 14924 5840
rect 14976 5788 14982 5840
rect 16868 5828 16896 5868
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 19426 5896 19432 5908
rect 17797 5868 19432 5896
rect 17797 5828 17825 5868
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 20257 5899 20315 5905
rect 20257 5865 20269 5899
rect 20303 5896 20315 5899
rect 20438 5896 20444 5908
rect 20303 5868 20444 5896
rect 20303 5865 20315 5868
rect 20257 5859 20315 5865
rect 20438 5856 20444 5868
rect 20496 5856 20502 5908
rect 24397 5899 24455 5905
rect 24397 5865 24409 5899
rect 24443 5896 24455 5899
rect 24762 5896 24768 5908
rect 24443 5868 24768 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 24762 5856 24768 5868
rect 24820 5856 24826 5908
rect 26973 5899 27031 5905
rect 26973 5865 26985 5899
rect 27019 5896 27031 5899
rect 27154 5896 27160 5908
rect 27019 5868 27160 5896
rect 27019 5865 27031 5868
rect 26973 5859 27031 5865
rect 27154 5856 27160 5868
rect 27212 5856 27218 5908
rect 30653 5899 30711 5905
rect 30653 5865 30665 5899
rect 30699 5896 30711 5899
rect 30834 5896 30840 5908
rect 30699 5868 30840 5896
rect 30699 5865 30711 5868
rect 30653 5859 30711 5865
rect 16868 5800 17825 5828
rect 17865 5831 17923 5837
rect 17865 5797 17877 5831
rect 17911 5828 17923 5831
rect 18506 5828 18512 5840
rect 17911 5800 18512 5828
rect 17911 5797 17923 5800
rect 17865 5791 17923 5797
rect 18506 5788 18512 5800
rect 18564 5828 18570 5840
rect 20898 5828 20904 5840
rect 18564 5800 20904 5828
rect 18564 5788 18570 5800
rect 20898 5788 20904 5800
rect 20956 5788 20962 5840
rect 12820 5732 13584 5760
rect 4522 5652 4528 5704
rect 4580 5692 4586 5704
rect 4890 5692 4896 5704
rect 4580 5664 4896 5692
rect 4580 5652 4586 5664
rect 4890 5652 4896 5664
rect 4948 5652 4954 5704
rect 5534 5692 5540 5704
rect 5495 5664 5540 5692
rect 5534 5652 5540 5664
rect 5592 5692 5598 5704
rect 6822 5692 6828 5704
rect 5592 5664 6828 5692
rect 5592 5652 5598 5664
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 6972 5664 7017 5692
rect 6972 5652 6978 5664
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7156 5664 7665 5692
rect 7156 5652 7162 5664
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 8386 5692 8392 5704
rect 8347 5664 8392 5692
rect 7653 5655 7711 5661
rect 8386 5652 8392 5664
rect 8444 5692 8450 5704
rect 9122 5692 9128 5704
rect 8444 5664 9128 5692
rect 8444 5652 8450 5664
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5692 9459 5695
rect 9674 5692 9680 5704
rect 9447 5664 9680 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 10042 5701 10048 5704
rect 10008 5695 10048 5701
rect 10008 5661 10020 5695
rect 10008 5655 10048 5661
rect 10042 5652 10048 5655
rect 10100 5652 10106 5704
rect 11330 5652 11336 5704
rect 11388 5692 11394 5704
rect 11425 5695 11483 5701
rect 11425 5692 11437 5695
rect 11388 5664 11437 5692
rect 11388 5652 11394 5664
rect 11425 5661 11437 5664
rect 11471 5661 11483 5695
rect 11425 5655 11483 5661
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5661 12127 5695
rect 13354 5692 13360 5704
rect 13315 5664 13360 5692
rect 12069 5655 12127 5661
rect 2124 5627 2182 5633
rect 2124 5593 2136 5627
rect 2170 5624 2182 5627
rect 2958 5624 2964 5636
rect 2170 5596 2964 5624
rect 2170 5593 2182 5596
rect 2124 5587 2182 5593
rect 2958 5584 2964 5596
rect 3016 5584 3022 5636
rect 4065 5627 4123 5633
rect 4065 5593 4077 5627
rect 4111 5624 4123 5627
rect 5442 5624 5448 5636
rect 4111 5596 5448 5624
rect 4111 5593 4123 5596
rect 4065 5587 4123 5593
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 6641 5627 6699 5633
rect 6641 5593 6653 5627
rect 6687 5624 6699 5627
rect 7374 5624 7380 5636
rect 6687 5596 7380 5624
rect 6687 5593 6699 5596
rect 6641 5587 6699 5593
rect 7374 5584 7380 5596
rect 7432 5624 7438 5636
rect 9858 5624 9864 5636
rect 7432 5596 9864 5624
rect 7432 5584 7438 5596
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 10226 5584 10232 5636
rect 10284 5624 10290 5636
rect 12084 5624 12112 5655
rect 13354 5652 13360 5664
rect 13412 5652 13418 5704
rect 13556 5701 13584 5732
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5661 13599 5695
rect 14826 5692 14832 5704
rect 14787 5664 14832 5692
rect 13541 5655 13599 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 14933 5701 14961 5788
rect 18693 5763 18751 5769
rect 18432 5732 18644 5760
rect 14918 5695 14976 5701
rect 14918 5661 14930 5695
rect 14964 5661 14976 5695
rect 14918 5655 14976 5661
rect 15013 5692 15071 5698
rect 15102 5692 15108 5704
rect 15013 5658 15025 5692
rect 15059 5664 15108 5692
rect 15059 5658 15071 5664
rect 15013 5652 15071 5658
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15197 5695 15255 5701
rect 15197 5661 15209 5695
rect 15243 5692 15255 5695
rect 15286 5692 15292 5704
rect 15243 5664 15292 5692
rect 15243 5661 15255 5664
rect 15197 5655 15255 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 10284 5596 12112 5624
rect 15672 5624 15700 5655
rect 15746 5652 15752 5704
rect 15804 5692 15810 5704
rect 15913 5695 15971 5701
rect 15913 5692 15925 5695
rect 15804 5664 15925 5692
rect 15804 5652 15810 5664
rect 15913 5661 15925 5664
rect 15959 5661 15971 5695
rect 18432 5692 18460 5732
rect 15913 5655 15971 5661
rect 16040 5664 18460 5692
rect 18616 5692 18644 5732
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 19334 5760 19340 5772
rect 18739 5732 19340 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 19334 5720 19340 5732
rect 19392 5720 19398 5772
rect 26970 5720 26976 5772
rect 27028 5760 27034 5772
rect 27028 5732 27384 5760
rect 27028 5720 27034 5732
rect 20622 5692 20628 5704
rect 18616 5664 20628 5692
rect 16040 5624 16068 5664
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 23474 5652 23480 5704
rect 23532 5692 23538 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 23532 5664 24593 5692
rect 23532 5652 23538 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 24765 5695 24823 5701
rect 24765 5661 24777 5695
rect 24811 5692 24823 5695
rect 25866 5692 25872 5704
rect 24811 5664 25872 5692
rect 24811 5661 24823 5664
rect 24765 5655 24823 5661
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 26234 5652 26240 5704
rect 26292 5692 26298 5704
rect 26513 5695 26571 5701
rect 26513 5692 26525 5695
rect 26292 5664 26525 5692
rect 26292 5652 26298 5664
rect 26513 5661 26525 5664
rect 26559 5692 26571 5695
rect 27246 5692 27252 5704
rect 26559 5664 27252 5692
rect 26559 5661 26571 5664
rect 26513 5655 26571 5661
rect 27246 5652 27252 5664
rect 27304 5652 27310 5704
rect 27356 5701 27384 5732
rect 27341 5695 27399 5701
rect 27341 5661 27353 5695
rect 27387 5661 27399 5695
rect 27341 5655 27399 5661
rect 27430 5652 27436 5704
rect 27488 5692 27494 5704
rect 27617 5695 27675 5701
rect 27488 5664 27533 5692
rect 27488 5652 27494 5664
rect 27617 5661 27629 5695
rect 27663 5661 27675 5695
rect 27617 5655 27675 5661
rect 15672 5596 16068 5624
rect 10284 5584 10290 5596
rect 17862 5584 17868 5636
rect 17920 5624 17926 5636
rect 18325 5627 18383 5633
rect 18325 5624 18337 5627
rect 17920 5596 18337 5624
rect 17920 5584 17926 5596
rect 18325 5593 18337 5596
rect 18371 5593 18383 5627
rect 18506 5624 18512 5636
rect 18467 5596 18512 5624
rect 18325 5587 18383 5593
rect 4617 5559 4675 5565
rect 4617 5525 4629 5559
rect 4663 5556 4675 5559
rect 4890 5556 4896 5568
rect 4663 5528 4896 5556
rect 4663 5525 4675 5528
rect 4617 5519 4675 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 5077 5559 5135 5565
rect 5077 5525 5089 5559
rect 5123 5556 5135 5559
rect 6270 5556 6276 5568
rect 5123 5528 6276 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 6822 5556 6828 5568
rect 6512 5528 6828 5556
rect 6512 5516 6518 5528
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7469 5559 7527 5565
rect 7469 5556 7481 5559
rect 7064 5528 7481 5556
rect 7064 5516 7070 5528
rect 7469 5525 7481 5528
rect 7515 5525 7527 5559
rect 14550 5556 14556 5568
rect 14511 5528 14556 5556
rect 7469 5519 7527 5525
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 18340 5556 18368 5587
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 19337 5627 19395 5633
rect 19337 5593 19349 5627
rect 19383 5593 19395 5627
rect 19337 5587 19395 5593
rect 19521 5627 19579 5633
rect 19521 5593 19533 5627
rect 19567 5624 19579 5627
rect 21266 5624 21272 5636
rect 19567 5596 21272 5624
rect 19567 5593 19579 5596
rect 19521 5587 19579 5593
rect 19352 5556 19380 5587
rect 21266 5584 21272 5596
rect 21324 5584 21330 5636
rect 27154 5584 27160 5636
rect 27212 5624 27218 5636
rect 27632 5624 27660 5655
rect 29270 5652 29276 5704
rect 29328 5692 29334 5704
rect 29825 5695 29883 5701
rect 29825 5692 29837 5695
rect 29328 5664 29837 5692
rect 29328 5652 29334 5664
rect 29825 5661 29837 5664
rect 29871 5661 29883 5695
rect 29825 5655 29883 5661
rect 30009 5695 30067 5701
rect 30009 5661 30021 5695
rect 30055 5692 30067 5695
rect 30668 5692 30696 5859
rect 30834 5856 30840 5868
rect 30892 5856 30898 5908
rect 34701 5899 34759 5905
rect 34701 5865 34713 5899
rect 34747 5896 34759 5899
rect 34790 5896 34796 5908
rect 34747 5868 34796 5896
rect 34747 5865 34759 5868
rect 34701 5859 34759 5865
rect 34790 5856 34796 5868
rect 34848 5856 34854 5908
rect 35894 5856 35900 5908
rect 35952 5896 35958 5908
rect 35989 5899 36047 5905
rect 35989 5896 36001 5899
rect 35952 5868 36001 5896
rect 35952 5856 35958 5868
rect 35989 5865 36001 5868
rect 36035 5865 36047 5899
rect 35989 5859 36047 5865
rect 37369 5899 37427 5905
rect 37369 5865 37381 5899
rect 37415 5896 37427 5899
rect 37458 5896 37464 5908
rect 37415 5868 37464 5896
rect 37415 5865 37427 5868
rect 37369 5859 37427 5865
rect 37458 5856 37464 5868
rect 37516 5856 37522 5908
rect 32033 5763 32091 5769
rect 32033 5729 32045 5763
rect 32079 5760 32091 5763
rect 32766 5760 32772 5772
rect 32079 5732 32772 5760
rect 32079 5729 32091 5732
rect 32033 5723 32091 5729
rect 32766 5720 32772 5732
rect 32824 5720 32830 5772
rect 30055 5664 30696 5692
rect 34885 5695 34943 5701
rect 30055 5661 30067 5664
rect 30009 5655 30067 5661
rect 34885 5661 34897 5695
rect 34931 5692 34943 5695
rect 35342 5692 35348 5704
rect 34931 5664 35348 5692
rect 34931 5661 34943 5664
rect 34885 5655 34943 5661
rect 35342 5652 35348 5664
rect 35400 5652 35406 5704
rect 35805 5695 35863 5701
rect 35805 5661 35817 5695
rect 35851 5692 35863 5695
rect 35986 5692 35992 5704
rect 35851 5664 35992 5692
rect 35851 5661 35863 5664
rect 35805 5655 35863 5661
rect 35986 5652 35992 5664
rect 36044 5652 36050 5704
rect 37182 5692 37188 5704
rect 37143 5664 37188 5692
rect 37182 5652 37188 5664
rect 37240 5652 37246 5704
rect 27212 5596 27660 5624
rect 27212 5584 27218 5596
rect 30834 5584 30840 5636
rect 30892 5624 30898 5636
rect 31766 5627 31824 5633
rect 31766 5624 31778 5627
rect 30892 5596 31778 5624
rect 30892 5584 30898 5596
rect 31766 5593 31778 5596
rect 31812 5593 31824 5627
rect 31766 5587 31824 5593
rect 35069 5627 35127 5633
rect 35069 5593 35081 5627
rect 35115 5624 35127 5627
rect 35526 5624 35532 5636
rect 35115 5596 35532 5624
rect 35115 5593 35127 5596
rect 35069 5587 35127 5593
rect 35526 5584 35532 5596
rect 35584 5624 35590 5636
rect 35621 5627 35679 5633
rect 35621 5624 35633 5627
rect 35584 5596 35633 5624
rect 35584 5584 35590 5596
rect 35621 5593 35633 5596
rect 35667 5593 35679 5627
rect 35621 5587 35679 5593
rect 37001 5627 37059 5633
rect 37001 5593 37013 5627
rect 37047 5624 37059 5627
rect 38378 5624 38384 5636
rect 37047 5596 38384 5624
rect 37047 5593 37059 5596
rect 37001 5587 37059 5593
rect 38378 5584 38384 5596
rect 38436 5584 38442 5636
rect 18340 5528 19380 5556
rect 19426 5516 19432 5568
rect 19484 5556 19490 5568
rect 19705 5559 19763 5565
rect 19705 5556 19717 5559
rect 19484 5528 19717 5556
rect 19484 5516 19490 5528
rect 19705 5525 19717 5528
rect 19751 5525 19763 5559
rect 19705 5519 19763 5525
rect 30193 5559 30251 5565
rect 30193 5525 30205 5559
rect 30239 5556 30251 5559
rect 30374 5556 30380 5568
rect 30239 5528 30380 5556
rect 30239 5525 30251 5528
rect 30193 5519 30251 5525
rect 30374 5516 30380 5528
rect 30432 5516 30438 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 6362 5312 6368 5364
rect 6420 5352 6426 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 6420 5324 6561 5352
rect 6420 5312 6426 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 8628 5324 8677 5352
rect 8628 5312 8634 5324
rect 8665 5321 8677 5324
rect 8711 5352 8723 5355
rect 14277 5355 14335 5361
rect 8711 5324 12434 5352
rect 8711 5321 8723 5324
rect 8665 5315 8723 5321
rect 1578 5244 1584 5296
rect 1636 5284 1642 5296
rect 1636 5256 2084 5284
rect 1636 5244 1642 5256
rect 2056 5225 2084 5256
rect 2130 5244 2136 5296
rect 2188 5284 2194 5296
rect 2777 5287 2835 5293
rect 2777 5284 2789 5287
rect 2188 5256 2789 5284
rect 2188 5244 2194 5256
rect 2777 5253 2789 5256
rect 2823 5253 2835 5287
rect 2777 5247 2835 5253
rect 4341 5287 4399 5293
rect 4341 5253 4353 5287
rect 4387 5284 4399 5287
rect 4614 5284 4620 5296
rect 4387 5256 4620 5284
rect 4387 5253 4399 5256
rect 4341 5247 4399 5253
rect 4614 5244 4620 5256
rect 4672 5244 4678 5296
rect 6454 5244 6460 5296
rect 6512 5284 6518 5296
rect 7101 5287 7159 5293
rect 7101 5284 7113 5287
rect 6512 5256 7113 5284
rect 6512 5244 6518 5256
rect 7101 5253 7113 5256
rect 7147 5284 7159 5287
rect 7653 5287 7711 5293
rect 7653 5284 7665 5287
rect 7147 5256 7665 5284
rect 7147 5253 7159 5256
rect 7101 5247 7159 5253
rect 7653 5253 7665 5256
rect 7699 5253 7711 5287
rect 7653 5247 7711 5253
rect 10965 5287 11023 5293
rect 10965 5253 10977 5287
rect 11011 5284 11023 5287
rect 11698 5284 11704 5296
rect 11011 5256 11704 5284
rect 11011 5253 11023 5256
rect 10965 5247 11023 5253
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 12406 5284 12434 5324
rect 14277 5321 14289 5355
rect 14323 5352 14335 5355
rect 14826 5352 14832 5364
rect 14323 5324 14832 5352
rect 14323 5321 14335 5324
rect 14277 5315 14335 5321
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 16117 5355 16175 5361
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 16666 5352 16672 5364
rect 16163 5324 16672 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 23109 5355 23167 5361
rect 19392 5324 19840 5352
rect 19392 5312 19398 5324
rect 12406 5256 13768 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5185 2007 5219
rect 1949 5179 2007 5185
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5185 2099 5219
rect 4890 5216 4896 5228
rect 4851 5188 4896 5216
rect 2041 5179 2099 5185
rect 1964 5148 1992 5179
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 5166 5176 5172 5228
rect 5224 5216 5230 5228
rect 5537 5219 5595 5225
rect 5537 5216 5549 5219
rect 5224 5188 5549 5216
rect 5224 5176 5230 5188
rect 5537 5185 5549 5188
rect 5583 5185 5595 5219
rect 5537 5179 5595 5185
rect 6270 5176 6276 5228
rect 6328 5216 6334 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6328 5188 6377 5216
rect 6328 5176 6334 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7558 5216 7564 5228
rect 6972 5188 7564 5216
rect 6972 5176 6978 5188
rect 7558 5176 7564 5188
rect 7616 5216 7622 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7616 5188 7849 5216
rect 7616 5176 7622 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 8018 5216 8024 5228
rect 7979 5188 8024 5216
rect 7837 5179 7895 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5216 8539 5219
rect 8662 5216 8668 5228
rect 8527 5188 8668 5216
rect 8527 5185 8539 5188
rect 8481 5179 8539 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5216 9643 5219
rect 10778 5216 10784 5228
rect 9631 5188 10784 5216
rect 9631 5185 9643 5188
rect 9585 5179 9643 5185
rect 10778 5176 10784 5188
rect 10836 5176 10842 5228
rect 6638 5148 6644 5160
rect 1964 5120 6644 5148
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 10410 5108 10416 5160
rect 10468 5108 10474 5160
rect 10594 5148 10600 5160
rect 10555 5120 10600 5148
rect 10594 5108 10600 5120
rect 10652 5148 10658 5160
rect 10870 5148 10876 5160
rect 10652 5120 10876 5148
rect 10652 5108 10658 5120
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 12621 5151 12679 5157
rect 12621 5148 12633 5151
rect 11112 5120 12633 5148
rect 11112 5108 11118 5120
rect 12621 5117 12633 5120
rect 12667 5117 12679 5151
rect 12621 5111 12679 5117
rect 7098 5080 7104 5092
rect 7059 5052 7104 5080
rect 7098 5040 7104 5052
rect 7156 5040 7162 5092
rect 10042 5080 10048 5092
rect 10003 5052 10048 5080
rect 10042 5040 10048 5052
rect 10100 5040 10106 5092
rect 10428 5080 10456 5108
rect 10505 5083 10563 5089
rect 10505 5080 10517 5083
rect 10428 5052 10517 5080
rect 10505 5049 10517 5052
rect 10551 5049 10563 5083
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 10505 5043 10563 5049
rect 12544 5052 13277 5080
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 1728 4984 1777 5012
rect 1728 4972 1734 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 1765 4975 1823 4981
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5626 5012 5632 5024
rect 5123 4984 5632 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 5721 5015 5779 5021
rect 5721 4981 5733 5015
rect 5767 5012 5779 5015
rect 6178 5012 6184 5024
rect 5767 4984 6184 5012
rect 5767 4981 5779 4984
rect 5721 4975 5779 4981
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10410 5012 10416 5024
rect 9916 4984 10416 5012
rect 9916 4972 9922 4984
rect 10410 4972 10416 4984
rect 10468 4972 10474 5024
rect 10520 5012 10548 5043
rect 10594 5012 10600 5024
rect 10520 4984 10600 5012
rect 10594 4972 10600 4984
rect 10652 5012 10658 5024
rect 11790 5012 11796 5024
rect 10652 4984 11796 5012
rect 10652 4972 10658 4984
rect 11790 4972 11796 4984
rect 11848 4972 11854 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 11977 5015 12035 5021
rect 11977 5012 11989 5015
rect 11940 4984 11989 5012
rect 11940 4972 11946 4984
rect 11977 4981 11989 4984
rect 12023 4981 12035 5015
rect 11977 4975 12035 4981
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 12544 5012 12572 5052
rect 13265 5049 13277 5052
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 12124 4984 12572 5012
rect 13740 5012 13768 5256
rect 14550 5244 14556 5296
rect 14608 5284 14614 5296
rect 14982 5287 15040 5293
rect 14982 5284 14994 5287
rect 14608 5256 14994 5284
rect 14608 5244 14614 5256
rect 14982 5253 14994 5256
rect 15028 5253 15040 5287
rect 14982 5247 15040 5253
rect 18524 5256 19104 5284
rect 14458 5176 14464 5228
rect 14516 5216 14522 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14516 5188 14749 5216
rect 14516 5176 14522 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 15286 5176 15292 5228
rect 15344 5216 15350 5228
rect 18524 5225 18552 5256
rect 17681 5219 17739 5225
rect 17681 5216 17693 5219
rect 15344 5188 17693 5216
rect 15344 5176 15350 5188
rect 17681 5185 17693 5188
rect 17727 5216 17739 5219
rect 18509 5219 18567 5225
rect 18509 5216 18521 5219
rect 17727 5188 18521 5216
rect 17727 5185 17739 5188
rect 17681 5179 17739 5185
rect 18509 5185 18521 5188
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 18693 5219 18751 5225
rect 18693 5185 18705 5219
rect 18739 5185 18751 5219
rect 18693 5179 18751 5185
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 17862 5148 17868 5160
rect 17000 5120 17868 5148
rect 17000 5108 17006 5120
rect 17862 5108 17868 5120
rect 17920 5148 17926 5160
rect 17957 5151 18015 5157
rect 17957 5148 17969 5151
rect 17920 5120 17969 5148
rect 17920 5108 17926 5120
rect 17957 5117 17969 5120
rect 18003 5117 18015 5151
rect 17957 5111 18015 5117
rect 18708 5080 18736 5179
rect 18800 5148 18828 5179
rect 18874 5176 18880 5228
rect 18932 5216 18938 5228
rect 19076 5216 19104 5256
rect 19242 5244 19248 5296
rect 19300 5284 19306 5296
rect 19426 5284 19432 5296
rect 19300 5256 19432 5284
rect 19300 5244 19306 5256
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 19812 5225 19840 5324
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23474 5352 23480 5364
rect 23155 5324 23480 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23474 5312 23480 5324
rect 23532 5312 23538 5364
rect 30374 5312 30380 5364
rect 30432 5312 30438 5364
rect 30834 5352 30840 5364
rect 30795 5324 30840 5352
rect 30834 5312 30840 5324
rect 30892 5312 30898 5364
rect 35621 5355 35679 5361
rect 35621 5321 35633 5355
rect 35667 5352 35679 5355
rect 36078 5352 36084 5364
rect 35667 5324 36084 5352
rect 35667 5321 35679 5324
rect 35621 5315 35679 5321
rect 36078 5312 36084 5324
rect 36136 5312 36142 5364
rect 30392 5231 30420 5312
rect 19613 5219 19671 5225
rect 19613 5216 19625 5219
rect 18932 5188 18977 5216
rect 19076 5188 19625 5216
rect 18932 5176 18938 5188
rect 19613 5185 19625 5188
rect 19659 5185 19671 5219
rect 19613 5179 19671 5185
rect 19797 5219 19855 5225
rect 19797 5185 19809 5219
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 19889 5219 19947 5225
rect 19889 5185 19901 5219
rect 19935 5185 19947 5219
rect 19889 5179 19947 5185
rect 19058 5148 19064 5160
rect 18800 5120 19064 5148
rect 19058 5108 19064 5120
rect 19116 5148 19122 5160
rect 19904 5148 19932 5179
rect 19978 5176 19984 5228
rect 20036 5216 20042 5228
rect 20162 5216 20168 5228
rect 20036 5188 20168 5216
rect 20036 5176 20042 5188
rect 20162 5176 20168 5188
rect 20220 5216 20226 5228
rect 20717 5219 20775 5225
rect 20717 5216 20729 5219
rect 20220 5188 20729 5216
rect 20220 5176 20226 5188
rect 20717 5185 20729 5188
rect 20763 5185 20775 5219
rect 20717 5179 20775 5185
rect 24210 5176 24216 5228
rect 24268 5225 24274 5228
rect 24268 5216 24280 5225
rect 24489 5219 24547 5225
rect 24268 5188 24313 5216
rect 24268 5179 24280 5188
rect 24489 5185 24501 5219
rect 24535 5216 24547 5219
rect 24854 5216 24860 5228
rect 24535 5188 24860 5216
rect 24535 5185 24547 5188
rect 24489 5179 24547 5185
rect 24268 5176 24274 5179
rect 24854 5176 24860 5188
rect 24912 5176 24918 5228
rect 30006 5176 30012 5228
rect 30064 5216 30070 5228
rect 30377 5225 30435 5231
rect 30193 5219 30251 5225
rect 30193 5216 30205 5219
rect 30064 5188 30205 5216
rect 30064 5176 30070 5188
rect 30193 5185 30205 5188
rect 30239 5185 30251 5219
rect 30377 5191 30389 5225
rect 30423 5191 30435 5225
rect 30377 5185 30435 5191
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5185 30527 5219
rect 30193 5179 30251 5185
rect 30469 5179 30527 5185
rect 30561 5219 30619 5225
rect 30561 5185 30573 5219
rect 30607 5191 30788 5219
rect 30607 5185 30619 5191
rect 30561 5179 30619 5185
rect 24946 5148 24952 5160
rect 19116 5120 19932 5148
rect 24907 5120 24952 5148
rect 19116 5108 19122 5120
rect 24946 5108 24952 5120
rect 25004 5108 25010 5160
rect 25225 5151 25283 5157
rect 25225 5117 25237 5151
rect 25271 5148 25283 5151
rect 27154 5148 27160 5160
rect 25271 5120 27160 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 27154 5108 27160 5120
rect 27212 5108 27218 5160
rect 30282 5108 30288 5160
rect 30340 5148 30346 5160
rect 30471 5148 30499 5179
rect 30340 5120 30499 5148
rect 30340 5108 30346 5120
rect 19242 5080 19248 5092
rect 18708 5052 19248 5080
rect 19242 5040 19248 5052
rect 19300 5040 19306 5092
rect 27430 5040 27436 5092
rect 27488 5080 27494 5092
rect 29641 5083 29699 5089
rect 29641 5080 29653 5083
rect 27488 5052 29653 5080
rect 27488 5040 27494 5052
rect 29641 5049 29653 5052
rect 29687 5080 29699 5083
rect 29730 5080 29736 5092
rect 29687 5052 29736 5080
rect 29687 5049 29699 5052
rect 29641 5043 29699 5049
rect 29730 5040 29736 5052
rect 29788 5080 29794 5092
rect 30760 5080 30788 5191
rect 53742 5108 53748 5160
rect 53800 5148 53806 5160
rect 54389 5151 54447 5157
rect 54389 5148 54401 5151
rect 53800 5120 54401 5148
rect 53800 5108 53806 5120
rect 54389 5117 54401 5120
rect 54435 5117 54447 5151
rect 54389 5111 54447 5117
rect 29788 5052 30788 5080
rect 29788 5040 29794 5052
rect 54110 5040 54116 5092
rect 54168 5080 54174 5092
rect 55033 5083 55091 5089
rect 55033 5080 55045 5083
rect 54168 5052 55045 5080
rect 54168 5040 54174 5052
rect 55033 5049 55045 5052
rect 55079 5049 55091 5083
rect 55033 5043 55091 5049
rect 17954 5012 17960 5024
rect 13740 4984 17960 5012
rect 12124 4972 12130 4984
rect 17954 4972 17960 4984
rect 18012 5012 18018 5024
rect 18322 5012 18328 5024
rect 18012 4984 18328 5012
rect 18012 4972 18018 4984
rect 18322 4972 18328 4984
rect 18380 5012 18386 5024
rect 18874 5012 18880 5024
rect 18380 4984 18880 5012
rect 18380 4972 18386 4984
rect 18874 4972 18880 4984
rect 18932 4972 18938 5024
rect 19150 5012 19156 5024
rect 19111 4984 19156 5012
rect 19150 4972 19156 4984
rect 19208 4972 19214 5024
rect 20254 5012 20260 5024
rect 20215 4984 20260 5012
rect 20254 4972 20260 4984
rect 20312 4972 20318 5024
rect 25774 4972 25780 5024
rect 25832 5012 25838 5024
rect 30558 5012 30564 5024
rect 25832 4984 30564 5012
rect 25832 4972 25838 4984
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 53650 4972 53656 5024
rect 53708 5012 53714 5024
rect 53745 5015 53803 5021
rect 53745 5012 53757 5015
rect 53708 4984 53757 5012
rect 53708 4972 53714 4984
rect 53745 4981 53757 4984
rect 53791 4981 53803 5015
rect 58158 5012 58164 5024
rect 58119 4984 58164 5012
rect 53745 4975 53803 4981
rect 58158 4972 58164 4984
rect 58216 4972 58222 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3936 4780 3985 4808
rect 3936 4768 3942 4780
rect 3973 4777 3985 4780
rect 4019 4777 4031 4811
rect 5350 4808 5356 4820
rect 5311 4780 5356 4808
rect 3973 4771 4031 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 6454 4808 6460 4820
rect 6415 4780 6460 4808
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 8205 4811 8263 4817
rect 8205 4777 8217 4811
rect 8251 4808 8263 4811
rect 8294 4808 8300 4820
rect 8251 4780 8300 4808
rect 8251 4777 8263 4780
rect 8205 4771 8263 4777
rect 8294 4768 8300 4780
rect 8352 4808 8358 4820
rect 9217 4811 9275 4817
rect 9217 4808 9229 4811
rect 8352 4780 9229 4808
rect 8352 4768 8358 4780
rect 9217 4777 9229 4780
rect 9263 4777 9275 4811
rect 9217 4771 9275 4777
rect 10134 4768 10140 4820
rect 10192 4808 10198 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 10192 4780 10241 4808
rect 10192 4768 10198 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 10229 4771 10287 4777
rect 10428 4780 10701 4808
rect 3237 4743 3295 4749
rect 3237 4709 3249 4743
rect 3283 4740 3295 4743
rect 5258 4740 5264 4752
rect 3283 4712 5264 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 5258 4700 5264 4712
rect 5316 4700 5322 4752
rect 7098 4700 7104 4752
rect 7156 4740 7162 4752
rect 7285 4743 7343 4749
rect 7285 4740 7297 4743
rect 7156 4712 7297 4740
rect 7156 4700 7162 4712
rect 7285 4709 7297 4712
rect 7331 4709 7343 4743
rect 7285 4703 7343 4709
rect 1946 4632 1952 4684
rect 2004 4632 2010 4684
rect 7300 4672 7328 4703
rect 10042 4700 10048 4752
rect 10100 4740 10106 4752
rect 10428 4740 10456 4780
rect 10689 4777 10701 4780
rect 10735 4808 10747 4811
rect 11514 4808 11520 4820
rect 10735 4780 11520 4808
rect 10735 4777 10747 4780
rect 10689 4771 10747 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 11848 4780 12081 4808
rect 11848 4768 11854 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 12069 4771 12127 4777
rect 12253 4811 12311 4817
rect 12253 4777 12265 4811
rect 12299 4808 12311 4811
rect 12710 4808 12716 4820
rect 12299 4780 12716 4808
rect 12299 4777 12311 4780
rect 12253 4771 12311 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 25774 4808 25780 4820
rect 15764 4780 25780 4808
rect 10594 4740 10600 4752
rect 10100 4712 10456 4740
rect 10555 4712 10600 4740
rect 10100 4700 10106 4712
rect 10594 4700 10600 4712
rect 10652 4700 10658 4752
rect 15764 4740 15792 4780
rect 25774 4768 25780 4780
rect 25832 4768 25838 4820
rect 31202 4808 31208 4820
rect 25884 4780 31208 4808
rect 16942 4740 16948 4752
rect 10888 4712 12112 4740
rect 10888 4684 10916 4712
rect 8113 4675 8171 4681
rect 8113 4672 8125 4675
rect 6380 4644 8125 4672
rect 1964 4604 1992 4632
rect 2590 4604 2596 4616
rect 1964 4576 2596 4604
rect 2590 4564 2596 4576
rect 2648 4564 2654 4616
rect 3050 4613 3056 4616
rect 3045 4604 3056 4613
rect 3011 4576 3056 4604
rect 3045 4567 3056 4576
rect 3050 4564 3056 4567
rect 3108 4564 3114 4616
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4798 4604 4804 4616
rect 4479 4576 4804 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 5442 4604 5448 4616
rect 5403 4576 5448 4604
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6270 4604 6276 4616
rect 6043 4576 6276 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6380 4613 6408 4644
rect 8113 4641 8125 4644
rect 8159 4672 8171 4675
rect 8938 4672 8944 4684
rect 8159 4644 8944 4672
rect 8159 4641 8171 4644
rect 8113 4635 8171 4641
rect 8938 4632 8944 4644
rect 8996 4672 9002 4684
rect 9088 4675 9146 4681
rect 9088 4672 9100 4675
rect 8996 4644 9100 4672
rect 8996 4632 9002 4644
rect 9088 4641 9100 4644
rect 9134 4641 9146 4675
rect 9306 4672 9312 4684
rect 9267 4644 9312 4672
rect 9088 4635 9146 4641
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4641 9459 4675
rect 9401 4635 9459 4641
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4672 10563 4675
rect 10870 4672 10876 4684
rect 10551 4644 10876 4672
rect 10551 4641 10563 4644
rect 10505 4635 10563 4641
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 6730 4604 6736 4616
rect 6687 4576 6736 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 7098 4604 7104 4616
rect 7059 4576 7104 4604
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4604 7803 4607
rect 8018 4604 8024 4616
rect 7791 4576 8024 4604
rect 7791 4573 7803 4576
rect 7745 4567 7803 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4604 8263 4607
rect 8386 4604 8392 4616
rect 8251 4576 8392 4604
rect 8251 4573 8263 4576
rect 8205 4567 8263 4573
rect 8386 4564 8392 4576
rect 8444 4604 8450 4616
rect 9324 4604 9352 4632
rect 8444 4576 9352 4604
rect 8444 4564 8450 4576
rect 1949 4539 2007 4545
rect 1949 4505 1961 4539
rect 1995 4536 2007 4539
rect 5258 4536 5264 4548
rect 1995 4508 5264 4536
rect 1995 4505 2007 4508
rect 1949 4499 2007 4505
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 8036 4536 8064 4564
rect 8846 4536 8852 4548
rect 8036 4508 8852 4536
rect 8846 4496 8852 4508
rect 8904 4536 8910 4548
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 8904 4508 8953 4536
rect 8904 4496 8910 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 9214 4496 9220 4548
rect 9272 4536 9278 4548
rect 9416 4536 9444 4635
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 11072 4644 11744 4672
rect 10410 4564 10416 4616
rect 10468 4604 10474 4616
rect 11072 4613 11100 4644
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10468 4576 11069 4604
rect 10468 4564 10474 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11514 4564 11520 4616
rect 11572 4604 11578 4616
rect 11716 4613 11744 4644
rect 12084 4613 12112 4712
rect 12268 4712 15792 4740
rect 16903 4712 16948 4740
rect 12268 4684 12296 4712
rect 16942 4700 16948 4712
rect 17000 4700 17006 4752
rect 18322 4740 18328 4752
rect 18283 4712 18328 4740
rect 18322 4700 18328 4712
rect 18380 4700 18386 4752
rect 21266 4740 21272 4752
rect 21227 4712 21272 4740
rect 21266 4700 21272 4712
rect 21324 4700 21330 4752
rect 12250 4632 12256 4684
rect 12308 4632 12314 4684
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11572 4576 11621 4604
rect 11572 4564 11578 4576
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4573 11759 4607
rect 11701 4567 11759 4573
rect 12069 4607 12127 4613
rect 12069 4573 12081 4607
rect 12115 4573 12127 4607
rect 12069 4567 12127 4573
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12768 4576 12817 4604
rect 12768 4564 12774 4576
rect 12805 4573 12817 4576
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 14148 4576 14197 4604
rect 14148 4564 14154 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19889 4607 19947 4613
rect 19889 4604 19901 4607
rect 19392 4576 19901 4604
rect 19392 4564 19398 4576
rect 19889 4573 19901 4576
rect 19935 4604 19947 4607
rect 20622 4604 20628 4616
rect 19935 4576 20628 4604
rect 19935 4573 19947 4576
rect 19889 4567 19947 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 24857 4607 24915 4613
rect 24857 4604 24869 4607
rect 20732 4576 24869 4604
rect 9272 4508 9444 4536
rect 9508 4508 12434 4536
rect 9272 4496 9278 4508
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2409 4471 2467 4477
rect 2409 4468 2421 4471
rect 2372 4440 2421 4468
rect 2372 4428 2378 4440
rect 2409 4437 2421 4440
rect 2455 4437 2467 4471
rect 4614 4468 4620 4480
rect 4575 4440 4620 4468
rect 2409 4431 2467 4437
rect 4614 4428 4620 4440
rect 4672 4428 4678 4480
rect 5534 4428 5540 4480
rect 5592 4468 5598 4480
rect 6181 4471 6239 4477
rect 6181 4468 6193 4471
rect 5592 4440 6193 4468
rect 5592 4428 5598 4440
rect 6181 4437 6193 4440
rect 6227 4437 6239 4471
rect 6181 4431 6239 4437
rect 8389 4471 8447 4477
rect 8389 4437 8401 4471
rect 8435 4468 8447 4471
rect 9508 4468 9536 4508
rect 8435 4440 9536 4468
rect 12406 4468 12434 4508
rect 19150 4496 19156 4548
rect 19208 4536 19214 4548
rect 20134 4539 20192 4545
rect 20134 4536 20146 4539
rect 19208 4508 20146 4536
rect 19208 4496 19214 4508
rect 20134 4505 20146 4508
rect 20180 4505 20192 4539
rect 20134 4499 20192 4505
rect 13354 4468 13360 4480
rect 12406 4440 13360 4468
rect 8435 4437 8447 4440
rect 8389 4431 8447 4437
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 13446 4428 13452 4480
rect 13504 4468 13510 4480
rect 13504 4440 13549 4468
rect 13504 4428 13510 4440
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 20732 4468 20760 4576
rect 24857 4573 24869 4576
rect 24903 4604 24915 4607
rect 24946 4604 24952 4616
rect 24903 4576 24952 4604
rect 24903 4573 24915 4576
rect 24857 4567 24915 4573
rect 24946 4564 24952 4576
rect 25004 4564 25010 4616
rect 21266 4496 21272 4548
rect 21324 4536 21330 4548
rect 25884 4536 25912 4780
rect 31202 4768 31208 4780
rect 31260 4768 31266 4820
rect 35897 4811 35955 4817
rect 35897 4777 35909 4811
rect 35943 4808 35955 4811
rect 35986 4808 35992 4820
rect 35943 4780 35992 4808
rect 35943 4777 35955 4780
rect 35897 4771 35955 4777
rect 35986 4768 35992 4780
rect 36044 4768 36050 4820
rect 27154 4700 27160 4752
rect 27212 4740 27218 4752
rect 27212 4712 29408 4740
rect 27212 4700 27218 4712
rect 27614 4632 27620 4684
rect 27672 4632 27678 4684
rect 29270 4672 29276 4684
rect 28000 4644 29276 4672
rect 26050 4604 26056 4616
rect 25963 4576 26056 4604
rect 26050 4564 26056 4576
rect 26108 4604 26114 4616
rect 26510 4604 26516 4616
rect 26108 4576 26516 4604
rect 26108 4564 26114 4576
rect 26510 4564 26516 4576
rect 26568 4604 26574 4616
rect 26743 4607 26801 4613
rect 26743 4604 26755 4607
rect 26568 4576 26755 4604
rect 26568 4564 26574 4576
rect 26743 4573 26755 4576
rect 26789 4573 26801 4607
rect 26878 4604 26884 4616
rect 26839 4576 26884 4604
rect 26743 4567 26801 4573
rect 26878 4564 26884 4576
rect 26936 4564 26942 4616
rect 26973 4607 27031 4613
rect 26973 4573 26985 4607
rect 27019 4573 27031 4607
rect 27154 4604 27160 4616
rect 27115 4576 27160 4604
rect 26973 4567 27031 4573
rect 21324 4508 25912 4536
rect 21324 4496 21330 4508
rect 17920 4440 20760 4468
rect 17920 4428 17926 4440
rect 26326 4428 26332 4480
rect 26384 4468 26390 4480
rect 26513 4471 26571 4477
rect 26513 4468 26525 4471
rect 26384 4440 26525 4468
rect 26384 4428 26390 4440
rect 26513 4437 26525 4440
rect 26559 4437 26571 4471
rect 26896 4468 26924 4564
rect 26988 4536 27016 4567
rect 27154 4564 27160 4576
rect 27212 4564 27218 4616
rect 27632 4604 27660 4632
rect 28000 4613 28028 4644
rect 29270 4632 29276 4644
rect 29328 4632 29334 4684
rect 27801 4607 27859 4613
rect 27801 4604 27813 4607
rect 27632 4576 27813 4604
rect 27801 4573 27813 4576
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 27985 4607 28043 4613
rect 27985 4573 27997 4607
rect 28031 4573 28043 4607
rect 29380 4604 29408 4712
rect 30558 4700 30564 4752
rect 30616 4740 30622 4752
rect 30653 4743 30711 4749
rect 30653 4740 30665 4743
rect 30616 4712 30665 4740
rect 30616 4700 30622 4712
rect 30653 4709 30665 4712
rect 30699 4709 30711 4743
rect 30653 4703 30711 4709
rect 52178 4700 52184 4752
rect 52236 4740 52242 4752
rect 52825 4743 52883 4749
rect 52825 4740 52837 4743
rect 52236 4712 52837 4740
rect 52236 4700 52242 4712
rect 52825 4709 52837 4712
rect 52871 4709 52883 4743
rect 52825 4703 52883 4709
rect 53926 4700 53932 4752
rect 53984 4740 53990 4752
rect 55309 4743 55367 4749
rect 55309 4740 55321 4743
rect 53984 4712 55321 4740
rect 53984 4700 53990 4712
rect 55309 4709 55321 4712
rect 55355 4709 55367 4743
rect 55309 4703 55367 4709
rect 31481 4675 31539 4681
rect 31481 4672 31493 4675
rect 30208 4644 31493 4672
rect 30006 4604 30012 4616
rect 29380 4576 30012 4604
rect 27985 4567 28043 4573
rect 30006 4564 30012 4576
rect 30064 4564 30070 4616
rect 30208 4613 30236 4644
rect 31481 4641 31493 4644
rect 31527 4641 31539 4675
rect 37274 4672 37280 4684
rect 37235 4644 37280 4672
rect 31481 4635 31539 4641
rect 37274 4632 37280 4644
rect 37332 4632 37338 4684
rect 53190 4632 53196 4684
rect 53248 4672 53254 4684
rect 54113 4675 54171 4681
rect 54113 4672 54125 4675
rect 53248 4644 54125 4672
rect 53248 4632 53254 4644
rect 54113 4641 54125 4644
rect 54159 4641 54171 4675
rect 54113 4635 54171 4641
rect 54294 4632 54300 4684
rect 54352 4672 54358 4684
rect 55953 4675 56011 4681
rect 55953 4672 55965 4675
rect 54352 4644 55965 4672
rect 54352 4632 54358 4644
rect 55953 4641 55965 4644
rect 55999 4641 56011 4675
rect 55953 4635 56011 4641
rect 30193 4607 30251 4613
rect 30193 4573 30205 4607
rect 30239 4573 30251 4607
rect 30193 4567 30251 4573
rect 30285 4607 30343 4613
rect 30285 4573 30297 4607
rect 30331 4573 30343 4607
rect 30285 4567 30343 4573
rect 27617 4539 27675 4545
rect 27617 4536 27629 4539
rect 26988 4508 27629 4536
rect 27617 4505 27629 4508
rect 27663 4505 27675 4539
rect 30300 4536 30328 4567
rect 30374 4564 30380 4616
rect 30432 4604 30438 4616
rect 30650 4604 30656 4616
rect 30432 4576 30656 4604
rect 30432 4564 30438 4576
rect 30650 4564 30656 4576
rect 30708 4564 30714 4616
rect 30926 4564 30932 4616
rect 30984 4604 30990 4616
rect 31297 4607 31355 4613
rect 31297 4604 31309 4607
rect 30984 4576 31309 4604
rect 30984 4564 30990 4576
rect 31297 4573 31309 4576
rect 31343 4604 31355 4607
rect 31570 4604 31576 4616
rect 31343 4576 31576 4604
rect 31343 4573 31355 4576
rect 31297 4567 31355 4573
rect 31570 4564 31576 4576
rect 31628 4564 31634 4616
rect 36998 4564 37004 4616
rect 37056 4613 37062 4616
rect 37056 4604 37068 4613
rect 37056 4576 37101 4604
rect 37056 4567 37068 4576
rect 37056 4564 37062 4567
rect 52086 4564 52092 4616
rect 52144 4604 52150 4616
rect 52181 4607 52239 4613
rect 52181 4604 52193 4607
rect 52144 4576 52193 4604
rect 52144 4564 52150 4576
rect 52181 4573 52193 4576
rect 52227 4573 52239 4607
rect 52181 4567 52239 4573
rect 52638 4564 52644 4616
rect 52696 4604 52702 4616
rect 53469 4607 53527 4613
rect 53469 4604 53481 4607
rect 52696 4576 53481 4604
rect 52696 4564 52702 4576
rect 53469 4573 53481 4576
rect 53515 4573 53527 4607
rect 53469 4567 53527 4573
rect 30466 4536 30472 4548
rect 27617 4499 27675 4505
rect 28828 4508 30472 4536
rect 28828 4468 28856 4508
rect 30466 4496 30472 4508
rect 30524 4496 30530 4548
rect 31113 4539 31171 4545
rect 31113 4536 31125 4539
rect 30576 4508 31125 4536
rect 28994 4468 29000 4480
rect 26896 4440 28856 4468
rect 28955 4440 29000 4468
rect 26513 4431 26571 4437
rect 28994 4428 29000 4440
rect 29052 4428 29058 4480
rect 29270 4428 29276 4480
rect 29328 4468 29334 4480
rect 30576 4468 30604 4508
rect 31113 4505 31125 4508
rect 31159 4505 31171 4539
rect 31113 4499 31171 4505
rect 29328 4440 30604 4468
rect 29328 4428 29334 4440
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 3786 4264 3792 4276
rect 2746 4236 3792 4264
rect 2590 4156 2596 4208
rect 2648 4196 2654 4208
rect 2746 4196 2774 4236
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 6575 4267 6633 4273
rect 4028 4236 6500 4264
rect 4028 4224 4034 4236
rect 5000 4205 5028 4236
rect 2648 4168 2774 4196
rect 4985 4199 5043 4205
rect 2648 4156 2654 4168
rect 4985 4165 4997 4199
rect 5031 4165 5043 4199
rect 4985 4159 5043 4165
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 6365 4199 6423 4205
rect 6365 4196 6377 4199
rect 5408 4168 6377 4196
rect 5408 4156 5414 4168
rect 6365 4165 6377 4168
rect 6411 4165 6423 4199
rect 6472 4196 6500 4236
rect 6575 4233 6587 4267
rect 6621 4264 6633 4267
rect 6822 4264 6828 4276
rect 6621 4236 6828 4264
rect 6621 4233 6633 4236
rect 6575 4227 6633 4233
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 7558 4264 7564 4276
rect 7519 4236 7564 4264
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 28994 4224 29000 4276
rect 29052 4264 29058 4276
rect 30374 4264 30380 4276
rect 29052 4236 30380 4264
rect 29052 4224 29058 4236
rect 30374 4224 30380 4236
rect 30432 4224 30438 4276
rect 31570 4264 31576 4276
rect 31531 4236 31576 4264
rect 31570 4224 31576 4236
rect 31628 4224 31634 4276
rect 6914 4196 6920 4208
rect 6472 4168 6920 4196
rect 6365 4159 6423 4165
rect 6914 4156 6920 4168
rect 6972 4156 6978 4208
rect 19604 4199 19662 4205
rect 19604 4165 19616 4199
rect 19650 4196 19662 4199
rect 20254 4196 20260 4208
rect 19650 4168 20260 4196
rect 19650 4165 19662 4168
rect 19604 4159 19662 4165
rect 20254 4156 20260 4168
rect 20312 4156 20318 4208
rect 30460 4199 30518 4205
rect 30460 4165 30472 4199
rect 30506 4196 30518 4199
rect 30558 4196 30564 4208
rect 30506 4168 30564 4196
rect 30506 4165 30518 4168
rect 30460 4159 30518 4165
rect 30558 4156 30564 4168
rect 30616 4156 30622 4208
rect 1670 4128 1676 4140
rect 1631 4100 1676 4128
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4088 2378 4140
rect 2406 4088 2412 4140
rect 2464 4128 2470 4140
rect 2464 4100 2509 4128
rect 2464 4088 2470 4100
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 2924 4100 3157 4128
rect 2924 4088 2930 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4120 4100 4353 4128
rect 4120 4088 4126 4100
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6546 4128 6552 4140
rect 5859 4100 6552 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6546 4088 6552 4100
rect 6604 4128 6610 4140
rect 7282 4128 7288 4140
rect 6604 4100 7288 4128
rect 6604 4088 6610 4100
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7524 4100 7757 4128
rect 7524 4088 7530 4100
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4128 7987 4131
rect 8294 4128 8300 4140
rect 7975 4100 8300 4128
rect 7975 4097 7987 4100
rect 7929 4091 7987 4097
rect 3510 4020 3516 4072
rect 3568 4060 3574 4072
rect 4801 4063 4859 4069
rect 4801 4060 4813 4063
rect 3568 4032 4813 4060
rect 3568 4020 3574 4032
rect 4801 4029 4813 4032
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 6362 4060 6368 4072
rect 4948 4032 6368 4060
rect 4948 4020 4954 4032
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 2958 3992 2964 4004
rect 2919 3964 2964 3992
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3992 4215 3995
rect 4522 3992 4528 4004
rect 4203 3964 4528 3992
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 4614 3952 4620 4004
rect 4672 3992 4678 4004
rect 4672 3964 6592 3992
rect 4672 3952 4678 3964
rect 1857 3927 1915 3933
rect 1857 3893 1869 3927
rect 1903 3924 1915 3927
rect 1946 3924 1952 3936
rect 1903 3896 1952 3924
rect 1903 3893 1915 3896
rect 1857 3887 1915 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 5350 3884 5356 3936
rect 5408 3924 5414 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5408 3896 5641 3924
rect 5408 3884 5414 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 6270 3924 6276 3936
rect 5776 3896 6276 3924
rect 5776 3884 5782 3896
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6564 3933 6592 3964
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 6733 3995 6791 4001
rect 6733 3992 6745 3995
rect 6696 3964 6745 3992
rect 6696 3952 6702 3964
rect 6733 3961 6745 3964
rect 6779 3961 6791 3995
rect 7760 3992 7788 4091
rect 8294 4088 8300 4100
rect 8352 4128 8358 4140
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8352 4100 8585 4128
rect 8352 4088 8358 4100
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 8938 4128 8944 4140
rect 8899 4100 8944 4128
rect 8573 4091 8631 4097
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4128 10011 4131
rect 11606 4128 11612 4140
rect 9999 4100 11612 4128
rect 9999 4097 10011 4100
rect 9953 4091 10011 4097
rect 11606 4088 11612 4100
rect 11664 4088 11670 4140
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 15013 4131 15071 4137
rect 15013 4128 15025 4131
rect 14792 4100 15025 4128
rect 14792 4088 14798 4100
rect 15013 4097 15025 4100
rect 15059 4128 15071 4131
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 15059 4100 15485 4128
rect 15059 4097 15071 4100
rect 15013 4091 15071 4097
rect 15473 4097 15485 4100
rect 15519 4097 15531 4131
rect 19334 4128 19340 4140
rect 19295 4100 19340 4128
rect 15473 4091 15531 4097
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 30190 4128 30196 4140
rect 30151 4100 30196 4128
rect 30190 4088 30196 4100
rect 30248 4088 30254 4140
rect 32766 4088 32772 4140
rect 32824 4128 32830 4140
rect 33505 4131 33563 4137
rect 33505 4128 33517 4131
rect 32824 4100 33517 4128
rect 32824 4088 32830 4100
rect 33505 4097 33517 4100
rect 33551 4097 33563 4131
rect 33505 4091 33563 4097
rect 33772 4131 33830 4137
rect 33772 4097 33784 4131
rect 33818 4128 33830 4131
rect 34330 4128 34336 4140
rect 33818 4100 34336 4128
rect 33818 4097 33830 4100
rect 33772 4091 33830 4097
rect 34330 4088 34336 4100
rect 34388 4088 34394 4140
rect 53006 4088 53012 4140
rect 53064 4128 53070 4140
rect 54665 4131 54723 4137
rect 54665 4128 54677 4131
rect 53064 4100 54677 4128
rect 53064 4088 53070 4100
rect 54665 4097 54677 4100
rect 54711 4097 54723 4131
rect 54665 4091 54723 4097
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8444 4032 8493 4060
rect 8444 4020 8450 4032
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 10042 4060 10048 4072
rect 8481 4023 8539 4029
rect 9048 4032 10048 4060
rect 9048 3992 9076 4032
rect 10042 4020 10048 4032
rect 10100 4020 10106 4072
rect 51810 4020 51816 4072
rect 51868 4060 51874 4072
rect 52733 4063 52791 4069
rect 52733 4060 52745 4063
rect 51868 4032 52745 4060
rect 51868 4020 51874 4032
rect 52733 4029 52745 4032
rect 52779 4029 52791 4063
rect 52733 4023 52791 4029
rect 54018 4020 54024 4072
rect 54076 4060 54082 4072
rect 55953 4063 56011 4069
rect 55953 4060 55965 4063
rect 54076 4032 55965 4060
rect 54076 4020 54082 4032
rect 55953 4029 55965 4032
rect 55999 4029 56011 4063
rect 55953 4023 56011 4029
rect 7760 3964 9076 3992
rect 9125 3995 9183 4001
rect 6733 3955 6791 3961
rect 9125 3961 9137 3995
rect 9171 3992 9183 3995
rect 9306 3992 9312 4004
rect 9171 3964 9312 3992
rect 9171 3961 9183 3964
rect 9125 3955 9183 3961
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 34885 3995 34943 4001
rect 34885 3961 34897 3995
rect 34931 3992 34943 3995
rect 35342 3992 35348 4004
rect 34931 3964 35348 3992
rect 34931 3961 34943 3964
rect 34885 3955 34943 3961
rect 35342 3952 35348 3964
rect 35400 3952 35406 4004
rect 52822 3952 52828 4004
rect 52880 3992 52886 4004
rect 52880 3964 54064 3992
rect 52880 3952 52886 3964
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3893 6607 3927
rect 6549 3887 6607 3893
rect 7929 3927 7987 3933
rect 7929 3893 7941 3927
rect 7975 3924 7987 3927
rect 8386 3924 8392 3936
rect 7975 3896 8392 3924
rect 7975 3893 7987 3896
rect 7929 3887 7987 3893
rect 8386 3884 8392 3896
rect 8444 3924 8450 3936
rect 8570 3924 8576 3936
rect 8444 3896 8576 3924
rect 8444 3884 8450 3896
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 8941 3927 8999 3933
rect 8941 3924 8953 3927
rect 8904 3896 8953 3924
rect 8904 3884 8910 3896
rect 8941 3893 8953 3896
rect 8987 3893 8999 3927
rect 8941 3887 8999 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9272 3896 9781 3924
rect 9272 3884 9278 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 9769 3887 9827 3893
rect 10965 3927 11023 3933
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 11606 3924 11612 3936
rect 11011 3896 11612 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 11606 3884 11612 3896
rect 11664 3884 11670 3936
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 12158 3924 12164 3936
rect 11839 3896 12164 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13081 3927 13139 3933
rect 12492 3896 12537 3924
rect 12492 3884 12498 3896
rect 13081 3893 13093 3927
rect 13127 3924 13139 3927
rect 13262 3924 13268 3936
rect 13127 3896 13268 3924
rect 13127 3893 13139 3896
rect 13081 3887 13139 3893
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13725 3927 13783 3933
rect 13725 3893 13737 3927
rect 13771 3924 13783 3927
rect 13814 3924 13820 3936
rect 13771 3896 13820 3924
rect 13771 3893 13783 3896
rect 13725 3887 13783 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14366 3924 14372 3936
rect 14327 3896 14372 3924
rect 14366 3884 14372 3896
rect 14424 3884 14430 3936
rect 14826 3924 14832 3936
rect 14787 3896 14832 3924
rect 14826 3884 14832 3896
rect 14884 3884 14890 3936
rect 20717 3927 20775 3933
rect 20717 3893 20729 3927
rect 20763 3924 20775 3927
rect 20898 3924 20904 3936
rect 20763 3896 20904 3924
rect 20763 3893 20775 3896
rect 20717 3887 20775 3893
rect 20898 3884 20904 3896
rect 20956 3924 20962 3936
rect 29454 3924 29460 3936
rect 20956 3896 29460 3924
rect 20956 3884 20962 3896
rect 29454 3884 29460 3896
rect 29512 3884 29518 3936
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 51169 3927 51227 3933
rect 51169 3924 51181 3927
rect 51132 3896 51181 3924
rect 51132 3884 51138 3896
rect 51169 3893 51181 3896
rect 51215 3893 51227 3927
rect 51169 3887 51227 3893
rect 51350 3884 51356 3936
rect 51408 3924 51414 3936
rect 51813 3927 51871 3933
rect 51813 3924 51825 3927
rect 51408 3896 51825 3924
rect 51408 3884 51414 3896
rect 51813 3893 51825 3896
rect 51859 3893 51871 3927
rect 51813 3887 51871 3893
rect 52454 3884 52460 3936
rect 52512 3924 52518 3936
rect 54036 3933 54064 3964
rect 53377 3927 53435 3933
rect 53377 3924 53389 3927
rect 52512 3896 53389 3924
rect 52512 3884 52518 3896
rect 53377 3893 53389 3896
rect 53423 3893 53435 3927
rect 53377 3887 53435 3893
rect 54021 3927 54079 3933
rect 54021 3893 54033 3927
rect 54067 3893 54079 3927
rect 55306 3924 55312 3936
rect 55267 3896 55312 3924
rect 54021 3887 54079 3893
rect 55306 3884 55312 3896
rect 55364 3884 55370 3936
rect 58161 3927 58219 3933
rect 58161 3893 58173 3927
rect 58207 3924 58219 3927
rect 58434 3924 58440 3936
rect 58207 3896 58440 3924
rect 58207 3893 58219 3896
rect 58161 3887 58219 3893
rect 58434 3884 58440 3896
rect 58492 3884 58498 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 2130 3720 2136 3732
rect 1872 3692 2136 3720
rect 1872 3593 1900 3692
rect 2130 3680 2136 3692
rect 2188 3720 2194 3732
rect 5166 3720 5172 3732
rect 2188 3692 3832 3720
rect 5127 3692 5172 3720
rect 2188 3680 2194 3692
rect 3804 3593 3832 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 5905 3723 5963 3729
rect 5905 3720 5917 3723
rect 5684 3692 5917 3720
rect 5684 3680 5690 3692
rect 5905 3689 5917 3692
rect 5951 3689 5963 3723
rect 5905 3683 5963 3689
rect 6089 3723 6147 3729
rect 6089 3689 6101 3723
rect 6135 3720 6147 3723
rect 7558 3720 7564 3732
rect 6135 3692 7564 3720
rect 6135 3689 6147 3692
rect 6089 3683 6147 3689
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 8662 3720 8668 3732
rect 7708 3692 8668 3720
rect 7708 3680 7714 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 9309 3723 9367 3729
rect 9309 3720 9321 3723
rect 9180 3692 9321 3720
rect 9180 3680 9186 3692
rect 9309 3689 9321 3692
rect 9355 3689 9367 3723
rect 9766 3720 9772 3732
rect 9727 3692 9772 3720
rect 9309 3683 9367 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 10505 3723 10563 3729
rect 10505 3689 10517 3723
rect 10551 3720 10563 3723
rect 10962 3720 10968 3732
rect 10551 3692 10968 3720
rect 10551 3689 10563 3692
rect 10505 3683 10563 3689
rect 10962 3680 10968 3692
rect 11020 3720 11026 3732
rect 26050 3720 26056 3732
rect 11020 3692 26056 3720
rect 11020 3680 11026 3692
rect 26050 3680 26056 3692
rect 26108 3680 26114 3732
rect 27433 3723 27491 3729
rect 27433 3689 27445 3723
rect 27479 3720 27491 3723
rect 27614 3720 27620 3732
rect 27479 3692 27620 3720
rect 27479 3689 27491 3692
rect 27433 3683 27491 3689
rect 27614 3680 27620 3692
rect 27672 3680 27678 3732
rect 52730 3680 52736 3732
rect 52788 3720 52794 3732
rect 52788 3692 55214 3720
rect 52788 3680 52794 3692
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 6546 3652 6552 3664
rect 5500 3624 6552 3652
rect 5500 3612 5506 3624
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 8294 3612 8300 3664
rect 8352 3652 8358 3664
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 8352 3624 8953 3652
rect 8352 3612 8358 3624
rect 8941 3621 8953 3624
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 9401 3655 9459 3661
rect 9401 3621 9413 3655
rect 9447 3621 9459 3655
rect 9401 3615 9459 3621
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 6730 3544 6736 3596
rect 6788 3584 6794 3596
rect 6825 3587 6883 3593
rect 6825 3584 6837 3587
rect 6788 3556 6837 3584
rect 6788 3544 6794 3556
rect 6825 3553 6837 3556
rect 6871 3553 6883 3587
rect 6825 3547 6883 3553
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 9416 3584 9444 3615
rect 11238 3612 11244 3664
rect 11296 3652 11302 3664
rect 12250 3652 12256 3664
rect 11296 3624 12256 3652
rect 11296 3612 11302 3624
rect 12250 3612 12256 3624
rect 12308 3612 12314 3664
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14093 3655 14151 3661
rect 14093 3652 14105 3655
rect 14056 3624 14105 3652
rect 14056 3612 14062 3624
rect 14093 3621 14105 3624
rect 14139 3621 14151 3655
rect 14093 3615 14151 3621
rect 14829 3655 14887 3661
rect 14829 3621 14841 3655
rect 14875 3621 14887 3655
rect 14829 3615 14887 3621
rect 8720 3556 9444 3584
rect 8720 3544 8726 3556
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 12897 3587 12955 3593
rect 9548 3556 9593 3584
rect 9548 3544 9554 3556
rect 12897 3553 12909 3587
rect 12943 3584 12955 3587
rect 13538 3584 13544 3596
rect 12943 3556 13544 3584
rect 12943 3553 12955 3556
rect 12897 3547 12955 3553
rect 13538 3544 13544 3556
rect 13596 3544 13602 3596
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 14844 3584 14872 3615
rect 46290 3612 46296 3664
rect 46348 3652 46354 3664
rect 46937 3655 46995 3661
rect 46937 3652 46949 3655
rect 46348 3624 46949 3652
rect 46348 3612 46354 3624
rect 46937 3621 46949 3624
rect 46983 3621 46995 3655
rect 46937 3615 46995 3621
rect 51442 3612 51448 3664
rect 51500 3652 51506 3664
rect 52825 3655 52883 3661
rect 52825 3652 52837 3655
rect 51500 3624 52837 3652
rect 51500 3612 51506 3624
rect 52825 3621 52837 3624
rect 52871 3621 52883 3655
rect 55186 3652 55214 3692
rect 55309 3655 55367 3661
rect 55309 3652 55321 3655
rect 55186 3624 55321 3652
rect 52825 3615 52883 3621
rect 55309 3621 55321 3624
rect 55355 3621 55367 3655
rect 55309 3615 55367 3621
rect 13964 3556 14872 3584
rect 13964 3544 13970 3556
rect 24854 3544 24860 3596
rect 24912 3584 24918 3596
rect 26053 3587 26111 3593
rect 26053 3584 26065 3587
rect 24912 3556 26065 3584
rect 24912 3544 24918 3556
rect 26053 3553 26065 3556
rect 26099 3553 26111 3587
rect 26053 3547 26111 3553
rect 50798 3544 50804 3596
rect 50856 3584 50862 3596
rect 51537 3587 51595 3593
rect 51537 3584 51549 3587
rect 50856 3556 51549 3584
rect 50856 3544 50862 3556
rect 51537 3553 51549 3556
rect 51583 3553 51595 3587
rect 51537 3547 51595 3553
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 53469 3587 53527 3593
rect 53469 3584 53481 3587
rect 51684 3556 53481 3584
rect 51684 3544 51690 3556
rect 53469 3553 53481 3556
rect 53515 3553 53527 3587
rect 53469 3547 53527 3553
rect 53834 3544 53840 3596
rect 53892 3584 53898 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 53892 3556 56609 3584
rect 53892 3544 53898 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 1946 3476 1952 3528
rect 2004 3516 2010 3528
rect 2113 3519 2171 3525
rect 2113 3516 2125 3519
rect 2004 3488 2125 3516
rect 2004 3476 2010 3488
rect 2113 3485 2125 3488
rect 2159 3485 2171 3519
rect 2113 3479 2171 3485
rect 4056 3519 4114 3525
rect 4056 3485 4068 3519
rect 4102 3516 4114 3519
rect 5074 3516 5080 3528
rect 4102 3488 5080 3516
rect 4102 3485 4114 3488
rect 4056 3479 4114 3485
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 6454 3516 6460 3528
rect 5316 3488 6460 3516
rect 5316 3476 5322 3488
rect 6454 3476 6460 3488
rect 6512 3516 6518 3528
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 6512 3488 6561 3516
rect 6512 3476 6518 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3516 8355 3519
rect 8478 3516 8484 3528
rect 8343 3488 8484 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 10318 3516 10324 3528
rect 9088 3488 10324 3516
rect 9088 3476 9094 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3516 11115 3519
rect 11146 3516 11152 3528
rect 11103 3488 11152 3516
rect 11103 3485 11115 3488
rect 11057 3479 11115 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12986 3516 12992 3528
rect 12299 3488 12992 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 14182 3516 14188 3528
rect 13403 3488 14188 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 15381 3519 15439 3525
rect 15381 3516 15393 3519
rect 15252 3488 15393 3516
rect 15252 3476 15258 3488
rect 15381 3485 15393 3488
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15988 3488 16037 3516
rect 15988 3476 15994 3488
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 16025 3479 16083 3485
rect 16758 3476 16764 3528
rect 16816 3516 16822 3528
rect 16853 3519 16911 3525
rect 16853 3516 16865 3519
rect 16816 3488 16865 3516
rect 16816 3476 16822 3488
rect 16853 3485 16865 3488
rect 16899 3485 16911 3519
rect 16853 3479 16911 3485
rect 17586 3476 17592 3528
rect 17644 3516 17650 3528
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17644 3488 17693 3516
rect 17644 3476 17650 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18472 3488 18521 3516
rect 18472 3476 18478 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 19484 3488 19625 3516
rect 19484 3476 19490 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 20441 3519 20499 3525
rect 20441 3516 20453 3519
rect 20404 3488 20453 3516
rect 20404 3476 20410 3488
rect 20441 3485 20453 3488
rect 20487 3485 20499 3519
rect 20441 3479 20499 3485
rect 21174 3476 21180 3528
rect 21232 3516 21238 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21232 3488 21281 3516
rect 21232 3476 21238 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21269 3479 21327 3485
rect 22189 3519 22247 3525
rect 22189 3485 22201 3519
rect 22235 3516 22247 3519
rect 22278 3516 22284 3528
rect 22235 3488 22284 3516
rect 22235 3485 22247 3488
rect 22189 3479 22247 3485
rect 22278 3476 22284 3488
rect 22336 3476 22342 3528
rect 22554 3476 22560 3528
rect 22612 3516 22618 3528
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 22612 3488 22661 3516
rect 22612 3476 22618 3488
rect 22649 3485 22661 3488
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 23382 3476 23388 3528
rect 23440 3516 23446 3528
rect 23477 3519 23535 3525
rect 23477 3516 23489 3519
rect 23440 3488 23489 3516
rect 23440 3476 23446 3488
rect 23477 3485 23489 3488
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 24486 3476 24492 3528
rect 24544 3516 24550 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 24544 3488 24593 3516
rect 24544 3476 24550 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 25590 3516 25596 3528
rect 25551 3488 25596 3516
rect 24581 3479 24639 3485
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 26326 3525 26332 3528
rect 26320 3516 26332 3525
rect 26287 3488 26332 3516
rect 26320 3479 26332 3488
rect 26326 3476 26332 3479
rect 26384 3476 26390 3528
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 27893 3519 27951 3525
rect 27893 3516 27905 3519
rect 27580 3488 27905 3516
rect 27580 3476 27586 3488
rect 27893 3485 27905 3488
rect 27939 3485 27951 3519
rect 27893 3479 27951 3485
rect 28626 3476 28632 3528
rect 28684 3516 28690 3528
rect 28721 3519 28779 3525
rect 28721 3516 28733 3519
rect 28684 3488 28733 3516
rect 28684 3476 28690 3488
rect 28721 3485 28733 3488
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34793 3519 34851 3525
rect 34793 3516 34805 3519
rect 34756 3488 34805 3516
rect 34756 3476 34762 3488
rect 34793 3485 34805 3488
rect 34839 3485 34851 3519
rect 34793 3479 34851 3485
rect 35342 3476 35348 3528
rect 35400 3516 35406 3528
rect 35437 3519 35495 3525
rect 35437 3516 35449 3519
rect 35400 3488 35449 3516
rect 35400 3476 35406 3488
rect 35437 3485 35449 3488
rect 35483 3485 35495 3519
rect 35437 3479 35495 3485
rect 35802 3476 35808 3528
rect 35860 3516 35866 3528
rect 36081 3519 36139 3525
rect 36081 3516 36093 3519
rect 35860 3488 36093 3516
rect 35860 3476 35866 3488
rect 36081 3485 36093 3488
rect 36127 3485 36139 3519
rect 36081 3479 36139 3485
rect 36630 3476 36636 3528
rect 36688 3516 36694 3528
rect 36725 3519 36783 3525
rect 36725 3516 36737 3519
rect 36688 3488 36737 3516
rect 36688 3476 36694 3488
rect 36725 3485 36737 3488
rect 36771 3485 36783 3519
rect 36725 3479 36783 3485
rect 37458 3476 37464 3528
rect 37516 3516 37522 3528
rect 37553 3519 37611 3525
rect 37553 3516 37565 3519
rect 37516 3488 37565 3516
rect 37516 3476 37522 3488
rect 37553 3485 37565 3488
rect 37599 3485 37611 3519
rect 37553 3479 37611 3485
rect 38562 3476 38568 3528
rect 38620 3516 38626 3528
rect 38657 3519 38715 3525
rect 38657 3516 38669 3519
rect 38620 3488 38669 3516
rect 38620 3476 38626 3488
rect 38657 3485 38669 3488
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 40000 3488 40049 3516
rect 40000 3476 40006 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40494 3476 40500 3528
rect 40552 3516 40558 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40552 3488 40693 3516
rect 40552 3476 40558 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 40681 3479 40739 3485
rect 41046 3476 41052 3528
rect 41104 3516 41110 3528
rect 41325 3519 41383 3525
rect 41325 3516 41337 3519
rect 41104 3488 41337 3516
rect 41104 3476 41110 3488
rect 41325 3485 41337 3488
rect 41371 3485 41383 3519
rect 41325 3479 41383 3485
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 42521 3519 42579 3525
rect 42521 3516 42533 3519
rect 42484 3488 42533 3516
rect 42484 3476 42490 3488
rect 42521 3485 42533 3488
rect 42567 3485 42579 3519
rect 42521 3479 42579 3485
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 43165 3519 43223 3525
rect 43165 3516 43177 3519
rect 42760 3488 43177 3516
rect 42760 3476 42766 3488
rect 43165 3485 43177 3488
rect 43211 3485 43223 3519
rect 43165 3479 43223 3485
rect 44358 3476 44364 3528
rect 44416 3516 44422 3528
rect 45005 3519 45063 3525
rect 45005 3516 45017 3519
rect 44416 3488 45017 3516
rect 44416 3476 44422 3488
rect 45005 3485 45017 3488
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 45186 3476 45192 3528
rect 45244 3516 45250 3528
rect 45649 3519 45707 3525
rect 45649 3516 45661 3519
rect 45244 3488 45661 3516
rect 45244 3476 45250 3488
rect 45649 3485 45661 3488
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 46014 3476 46020 3528
rect 46072 3516 46078 3528
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 46072 3488 46305 3516
rect 46072 3476 46078 3488
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 47670 3476 47676 3528
rect 47728 3516 47734 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47728 3488 47777 3516
rect 47728 3476 47734 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 48222 3476 48228 3528
rect 48280 3516 48286 3528
rect 48409 3519 48467 3525
rect 48409 3516 48421 3519
rect 48280 3488 48421 3516
rect 48280 3476 48286 3488
rect 48409 3485 48421 3488
rect 48455 3485 48467 3519
rect 48409 3479 48467 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50249 3519 50307 3525
rect 50249 3516 50261 3519
rect 50212 3488 50261 3516
rect 50212 3476 50218 3488
rect 50249 3485 50261 3488
rect 50295 3485 50307 3519
rect 50249 3479 50307 3485
rect 50614 3476 50620 3528
rect 50672 3516 50678 3528
rect 50893 3519 50951 3525
rect 50893 3516 50905 3519
rect 50672 3488 50905 3516
rect 50672 3476 50678 3488
rect 50893 3485 50905 3488
rect 50939 3485 50951 3519
rect 50893 3479 50951 3485
rect 51166 3476 51172 3528
rect 51224 3516 51230 3528
rect 52181 3519 52239 3525
rect 52181 3516 52193 3519
rect 51224 3488 52193 3516
rect 51224 3476 51230 3488
rect 52181 3485 52193 3488
rect 52227 3485 52239 3519
rect 52181 3479 52239 3485
rect 52270 3476 52276 3528
rect 52328 3516 52334 3528
rect 54113 3519 54171 3525
rect 54113 3516 54125 3519
rect 52328 3488 54125 3516
rect 52328 3476 52334 3488
rect 54113 3485 54125 3488
rect 54159 3485 54171 3519
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 54113 3479 54171 3485
rect 55186 3488 55965 3516
rect 5718 3448 5724 3460
rect 5679 3420 5724 3448
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 5937 3451 5995 3457
rect 5937 3417 5949 3451
rect 5983 3448 5995 3451
rect 6638 3448 6644 3460
rect 5983 3420 6644 3448
rect 5983 3417 5995 3420
rect 5937 3411 5995 3417
rect 6638 3408 6644 3420
rect 6696 3408 6702 3460
rect 8386 3408 8392 3460
rect 8444 3448 8450 3460
rect 14369 3451 14427 3457
rect 14369 3448 14381 3451
rect 8444 3420 11284 3448
rect 8444 3408 8450 3420
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 3237 3383 3295 3389
rect 3237 3380 3249 3383
rect 2648 3352 3249 3380
rect 2648 3340 2654 3352
rect 3237 3349 3249 3352
rect 3283 3349 3295 3383
rect 3237 3343 3295 3349
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 5626 3380 5632 3392
rect 4120 3352 5632 3380
rect 4120 3340 4126 3352
rect 5626 3340 5632 3352
rect 5684 3340 5690 3392
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8205 3383 8263 3389
rect 8205 3380 8217 3383
rect 8076 3352 8217 3380
rect 8076 3340 8082 3352
rect 8205 3349 8217 3352
rect 8251 3380 8263 3383
rect 11146 3380 11152 3392
rect 8251 3352 11152 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 11146 3340 11152 3352
rect 11204 3340 11210 3392
rect 11256 3389 11284 3420
rect 13556 3420 14381 3448
rect 13556 3389 13584 3420
rect 14369 3417 14381 3420
rect 14415 3417 14427 3451
rect 14826 3448 14832 3460
rect 14787 3420 14832 3448
rect 14369 3411 14427 3417
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 53282 3408 53288 3460
rect 53340 3448 53346 3460
rect 55186 3448 55214 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 57514 3516 57520 3528
rect 57475 3488 57520 3516
rect 55953 3479 56011 3485
rect 57514 3476 57520 3488
rect 57572 3476 57578 3528
rect 58158 3516 58164 3528
rect 58119 3488 58164 3516
rect 58158 3476 58164 3488
rect 58216 3476 58222 3528
rect 53340 3420 55214 3448
rect 53340 3408 53346 3420
rect 11241 3383 11299 3389
rect 11241 3349 11253 3383
rect 11287 3349 11299 3383
rect 11241 3343 11299 3349
rect 13541 3383 13599 3389
rect 13541 3349 13553 3383
rect 13587 3349 13599 3383
rect 14274 3380 14280 3392
rect 14235 3352 14280 3380
rect 13541 3343 13599 3349
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1857 3179 1915 3185
rect 1857 3145 1869 3179
rect 1903 3176 1915 3179
rect 5718 3176 5724 3188
rect 1903 3148 5724 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 7558 3176 7564 3188
rect 5960 3148 7564 3176
rect 5960 3136 5966 3148
rect 7558 3136 7564 3148
rect 7616 3136 7622 3188
rect 7834 3136 7840 3188
rect 7892 3176 7898 3188
rect 12066 3176 12072 3188
rect 7892 3148 12072 3176
rect 7892 3136 7898 3148
rect 3326 3117 3332 3120
rect 3320 3108 3332 3117
rect 3287 3080 3332 3108
rect 3320 3071 3332 3080
rect 3326 3068 3332 3071
rect 3384 3068 3390 3120
rect 5074 3068 5080 3120
rect 5132 3108 5138 3120
rect 7098 3108 7104 3120
rect 5132 3080 7104 3108
rect 5132 3068 5138 3080
rect 7098 3068 7104 3080
rect 7156 3108 7162 3120
rect 7156 3080 7880 3108
rect 7156 3068 7162 3080
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 2590 3040 2596 3052
rect 2551 3012 2596 3040
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 4982 3040 4988 3052
rect 4939 3012 4988 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 4982 3000 4988 3012
rect 5040 3000 5046 3052
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6270 3040 6276 3052
rect 5960 3012 6276 3040
rect 5960 3000 5966 3012
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6822 3000 6828 3052
rect 6880 3040 6886 3052
rect 7653 3043 7711 3049
rect 7653 3040 7665 3043
rect 6880 3012 7665 3040
rect 6880 3000 6886 3012
rect 7653 3009 7665 3012
rect 7699 3040 7711 3043
rect 7742 3040 7748 3052
rect 7699 3012 7748 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 3053 2975 3111 2981
rect 3053 2972 3065 2975
rect 2188 2944 3065 2972
rect 2188 2932 2194 2944
rect 3053 2941 3065 2944
rect 3099 2941 3111 2975
rect 3053 2935 3111 2941
rect 4798 2932 4804 2984
rect 4856 2972 4862 2984
rect 7374 2972 7380 2984
rect 4856 2944 5856 2972
rect 7335 2944 7380 2972
rect 4856 2932 4862 2944
rect 5828 2916 5856 2944
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 5718 2904 5724 2916
rect 4264 2876 5724 2904
rect 2409 2839 2467 2845
rect 2409 2805 2421 2839
rect 2455 2836 2467 2839
rect 4264 2836 4292 2876
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 5810 2864 5816 2916
rect 5868 2864 5874 2916
rect 7852 2904 7880 3080
rect 8754 3068 8760 3120
rect 8812 3108 8818 3120
rect 9398 3108 9404 3120
rect 8812 3080 9404 3108
rect 8812 3068 8818 3080
rect 9398 3068 9404 3080
rect 9456 3108 9462 3120
rect 9585 3111 9643 3117
rect 9585 3108 9597 3111
rect 9456 3080 9597 3108
rect 9456 3068 9462 3080
rect 9585 3077 9597 3080
rect 9631 3077 9643 3111
rect 10410 3108 10416 3120
rect 10371 3080 10416 3108
rect 9585 3071 9643 3077
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 10796 3117 10824 3148
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 12897 3179 12955 3185
rect 12406 3148 12848 3176
rect 10781 3111 10839 3117
rect 10781 3077 10793 3111
rect 10827 3077 10839 3111
rect 10781 3071 10839 3077
rect 10962 3068 10968 3120
rect 11020 3108 11026 3120
rect 12406 3108 12434 3148
rect 11020 3080 12434 3108
rect 12820 3108 12848 3148
rect 12897 3145 12909 3179
rect 12943 3176 12955 3179
rect 14274 3176 14280 3188
rect 12943 3148 14280 3176
rect 12943 3145 12955 3148
rect 12897 3139 12955 3145
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 26234 3108 26240 3120
rect 12820 3080 26240 3108
rect 11020 3068 11026 3080
rect 26234 3068 26240 3080
rect 26292 3068 26298 3120
rect 51902 3068 51908 3120
rect 51960 3108 51966 3120
rect 51960 3080 54708 3108
rect 51960 3068 51966 3080
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8570 3040 8576 3052
rect 8159 3012 8576 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 8570 3000 8576 3012
rect 8628 3000 8634 3052
rect 8846 3040 8852 3052
rect 8680 3012 8852 3040
rect 8680 2981 8708 3012
rect 8846 3000 8852 3012
rect 8904 3000 8910 3052
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9490 3040 9496 3052
rect 9079 3012 9496 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10980 3040 11008 3068
rect 9999 3012 11008 3040
rect 11793 3043 11851 3049
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 11793 3009 11805 3043
rect 11839 3040 11851 3043
rect 12618 3040 12624 3052
rect 11839 3012 12624 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 12618 3000 12624 3012
rect 12676 3000 12682 3052
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 13446 3040 13452 3052
rect 12759 3012 13452 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 13446 3000 13452 3012
rect 13504 3040 13510 3052
rect 14458 3040 14464 3052
rect 13504 3012 14464 3040
rect 13504 3000 13510 3012
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 51718 3000 51724 3052
rect 51776 3040 51782 3052
rect 54680 3049 54708 3080
rect 54021 3043 54079 3049
rect 54021 3040 54033 3043
rect 51776 3012 54033 3040
rect 51776 3000 51782 3012
rect 54021 3009 54033 3012
rect 54067 3009 54079 3043
rect 54021 3003 54079 3009
rect 54665 3043 54723 3049
rect 54665 3009 54677 3043
rect 54711 3009 54723 3043
rect 54665 3003 54723 3009
rect 54754 3000 54760 3052
rect 54812 3040 54818 3052
rect 55309 3043 55367 3049
rect 55309 3040 55321 3043
rect 54812 3012 55321 3040
rect 54812 3000 54818 3012
rect 55309 3009 55321 3012
rect 55355 3009 55367 3043
rect 55309 3003 55367 3009
rect 8665 2975 8723 2981
rect 8665 2941 8677 2975
rect 8711 2941 8723 2975
rect 9122 2972 9128 2984
rect 8665 2935 8723 2941
rect 8772 2944 9128 2972
rect 8481 2907 8539 2913
rect 7852 2876 8156 2904
rect 2455 2808 4292 2836
rect 4433 2839 4491 2845
rect 2455 2805 2467 2808
rect 2409 2799 2467 2805
rect 4433 2805 4445 2839
rect 4479 2836 4491 2839
rect 4706 2836 4712 2848
rect 4479 2808 4712 2836
rect 4479 2805 4491 2808
rect 4433 2799 4491 2805
rect 4706 2796 4712 2808
rect 4764 2836 4770 2848
rect 4982 2836 4988 2848
rect 4764 2808 4988 2836
rect 4764 2796 4770 2808
rect 4982 2796 4988 2808
rect 5040 2796 5046 2848
rect 5074 2796 5080 2848
rect 5132 2836 5138 2848
rect 5629 2839 5687 2845
rect 5132 2808 5177 2836
rect 5132 2796 5138 2808
rect 5629 2805 5641 2839
rect 5675 2836 5687 2839
rect 8018 2836 8024 2848
rect 5675 2808 8024 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8128 2836 8156 2876
rect 8481 2873 8493 2907
rect 8527 2904 8539 2907
rect 8772 2904 8800 2944
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 9306 2932 9312 2984
rect 9364 2972 9370 2984
rect 11698 2972 11704 2984
rect 9364 2944 11704 2972
rect 9364 2932 9370 2944
rect 11698 2932 11704 2944
rect 11756 2972 11762 2984
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 11756 2944 16681 2972
rect 11756 2932 11762 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 18049 2975 18107 2981
rect 18049 2941 18061 2975
rect 18095 2972 18107 2975
rect 18690 2972 18696 2984
rect 18095 2944 18696 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 19978 2972 19984 2984
rect 19383 2944 19984 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 25777 2975 25835 2981
rect 25777 2941 25789 2975
rect 25823 2972 25835 2975
rect 26418 2972 26424 2984
rect 25823 2944 26424 2972
rect 25823 2941 25835 2944
rect 25777 2935 25835 2941
rect 26418 2932 26424 2944
rect 26476 2932 26482 2984
rect 32766 2932 32772 2984
rect 32824 2972 32830 2984
rect 33413 2975 33471 2981
rect 33413 2972 33425 2975
rect 32824 2944 33425 2972
rect 32824 2932 32830 2944
rect 33413 2941 33425 2944
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 38286 2932 38292 2984
rect 38344 2972 38350 2984
rect 39209 2975 39267 2981
rect 39209 2972 39221 2975
rect 38344 2944 39221 2972
rect 38344 2932 38350 2944
rect 39209 2941 39221 2944
rect 39255 2941 39267 2975
rect 39209 2935 39267 2941
rect 42150 2932 42156 2984
rect 42208 2972 42214 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 42208 2944 43085 2972
rect 42208 2932 42214 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 53098 2932 53104 2984
rect 53156 2972 53162 2984
rect 55953 2975 56011 2981
rect 55953 2972 55965 2975
rect 53156 2944 55965 2972
rect 53156 2932 53162 2944
rect 55953 2941 55965 2944
rect 55999 2941 56011 2975
rect 56594 2972 56600 2984
rect 56555 2944 56600 2972
rect 55953 2935 56011 2941
rect 56594 2932 56600 2944
rect 56652 2932 56658 2984
rect 8527 2876 8800 2904
rect 8527 2873 8539 2876
rect 8481 2867 8539 2873
rect 8846 2864 8852 2916
rect 8904 2904 8910 2916
rect 11609 2907 11667 2913
rect 11609 2904 11621 2907
rect 8904 2876 11621 2904
rect 8904 2864 8910 2876
rect 11609 2873 11621 2876
rect 11655 2873 11667 2907
rect 11609 2867 11667 2873
rect 14185 2907 14243 2913
rect 14185 2873 14197 2907
rect 14231 2904 14243 2907
rect 14918 2904 14924 2916
rect 14231 2876 14924 2904
rect 14231 2873 14243 2876
rect 14185 2867 14243 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 33870 2864 33876 2916
rect 33928 2904 33934 2916
rect 34701 2907 34759 2913
rect 34701 2904 34713 2907
rect 33928 2876 34713 2904
rect 33928 2864 33934 2876
rect 34701 2873 34713 2876
rect 34747 2873 34759 2907
rect 34701 2867 34759 2873
rect 37182 2864 37188 2916
rect 37240 2904 37246 2916
rect 37921 2907 37979 2913
rect 37921 2904 37933 2907
rect 37240 2876 37933 2904
rect 37240 2864 37246 2876
rect 37921 2873 37933 2876
rect 37967 2873 37979 2907
rect 37921 2867 37979 2873
rect 39114 2864 39120 2916
rect 39172 2904 39178 2916
rect 39853 2907 39911 2913
rect 39853 2904 39865 2907
rect 39172 2876 39865 2904
rect 39172 2864 39178 2876
rect 39853 2873 39865 2876
rect 39899 2873 39911 2907
rect 39853 2867 39911 2873
rect 40218 2864 40224 2916
rect 40276 2904 40282 2916
rect 41141 2907 41199 2913
rect 41141 2904 41153 2907
rect 40276 2876 41153 2904
rect 40276 2864 40282 2876
rect 41141 2873 41153 2876
rect 41187 2873 41199 2907
rect 41141 2867 41199 2873
rect 42978 2864 42984 2916
rect 43036 2904 43042 2916
rect 43717 2907 43775 2913
rect 43717 2904 43729 2907
rect 43036 2876 43729 2904
rect 43036 2864 43042 2876
rect 43717 2873 43729 2876
rect 43763 2873 43775 2907
rect 43717 2867 43775 2873
rect 44082 2864 44088 2916
rect 44140 2904 44146 2916
rect 45005 2907 45063 2913
rect 45005 2904 45017 2907
rect 44140 2876 45017 2904
rect 44140 2864 44146 2876
rect 45005 2873 45017 2876
rect 45051 2873 45063 2907
rect 45649 2907 45707 2913
rect 45649 2904 45661 2907
rect 45005 2867 45063 2873
rect 45112 2876 45661 2904
rect 8573 2839 8631 2845
rect 8573 2836 8585 2839
rect 8128 2808 8585 2836
rect 8573 2805 8585 2808
rect 8619 2836 8631 2839
rect 8662 2836 8668 2848
rect 8619 2808 8668 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 13541 2839 13599 2845
rect 13541 2805 13553 2839
rect 13587 2836 13599 2839
rect 14642 2836 14648 2848
rect 13587 2808 14648 2836
rect 13587 2805 13599 2808
rect 13541 2799 13599 2805
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15378 2836 15384 2848
rect 14875 2808 15384 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15378 2796 15384 2808
rect 15436 2796 15442 2848
rect 15473 2839 15531 2845
rect 15473 2805 15485 2839
rect 15519 2836 15531 2839
rect 15654 2836 15660 2848
rect 15519 2808 15660 2836
rect 15519 2805 15531 2808
rect 15473 2799 15531 2805
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 16117 2839 16175 2845
rect 16117 2805 16129 2839
rect 16163 2836 16175 2839
rect 16482 2836 16488 2848
rect 16163 2808 16488 2836
rect 16163 2805 16175 2808
rect 16117 2799 16175 2805
rect 16482 2796 16488 2808
rect 16540 2796 16546 2848
rect 17405 2839 17463 2845
rect 17405 2805 17417 2839
rect 17451 2836 17463 2839
rect 17862 2836 17868 2848
rect 17451 2808 17868 2836
rect 17451 2805 17463 2808
rect 17405 2799 17463 2805
rect 17862 2796 17868 2808
rect 17920 2796 17926 2848
rect 18693 2839 18751 2845
rect 18693 2805 18705 2839
rect 18739 2836 18751 2839
rect 19242 2836 19248 2848
rect 18739 2808 19248 2836
rect 18739 2805 18751 2808
rect 18693 2799 18751 2805
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 19981 2839 20039 2845
rect 19981 2805 19993 2839
rect 20027 2836 20039 2839
rect 20530 2836 20536 2848
rect 20027 2808 20536 2836
rect 20027 2805 20039 2808
rect 19981 2799 20039 2805
rect 20530 2796 20536 2808
rect 20588 2796 20594 2848
rect 20625 2839 20683 2845
rect 20625 2805 20637 2839
rect 20671 2836 20683 2839
rect 20898 2836 20904 2848
rect 20671 2808 20904 2836
rect 20671 2805 20683 2808
rect 20625 2799 20683 2805
rect 20898 2796 20904 2808
rect 20956 2796 20962 2848
rect 21269 2839 21327 2845
rect 21269 2805 21281 2839
rect 21315 2836 21327 2839
rect 21726 2836 21732 2848
rect 21315 2808 21732 2836
rect 21315 2805 21327 2808
rect 21269 2799 21327 2805
rect 21726 2796 21732 2808
rect 21784 2796 21790 2848
rect 22557 2839 22615 2845
rect 22557 2805 22569 2839
rect 22603 2836 22615 2839
rect 23106 2836 23112 2848
rect 22603 2808 23112 2836
rect 22603 2805 22615 2808
rect 22557 2799 22615 2805
rect 23106 2796 23112 2808
rect 23164 2796 23170 2848
rect 23201 2839 23259 2845
rect 23201 2805 23213 2839
rect 23247 2836 23259 2839
rect 23658 2836 23664 2848
rect 23247 2808 23664 2836
rect 23247 2805 23259 2808
rect 23201 2799 23259 2805
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2836 23903 2839
rect 24210 2836 24216 2848
rect 23891 2808 24216 2836
rect 23891 2805 23903 2808
rect 23845 2799 23903 2805
rect 24210 2796 24216 2808
rect 24268 2796 24274 2848
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 25038 2836 25044 2848
rect 24535 2808 25044 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2836 25191 2839
rect 25866 2836 25872 2848
rect 25179 2808 25872 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 26970 2836 26976 2848
rect 26467 2808 26976 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 26970 2796 26976 2808
rect 27028 2796 27034 2848
rect 27617 2839 27675 2845
rect 27617 2805 27629 2839
rect 27663 2836 27675 2839
rect 27798 2836 27804 2848
rect 27663 2808 27804 2836
rect 27663 2805 27675 2808
rect 27617 2799 27675 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28074 2836 28080 2848
rect 28035 2808 28080 2836
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 28905 2839 28963 2845
rect 28905 2805 28917 2839
rect 28951 2836 28963 2839
rect 29178 2836 29184 2848
rect 28951 2808 29184 2836
rect 28951 2805 28963 2808
rect 28905 2799 28963 2805
rect 29178 2796 29184 2808
rect 29236 2796 29242 2848
rect 29549 2839 29607 2845
rect 29549 2805 29561 2839
rect 29595 2836 29607 2839
rect 29730 2836 29736 2848
rect 29595 2808 29736 2836
rect 29595 2805 29607 2808
rect 29549 2799 29607 2805
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 30006 2836 30012 2848
rect 29967 2808 30012 2836
rect 30006 2796 30012 2808
rect 30064 2796 30070 2848
rect 30558 2796 30564 2848
rect 30616 2836 30622 2848
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 30616 2808 30665 2836
rect 30616 2796 30622 2808
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 31662 2796 31668 2848
rect 31720 2836 31726 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31720 2808 32137 2836
rect 31720 2796 31726 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 32769 2839 32827 2845
rect 32769 2836 32781 2839
rect 32272 2808 32781 2836
rect 32272 2796 32278 2808
rect 32769 2805 32781 2808
rect 32815 2805 32827 2839
rect 32769 2799 32827 2805
rect 33318 2796 33324 2848
rect 33376 2836 33382 2848
rect 34057 2839 34115 2845
rect 34057 2836 34069 2839
rect 33376 2808 34069 2836
rect 33376 2796 33382 2808
rect 34057 2805 34069 2808
rect 34103 2805 34115 2839
rect 34057 2799 34115 2805
rect 34422 2796 34428 2848
rect 34480 2836 34486 2848
rect 35345 2839 35403 2845
rect 35345 2836 35357 2839
rect 34480 2808 35357 2836
rect 34480 2796 34486 2808
rect 35345 2805 35357 2808
rect 35391 2805 35403 2839
rect 35345 2799 35403 2805
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35989 2839 36047 2845
rect 35989 2836 36001 2839
rect 35492 2808 36001 2836
rect 35492 2796 35498 2808
rect 35989 2805 36001 2808
rect 36035 2805 36047 2839
rect 35989 2799 36047 2805
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36412 2808 37289 2836
rect 36412 2796 36418 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37734 2796 37740 2848
rect 37792 2836 37798 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 37792 2808 38577 2836
rect 37792 2796 37798 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 39666 2796 39672 2848
rect 39724 2836 39730 2848
rect 40497 2839 40555 2845
rect 40497 2836 40509 2839
rect 39724 2808 40509 2836
rect 39724 2796 39730 2808
rect 40497 2805 40509 2808
rect 40543 2805 40555 2839
rect 40497 2799 40555 2805
rect 41598 2796 41604 2848
rect 41656 2836 41662 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41656 2808 42441 2836
rect 41656 2796 41662 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 43530 2796 43536 2848
rect 43588 2836 43594 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 43588 2808 44373 2836
rect 43588 2796 43594 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 44910 2796 44916 2848
rect 44968 2836 44974 2848
rect 45112 2836 45140 2876
rect 45649 2873 45661 2876
rect 45695 2873 45707 2907
rect 45649 2867 45707 2873
rect 47394 2864 47400 2916
rect 47452 2904 47458 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 47452 2876 48237 2904
rect 47452 2864 47458 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 48774 2864 48780 2916
rect 48832 2904 48838 2916
rect 49513 2907 49571 2913
rect 49513 2904 49525 2907
rect 48832 2876 49525 2904
rect 48832 2864 48838 2876
rect 49513 2873 49525 2876
rect 49559 2873 49571 2907
rect 49513 2867 49571 2873
rect 49878 2864 49884 2916
rect 49936 2904 49942 2916
rect 50801 2907 50859 2913
rect 50801 2904 50813 2907
rect 49936 2876 50813 2904
rect 49936 2864 49942 2876
rect 50801 2873 50813 2876
rect 50847 2873 50859 2907
rect 50801 2867 50859 2873
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 52733 2907 52791 2913
rect 52733 2904 52745 2907
rect 51040 2876 52745 2904
rect 51040 2864 51046 2876
rect 52733 2873 52745 2876
rect 52779 2873 52791 2907
rect 52733 2867 52791 2873
rect 54202 2864 54208 2916
rect 54260 2904 54266 2916
rect 57885 2907 57943 2913
rect 57885 2904 57897 2907
rect 54260 2876 57897 2904
rect 54260 2864 54266 2876
rect 57885 2873 57897 2876
rect 57931 2873 57943 2907
rect 57885 2867 57943 2873
rect 44968 2808 45140 2836
rect 44968 2796 44974 2808
rect 45462 2796 45468 2848
rect 45520 2836 45526 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45520 2808 46305 2836
rect 45520 2796 45526 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 46842 2796 46848 2848
rect 46900 2836 46906 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46900 2808 47593 2836
rect 46900 2796 46906 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 47946 2796 47952 2848
rect 48004 2836 48010 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48004 2808 48881 2836
rect 48004 2796 48010 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49326 2796 49332 2848
rect 49384 2836 49390 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49384 2808 50169 2836
rect 49384 2796 49390 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 50706 2796 50712 2848
rect 50764 2836 50770 2848
rect 51445 2839 51503 2845
rect 51445 2836 51457 2839
rect 50764 2808 51457 2836
rect 50764 2796 50770 2808
rect 51445 2805 51457 2808
rect 51491 2805 51503 2839
rect 51445 2799 51503 2805
rect 51534 2796 51540 2848
rect 51592 2836 51598 2848
rect 53377 2839 53435 2845
rect 53377 2836 53389 2839
rect 51592 2808 53389 2836
rect 51592 2796 51598 2808
rect 53377 2805 53389 2808
rect 53423 2805 53435 2839
rect 53377 2799 53435 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 2774 2632 2780 2644
rect 1811 2604 2780 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 5583 2635 5641 2641
rect 5583 2601 5595 2635
rect 5629 2632 5641 2635
rect 5902 2632 5908 2644
rect 5629 2604 5908 2632
rect 5629 2601 5641 2604
rect 5583 2595 5641 2601
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 6638 2632 6644 2644
rect 6599 2604 6644 2632
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 12437 2635 12495 2641
rect 12437 2632 12449 2635
rect 8628 2604 12449 2632
rect 8628 2592 8634 2604
rect 12437 2601 12449 2604
rect 12483 2601 12495 2635
rect 12437 2595 12495 2601
rect 13541 2635 13599 2641
rect 13541 2601 13553 2635
rect 13587 2632 13599 2635
rect 13906 2632 13912 2644
rect 13587 2604 13912 2632
rect 13587 2601 13599 2604
rect 13541 2595 13599 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 19981 2635 20039 2641
rect 14016 2604 16574 2632
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 5258 2564 5264 2576
rect 2363 2536 5264 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 6656 2564 6684 2592
rect 9398 2564 9404 2576
rect 5368 2536 6040 2564
rect 6656 2536 9404 2564
rect 3786 2456 3792 2508
rect 3844 2496 3850 2508
rect 3844 2468 4844 2496
rect 3844 2456 3850 2468
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2280 2400 2513 2428
rect 2280 2388 2286 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2866 2388 2872 2440
rect 2924 2428 2930 2440
rect 2961 2431 3019 2437
rect 2961 2428 2973 2431
rect 2924 2400 2973 2428
rect 2924 2388 2930 2400
rect 2961 2397 2973 2400
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4525 2431 4583 2437
rect 4525 2428 4537 2431
rect 4120 2400 4537 2428
rect 4120 2388 4126 2400
rect 4525 2397 4537 2400
rect 4571 2397 4583 2431
rect 4816 2428 4844 2468
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 5368 2496 5396 2536
rect 5040 2468 5396 2496
rect 6012 2496 6040 2536
rect 9398 2524 9404 2536
rect 9456 2524 9462 2576
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 10781 2567 10839 2573
rect 10781 2564 10793 2567
rect 9732 2536 10793 2564
rect 9732 2524 9738 2536
rect 10781 2533 10793 2536
rect 10827 2533 10839 2567
rect 10781 2527 10839 2533
rect 11514 2524 11520 2576
rect 11572 2564 11578 2576
rect 11609 2567 11667 2573
rect 11609 2564 11621 2567
rect 11572 2536 11621 2564
rect 11572 2524 11578 2536
rect 11609 2533 11621 2536
rect 11655 2533 11667 2567
rect 11609 2527 11667 2533
rect 6012 2468 7420 2496
rect 5040 2456 5046 2468
rect 5626 2428 5632 2440
rect 4816 2400 5632 2428
rect 4525 2391 4583 2397
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6086 2428 6092 2440
rect 5859 2400 6092 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7248 2400 7297 2428
rect 7248 2388 7254 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7392 2428 7420 2468
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 7561 2499 7619 2505
rect 7561 2496 7573 2499
rect 7524 2468 7573 2496
rect 7524 2456 7530 2468
rect 7561 2465 7573 2468
rect 7607 2465 7619 2499
rect 7561 2459 7619 2465
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 14016 2496 14044 2604
rect 14829 2567 14887 2573
rect 14829 2533 14841 2567
rect 14875 2564 14887 2567
rect 16206 2564 16212 2576
rect 14875 2536 16212 2564
rect 14875 2533 14887 2536
rect 14829 2527 14887 2533
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 16546 2564 16574 2604
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 21450 2632 21456 2644
rect 20027 2604 21456 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 51994 2592 52000 2644
rect 52052 2632 52058 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 52052 2604 55321 2632
rect 52052 2592 52058 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 27430 2564 27436 2576
rect 16546 2536 27436 2564
rect 27430 2524 27436 2536
rect 27488 2524 27494 2576
rect 27709 2567 27767 2573
rect 27709 2533 27721 2567
rect 27755 2564 27767 2567
rect 28350 2564 28356 2576
rect 27755 2536 28356 2564
rect 27755 2533 27767 2536
rect 27709 2527 27767 2533
rect 28350 2524 28356 2536
rect 28408 2524 28414 2576
rect 34146 2524 34152 2576
rect 34204 2564 34210 2576
rect 35989 2567 36047 2573
rect 35989 2564 36001 2567
rect 34204 2536 36001 2564
rect 34204 2524 34210 2536
rect 35989 2533 36001 2536
rect 36035 2533 36047 2567
rect 35989 2527 36047 2533
rect 38010 2524 38016 2576
rect 38068 2564 38074 2576
rect 39853 2567 39911 2573
rect 39853 2564 39865 2567
rect 38068 2536 39865 2564
rect 38068 2524 38074 2536
rect 39853 2533 39865 2536
rect 39899 2533 39911 2567
rect 39853 2527 39911 2533
rect 41874 2524 41880 2576
rect 41932 2564 41938 2576
rect 43717 2567 43775 2573
rect 43717 2564 43729 2567
rect 41932 2536 43729 2564
rect 41932 2524 41938 2536
rect 43717 2533 43729 2536
rect 43763 2533 43775 2567
rect 43717 2527 43775 2533
rect 45738 2524 45744 2576
rect 45796 2564 45802 2576
rect 47581 2567 47639 2573
rect 47581 2564 47593 2567
rect 45796 2536 47593 2564
rect 45796 2524 45802 2536
rect 47581 2533 47593 2536
rect 47627 2533 47639 2567
rect 47581 2527 47639 2533
rect 49602 2524 49608 2576
rect 49660 2564 49666 2576
rect 51445 2567 51503 2573
rect 51445 2564 51457 2567
rect 49660 2536 51457 2564
rect 49660 2524 49666 2536
rect 51445 2533 51457 2536
rect 51491 2533 51503 2567
rect 51445 2527 51503 2533
rect 54021 2567 54079 2573
rect 54021 2533 54033 2567
rect 54067 2533 54079 2567
rect 54021 2527 54079 2533
rect 9548 2468 10640 2496
rect 9548 2456 9554 2468
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 7392 2400 8953 2428
rect 7285 2391 7343 2397
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9398 2388 9404 2440
rect 9456 2428 9462 2440
rect 10612 2437 10640 2468
rect 12406 2468 14044 2496
rect 15473 2499 15531 2505
rect 10597 2431 10655 2437
rect 9456 2400 9904 2428
rect 9456 2388 9462 2400
rect 6733 2363 6791 2369
rect 3160 2332 6684 2360
rect 3160 2301 3188 2332
rect 3145 2295 3203 2301
rect 3145 2261 3157 2295
rect 3191 2261 3203 2295
rect 3145 2255 3203 2261
rect 4341 2295 4399 2301
rect 4341 2261 4353 2295
rect 4387 2292 4399 2295
rect 5902 2292 5908 2304
rect 4387 2264 5908 2292
rect 4387 2261 4399 2264
rect 4341 2255 4399 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 6656 2292 6684 2332
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 7926 2360 7932 2372
rect 6779 2332 7932 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 7926 2320 7932 2332
rect 7984 2320 7990 2372
rect 8202 2320 8208 2372
rect 8260 2360 8266 2372
rect 9490 2360 9496 2372
rect 8260 2332 9496 2360
rect 8260 2320 8266 2332
rect 9490 2320 9496 2332
rect 9548 2320 9554 2372
rect 9582 2320 9588 2372
rect 9640 2360 9646 2372
rect 9769 2363 9827 2369
rect 9769 2360 9781 2363
rect 9640 2332 9781 2360
rect 9640 2320 9646 2332
rect 9769 2329 9781 2332
rect 9815 2329 9827 2363
rect 9876 2360 9904 2400
rect 10597 2397 10609 2431
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 11793 2431 11851 2437
rect 11793 2428 11805 2431
rect 11756 2400 11805 2428
rect 11756 2388 11762 2400
rect 11793 2397 11805 2400
rect 11839 2397 11851 2431
rect 12250 2428 12256 2440
rect 12211 2400 12256 2428
rect 11793 2391 11851 2397
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 12406 2360 12434 2468
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 17034 2496 17040 2508
rect 15519 2468 17040 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 17405 2499 17463 2505
rect 17405 2465 17417 2499
rect 17451 2496 17463 2499
rect 18138 2496 18144 2508
rect 17451 2468 18144 2496
rect 17451 2465 17463 2468
rect 17405 2459 17463 2465
rect 18138 2456 18144 2468
rect 18196 2456 18202 2508
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2496 18751 2499
rect 20070 2496 20076 2508
rect 18739 2468 20076 2496
rect 18739 2465 18751 2468
rect 18693 2459 18751 2465
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 22002 2496 22008 2508
rect 20671 2468 22008 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 23845 2499 23903 2505
rect 23845 2465 23857 2499
rect 23891 2496 23903 2499
rect 25314 2496 25320 2508
rect 23891 2468 25320 2496
rect 23891 2465 23903 2468
rect 23845 2459 23903 2465
rect 25314 2456 25320 2468
rect 25372 2456 25378 2508
rect 25777 2499 25835 2505
rect 25777 2465 25789 2499
rect 25823 2496 25835 2499
rect 26694 2496 26700 2508
rect 25823 2468 26700 2496
rect 25823 2465 25835 2468
rect 25777 2459 25835 2465
rect 26694 2456 26700 2468
rect 26752 2456 26758 2508
rect 31938 2456 31944 2508
rect 31996 2496 32002 2508
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 31996 2468 32781 2496
rect 31996 2456 32002 2468
rect 32769 2465 32781 2468
rect 32815 2465 32827 2499
rect 32769 2459 32827 2465
rect 33042 2456 33048 2508
rect 33100 2496 33106 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 33100 2468 34713 2496
rect 33100 2456 33106 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 35526 2456 35532 2508
rect 35584 2496 35590 2508
rect 37277 2499 37335 2505
rect 37277 2496 37289 2499
rect 35584 2468 37289 2496
rect 35584 2456 35590 2468
rect 37277 2465 37289 2468
rect 37323 2465 37335 2499
rect 37277 2459 37335 2465
rect 38838 2456 38844 2508
rect 38896 2496 38902 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 38896 2468 40509 2496
rect 38896 2456 38902 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 40770 2456 40776 2508
rect 40828 2496 40834 2508
rect 42429 2499 42487 2505
rect 42429 2496 42441 2499
rect 40828 2468 42441 2496
rect 40828 2456 40834 2468
rect 42429 2465 42441 2468
rect 42475 2465 42487 2499
rect 42429 2459 42487 2465
rect 43254 2456 43260 2508
rect 43312 2496 43318 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 43312 2468 45017 2496
rect 43312 2456 43318 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45005 2459 45063 2465
rect 46566 2456 46572 2508
rect 46624 2496 46630 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 46624 2468 48237 2496
rect 46624 2456 46630 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 48498 2456 48504 2508
rect 48556 2496 48562 2508
rect 50157 2499 50215 2505
rect 50157 2496 50169 2499
rect 48556 2468 50169 2496
rect 48556 2456 48562 2468
rect 50157 2465 50169 2468
rect 50203 2465 50215 2499
rect 52733 2499 52791 2505
rect 52733 2496 52745 2499
rect 50157 2459 50215 2465
rect 51046 2468 52745 2496
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 17310 2428 17316 2440
rect 16163 2400 17316 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 9876 2332 12434 2360
rect 13372 2360 13400 2391
rect 17310 2388 17316 2400
rect 17368 2388 17374 2440
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2428 22615 2431
rect 23201 2431 23259 2437
rect 22603 2400 23152 2428
rect 22603 2397 22615 2400
rect 22557 2391 22615 2397
rect 15010 2360 15016 2372
rect 13372 2332 15016 2360
rect 9769 2323 9827 2329
rect 15010 2320 15016 2332
rect 15068 2360 15074 2372
rect 18064 2360 18092 2391
rect 18966 2360 18972 2372
rect 15068 2332 16574 2360
rect 18064 2332 18972 2360
rect 15068 2320 15074 2332
rect 7374 2292 7380 2304
rect 6656 2264 7380 2292
rect 7374 2252 7380 2264
rect 7432 2252 7438 2304
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 9398 2292 9404 2304
rect 9171 2264 9404 2292
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 9858 2292 9864 2304
rect 9819 2264 9864 2292
rect 9858 2252 9864 2264
rect 9916 2252 9922 2304
rect 14182 2292 14188 2304
rect 14143 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 16546 2292 16574 2332
rect 18966 2320 18972 2332
rect 19024 2320 19030 2372
rect 21284 2360 21312 2391
rect 22830 2360 22836 2372
rect 21284 2332 22836 2360
rect 22830 2320 22836 2332
rect 22888 2320 22894 2372
rect 23124 2360 23152 2400
rect 23201 2397 23213 2431
rect 23247 2428 23259 2431
rect 24762 2428 24768 2440
rect 23247 2400 24768 2428
rect 23247 2397 23259 2400
rect 23201 2391 23259 2397
rect 24762 2388 24768 2400
rect 24820 2388 24826 2440
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2428 25191 2431
rect 26142 2428 26148 2440
rect 25179 2400 26148 2428
rect 25179 2397 25191 2400
rect 25133 2391 25191 2397
rect 26142 2388 26148 2400
rect 26200 2388 26206 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 27246 2428 27252 2440
rect 26467 2400 27252 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 27246 2388 27252 2400
rect 27304 2388 27310 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28902 2428 28908 2440
rect 28399 2400 28908 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28902 2388 28908 2400
rect 28960 2388 28966 2440
rect 28997 2431 29055 2437
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 29454 2428 29460 2440
rect 29043 2400 29460 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29454 2388 29460 2400
rect 29512 2388 29518 2440
rect 30101 2431 30159 2437
rect 30101 2397 30113 2431
rect 30147 2428 30159 2431
rect 30282 2428 30288 2440
rect 30147 2400 30288 2428
rect 30147 2397 30159 2400
rect 30101 2391 30159 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2428 30803 2431
rect 30834 2428 30840 2440
rect 30791 2400 30840 2428
rect 30791 2397 30803 2400
rect 30745 2391 30803 2397
rect 30834 2388 30840 2400
rect 30892 2388 30898 2440
rect 31110 2388 31116 2440
rect 31168 2428 31174 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 31168 2400 31217 2428
rect 31168 2388 31174 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31444 2400 32137 2428
rect 31444 2388 31450 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32490 2388 32496 2440
rect 32548 2428 32554 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 32548 2400 33425 2428
rect 32548 2388 32554 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 33594 2388 33600 2440
rect 33652 2428 33658 2440
rect 35345 2431 35403 2437
rect 35345 2428 35357 2431
rect 33652 2400 35357 2428
rect 33652 2388 33658 2400
rect 35345 2397 35357 2400
rect 35391 2397 35403 2431
rect 35345 2391 35403 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37921 2431 37979 2437
rect 37921 2428 37933 2431
rect 36136 2400 37933 2428
rect 36136 2388 36142 2400
rect 37921 2397 37933 2400
rect 37967 2397 37979 2431
rect 37921 2391 37979 2397
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 23934 2360 23940 2372
rect 23124 2332 23940 2360
rect 23934 2320 23940 2332
rect 23992 2320 23998 2372
rect 36906 2320 36912 2372
rect 36964 2360 36970 2372
rect 38580 2360 38608 2391
rect 39390 2388 39396 2440
rect 39448 2428 39454 2440
rect 41141 2431 41199 2437
rect 41141 2428 41153 2431
rect 39448 2400 41153 2428
rect 39448 2388 39454 2400
rect 41141 2397 41153 2400
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 41322 2388 41328 2440
rect 41380 2428 41386 2440
rect 43073 2431 43131 2437
rect 43073 2428 43085 2431
rect 41380 2400 43085 2428
rect 41380 2388 41386 2400
rect 43073 2397 43085 2400
rect 43119 2397 43131 2431
rect 43073 2391 43131 2397
rect 43806 2388 43812 2440
rect 43864 2428 43870 2440
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 43864 2400 45661 2428
rect 43864 2388 43870 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 46293 2431 46351 2437
rect 46293 2397 46305 2431
rect 46339 2397 46351 2431
rect 46293 2391 46351 2397
rect 36964 2332 38608 2360
rect 36964 2320 36970 2332
rect 44634 2320 44640 2372
rect 44692 2360 44698 2372
rect 46308 2360 46336 2391
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 48869 2431 48927 2437
rect 48869 2428 48881 2431
rect 47176 2400 48881 2428
rect 47176 2388 47182 2400
rect 48869 2397 48881 2400
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 49050 2388 49056 2440
rect 49108 2428 49114 2440
rect 50801 2431 50859 2437
rect 50801 2428 50813 2431
rect 49108 2400 50813 2428
rect 49108 2388 49114 2400
rect 50801 2397 50813 2400
rect 50847 2397 50859 2431
rect 50801 2391 50859 2397
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 51046 2428 51074 2468
rect 52733 2465 52745 2468
rect 52779 2465 52791 2499
rect 54036 2496 54064 2527
rect 57882 2496 57888 2508
rect 54036 2468 54156 2496
rect 57843 2468 57888 2496
rect 52733 2459 52791 2465
rect 50948 2400 51074 2428
rect 50948 2388 50954 2400
rect 52546 2388 52552 2440
rect 52604 2428 52610 2440
rect 53377 2431 53435 2437
rect 53377 2428 53389 2431
rect 52604 2400 53389 2428
rect 52604 2388 52610 2400
rect 53377 2397 53389 2400
rect 53423 2397 53435 2431
rect 53377 2391 53435 2397
rect 44692 2332 46336 2360
rect 44692 2320 44698 2332
rect 16669 2295 16727 2301
rect 16669 2292 16681 2295
rect 16546 2264 16681 2292
rect 16669 2261 16681 2264
rect 16715 2261 16727 2295
rect 16669 2255 16727 2261
rect 51258 2252 51264 2304
rect 51316 2292 51322 2304
rect 54128 2292 54156 2468
rect 57882 2456 57888 2468
rect 57940 2456 57946 2508
rect 55950 2428 55956 2440
rect 55911 2400 55956 2428
rect 55950 2388 55956 2400
rect 56008 2388 56014 2440
rect 56594 2428 56600 2440
rect 56555 2400 56600 2428
rect 56594 2388 56600 2400
rect 56652 2388 56658 2440
rect 51316 2264 54156 2292
rect 51316 2252 51322 2264
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 5258 2048 5264 2100
rect 5316 2088 5322 2100
rect 6638 2088 6644 2100
rect 5316 2060 6644 2088
rect 5316 2048 5322 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 52362 2048 52368 2100
rect 52420 2088 52426 2100
rect 55950 2088 55956 2100
rect 52420 2060 55956 2088
rect 52420 2048 52426 2060
rect 55950 2048 55956 2060
rect 56008 2048 56014 2100
rect 11514 1980 11520 2032
rect 11572 2020 11578 2032
rect 17218 2020 17224 2032
rect 11572 1992 17224 2020
rect 11572 1980 11578 1992
rect 17218 1980 17224 1992
rect 17276 1980 17282 2032
rect 53558 1980 53564 2032
rect 53616 2020 53622 2032
rect 57882 2020 57888 2032
rect 53616 1992 57888 2020
rect 53616 1980 53622 1992
rect 57882 1980 57888 1992
rect 57940 1980 57946 2032
rect 12342 1912 12348 1964
rect 12400 1952 12406 1964
rect 20162 1952 20168 1964
rect 12400 1924 20168 1952
rect 12400 1912 12406 1924
rect 20162 1912 20168 1924
rect 20220 1912 20226 1964
rect 1578 1844 1584 1896
rect 1636 1884 1642 1896
rect 7466 1884 7472 1896
rect 1636 1856 7472 1884
rect 1636 1844 1642 1856
rect 7466 1844 7472 1856
rect 7524 1844 7530 1896
rect 7926 1708 7932 1760
rect 7984 1748 7990 1760
rect 8202 1748 8208 1760
rect 7984 1720 8208 1748
rect 7984 1708 7990 1720
rect 8202 1708 8208 1720
rect 8260 1708 8266 1760
rect 5902 1504 5908 1556
rect 5960 1544 5966 1556
rect 7742 1544 7748 1556
rect 5960 1516 7748 1544
rect 5960 1504 5966 1516
rect 7742 1504 7748 1516
rect 7800 1504 7806 1556
rect 3050 1368 3056 1420
rect 3108 1408 3114 1420
rect 5902 1408 5908 1420
rect 3108 1380 5908 1408
rect 3108 1368 3114 1380
rect 5902 1368 5908 1380
rect 5960 1368 5966 1420
rect 7466 1368 7472 1420
rect 7524 1408 7530 1420
rect 7524 1380 7880 1408
rect 7524 1368 7530 1380
rect 7852 1352 7880 1380
rect 52730 1368 52736 1420
rect 52788 1408 52794 1420
rect 53006 1408 53012 1420
rect 52788 1380 53012 1408
rect 52788 1368 52794 1380
rect 53006 1368 53012 1380
rect 53064 1368 53070 1420
rect 56594 1408 56600 1420
rect 53116 1380 56600 1408
rect 5350 1300 5356 1352
rect 5408 1340 5414 1352
rect 5994 1340 6000 1352
rect 5408 1312 6000 1340
rect 5408 1300 5414 1312
rect 5994 1300 6000 1312
rect 6052 1300 6058 1352
rect 7834 1300 7840 1352
rect 7892 1300 7898 1352
rect 52546 1136 52552 1148
rect 51000 1108 52552 1136
rect 51000 944 51028 1108
rect 52546 1096 52552 1108
rect 52604 1096 52610 1148
rect 50982 892 50988 944
rect 51040 892 51046 944
rect 52546 892 52552 944
rect 52604 892 52610 944
rect 52914 892 52920 944
rect 52972 932 52978 944
rect 53116 932 53144 1380
rect 56594 1368 56600 1380
rect 56652 1368 56658 1420
rect 52972 904 53144 932
rect 52972 892 52978 904
rect 52564 864 52592 892
rect 54754 864 54760 876
rect 52564 836 54760 864
rect 54754 824 54760 836
rect 54812 824 54818 876
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 1768 57400 1820 57452
rect 3332 57400 3384 57452
rect 4896 57400 4948 57452
rect 6460 57400 6512 57452
rect 8024 57400 8076 57452
rect 9680 57443 9732 57452
rect 9680 57409 9689 57443
rect 9689 57409 9723 57443
rect 9723 57409 9732 57443
rect 9680 57400 9732 57409
rect 11152 57400 11204 57452
rect 12716 57400 12768 57452
rect 14280 57400 14332 57452
rect 15844 57400 15896 57452
rect 17408 57400 17460 57452
rect 18972 57400 19024 57452
rect 20536 57400 20588 57452
rect 22100 57400 22152 57452
rect 23664 57400 23716 57452
rect 25228 57400 25280 57452
rect 26792 57400 26844 57452
rect 28356 57400 28408 57452
rect 29920 57400 29972 57452
rect 31484 57400 31536 57452
rect 33140 57443 33192 57452
rect 33140 57409 33149 57443
rect 33149 57409 33183 57443
rect 33183 57409 33192 57443
rect 33140 57400 33192 57409
rect 34612 57400 34664 57452
rect 36176 57400 36228 57452
rect 37740 57400 37792 57452
rect 39304 57400 39356 57452
rect 40868 57400 40920 57452
rect 42432 57400 42484 57452
rect 43996 57400 44048 57452
rect 45560 57400 45612 57452
rect 47124 57400 47176 57452
rect 48688 57400 48740 57452
rect 50160 57400 50212 57452
rect 51816 57400 51868 57452
rect 53380 57400 53432 57452
rect 56600 57443 56652 57452
rect 56600 57409 56609 57443
rect 56609 57409 56643 57443
rect 56643 57409 56652 57443
rect 56600 57400 56652 57409
rect 58072 57400 58124 57452
rect 54944 57332 54996 57384
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 57520 57035 57572 57044
rect 57520 57001 57529 57035
rect 57529 57001 57563 57035
rect 57563 57001 57572 57035
rect 57520 56992 57572 57001
rect 57888 56788 57940 56840
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 58440 56312 58492 56364
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 58164 55131 58216 55140
rect 58164 55097 58173 55131
rect 58173 55097 58207 55131
rect 58207 55097 58216 55131
rect 58164 55088 58216 55097
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 57888 53932 57940 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 57888 52436 57940 52488
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 58164 51391 58216 51400
rect 58164 51357 58173 51391
rect 58173 51357 58207 51391
rect 58207 51357 58216 51391
rect 58164 51348 58216 51357
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 58164 49759 58216 49768
rect 58164 49725 58173 49759
rect 58173 49725 58207 49759
rect 58207 49725 58216 49759
rect 58164 49716 58216 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 58164 48535 58216 48544
rect 58164 48501 58173 48535
rect 58173 48501 58207 48535
rect 58207 48501 58216 48535
rect 58164 48492 58216 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 58164 47039 58216 47048
rect 58164 47005 58173 47039
rect 58173 47005 58207 47039
rect 58207 47005 58216 47039
rect 58164 46996 58216 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 58164 45951 58216 45960
rect 58164 45917 58173 45951
rect 58173 45917 58207 45951
rect 58207 45917 58216 45951
rect 58164 45908 58216 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 58164 44251 58216 44260
rect 58164 44217 58173 44251
rect 58173 44217 58207 44251
rect 58207 44217 58216 44251
rect 58164 44208 58216 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 58164 43095 58216 43104
rect 58164 43061 58173 43095
rect 58173 43061 58207 43095
rect 58207 43061 58216 43095
rect 58164 43052 58216 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 12716 42644 12768 42696
rect 20444 42644 20496 42696
rect 14648 42576 14700 42628
rect 16304 42576 16356 42628
rect 14924 42551 14976 42560
rect 14924 42517 14933 42551
rect 14933 42517 14967 42551
rect 14967 42517 14976 42551
rect 14924 42508 14976 42517
rect 15936 42508 15988 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 12164 42304 12216 42356
rect 14648 42279 14700 42288
rect 14648 42245 14657 42279
rect 14657 42245 14691 42279
rect 14691 42245 14700 42279
rect 14648 42236 14700 42245
rect 12716 42211 12768 42220
rect 12716 42177 12725 42211
rect 12725 42177 12759 42211
rect 12759 42177 12768 42211
rect 12716 42168 12768 42177
rect 12900 42211 12952 42220
rect 12900 42177 12914 42211
rect 12914 42177 12948 42211
rect 12948 42177 12952 42211
rect 12900 42168 12952 42177
rect 12716 42032 12768 42084
rect 12992 42032 13044 42084
rect 13912 42168 13964 42220
rect 15384 42168 15436 42220
rect 15476 42211 15528 42220
rect 15476 42177 15485 42211
rect 15485 42177 15519 42211
rect 15519 42177 15528 42211
rect 15476 42168 15528 42177
rect 15752 42211 15804 42220
rect 15752 42177 15761 42211
rect 15761 42177 15795 42211
rect 15795 42177 15804 42211
rect 15752 42168 15804 42177
rect 15476 42032 15528 42084
rect 12072 41964 12124 42016
rect 12440 42007 12492 42016
rect 12440 41973 12449 42007
rect 12449 41973 12483 42007
rect 12483 41973 12492 42007
rect 12440 41964 12492 41973
rect 14556 41964 14608 42016
rect 16120 42007 16172 42016
rect 16120 41973 16129 42007
rect 16129 41973 16163 42007
rect 16163 41973 16172 42007
rect 16120 41964 16172 41973
rect 19892 42100 19944 42152
rect 19524 41964 19576 42016
rect 24768 41964 24820 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 12900 41760 12952 41812
rect 15384 41760 15436 41812
rect 12716 41624 12768 41676
rect 12072 41599 12124 41608
rect 12072 41565 12081 41599
rect 12081 41565 12115 41599
rect 12115 41565 12124 41599
rect 12072 41556 12124 41565
rect 12992 41556 13044 41608
rect 15752 41624 15804 41676
rect 11244 41531 11296 41540
rect 11244 41497 11253 41531
rect 11253 41497 11287 41531
rect 11287 41497 11296 41531
rect 11244 41488 11296 41497
rect 11428 41531 11480 41540
rect 11428 41497 11437 41531
rect 11437 41497 11471 41531
rect 11471 41497 11480 41531
rect 11428 41488 11480 41497
rect 14556 41599 14608 41608
rect 14556 41565 14565 41599
rect 14565 41565 14599 41599
rect 14599 41565 14608 41599
rect 14556 41556 14608 41565
rect 15476 41556 15528 41608
rect 16120 41556 16172 41608
rect 16856 41599 16908 41608
rect 16856 41565 16865 41599
rect 16865 41565 16899 41599
rect 16899 41565 16908 41599
rect 16856 41556 16908 41565
rect 14924 41488 14976 41540
rect 20352 41760 20404 41812
rect 18696 41556 18748 41608
rect 19524 41599 19576 41608
rect 19524 41565 19533 41599
rect 19533 41565 19567 41599
rect 19567 41565 19576 41599
rect 19524 41556 19576 41565
rect 19892 41599 19944 41608
rect 18972 41488 19024 41540
rect 19340 41488 19392 41540
rect 19892 41565 19901 41599
rect 19901 41565 19935 41599
rect 19935 41565 19944 41599
rect 19892 41556 19944 41565
rect 58164 41599 58216 41608
rect 58164 41565 58173 41599
rect 58173 41565 58207 41599
rect 58207 41565 58216 41599
rect 58164 41556 58216 41565
rect 5172 41463 5224 41472
rect 5172 41429 5181 41463
rect 5181 41429 5215 41463
rect 5215 41429 5224 41463
rect 5172 41420 5224 41429
rect 14096 41463 14148 41472
rect 14096 41429 14105 41463
rect 14105 41429 14139 41463
rect 14139 41429 14148 41463
rect 14096 41420 14148 41429
rect 17960 41420 18012 41472
rect 19432 41420 19484 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 6368 41148 6420 41200
rect 12532 41216 12584 41268
rect 15752 41216 15804 41268
rect 11244 41148 11296 41200
rect 12164 41148 12216 41200
rect 12440 41148 12492 41200
rect 14096 41148 14148 41200
rect 6000 41080 6052 41132
rect 4620 40876 4672 40928
rect 9312 41123 9364 41132
rect 9312 41089 9321 41123
rect 9321 41089 9355 41123
rect 9355 41089 9364 41123
rect 9312 41080 9364 41089
rect 10140 41080 10192 41132
rect 14924 41080 14976 41132
rect 9956 41012 10008 41064
rect 12900 41055 12952 41064
rect 12900 41021 12909 41055
rect 12909 41021 12943 41055
rect 12943 41021 12952 41055
rect 12900 41012 12952 41021
rect 15476 41012 15528 41064
rect 15936 41123 15988 41132
rect 15936 41089 15950 41123
rect 15950 41089 15984 41123
rect 15984 41089 15988 41123
rect 15936 41080 15988 41089
rect 16120 41123 16172 41132
rect 16120 41089 16129 41123
rect 16129 41089 16163 41123
rect 16163 41089 16172 41123
rect 16120 41080 16172 41089
rect 17960 41216 18012 41268
rect 19340 41148 19392 41200
rect 19432 41148 19484 41200
rect 10968 40944 11020 40996
rect 16120 40944 16172 40996
rect 17960 41123 18012 41132
rect 17960 41089 17969 41123
rect 17969 41089 18003 41123
rect 18003 41089 18012 41123
rect 17960 41080 18012 41089
rect 23940 41080 23992 41132
rect 27804 41080 27856 41132
rect 18420 41012 18472 41064
rect 27712 41055 27764 41064
rect 17960 40944 18012 40996
rect 6920 40876 6972 40928
rect 8116 40919 8168 40928
rect 8116 40885 8125 40919
rect 8125 40885 8159 40919
rect 8159 40885 8168 40919
rect 8116 40876 8168 40885
rect 11428 40876 11480 40928
rect 11520 40919 11572 40928
rect 11520 40885 11529 40919
rect 11529 40885 11563 40919
rect 11563 40885 11572 40919
rect 11520 40876 11572 40885
rect 11704 40876 11756 40928
rect 13820 40876 13872 40928
rect 15476 40919 15528 40928
rect 15476 40885 15485 40919
rect 15485 40885 15519 40919
rect 15519 40885 15528 40919
rect 15476 40876 15528 40885
rect 18604 40876 18656 40928
rect 18696 40919 18748 40928
rect 18696 40885 18705 40919
rect 18705 40885 18739 40919
rect 18739 40885 18748 40919
rect 18696 40876 18748 40885
rect 19340 40876 19392 40928
rect 27712 41021 27721 41055
rect 27721 41021 27755 41055
rect 27755 41021 27764 41055
rect 27712 41012 27764 41021
rect 23112 40919 23164 40928
rect 23112 40885 23121 40919
rect 23121 40885 23155 40919
rect 23155 40885 23164 40919
rect 23112 40876 23164 40885
rect 29276 40876 29328 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 9312 40672 9364 40724
rect 27804 40715 27856 40724
rect 27804 40681 27813 40715
rect 27813 40681 27847 40715
rect 27847 40681 27856 40715
rect 27804 40672 27856 40681
rect 27712 40536 27764 40588
rect 29920 40579 29972 40588
rect 29920 40545 29929 40579
rect 29929 40545 29963 40579
rect 29963 40545 29972 40579
rect 29920 40536 29972 40545
rect 4436 40511 4488 40520
rect 4436 40477 4445 40511
rect 4445 40477 4479 40511
rect 4479 40477 4488 40511
rect 4436 40468 4488 40477
rect 4620 40511 4672 40520
rect 4620 40477 4629 40511
rect 4629 40477 4663 40511
rect 4663 40477 4672 40511
rect 4620 40468 4672 40477
rect 4712 40511 4764 40520
rect 4712 40477 4724 40511
rect 4724 40477 4758 40511
rect 4758 40477 4764 40511
rect 4712 40468 4764 40477
rect 5172 40468 5224 40520
rect 6920 40511 6972 40520
rect 6920 40477 6929 40511
rect 6929 40477 6963 40511
rect 6963 40477 6972 40511
rect 6920 40468 6972 40477
rect 8484 40468 8536 40520
rect 10508 40468 10560 40520
rect 12900 40511 12952 40520
rect 12900 40477 12909 40511
rect 12909 40477 12943 40511
rect 12943 40477 12952 40511
rect 14924 40511 14976 40520
rect 12900 40468 12952 40477
rect 14924 40477 14933 40511
rect 14933 40477 14967 40511
rect 14967 40477 14976 40511
rect 14924 40468 14976 40477
rect 16856 40468 16908 40520
rect 19340 40468 19392 40520
rect 25964 40468 26016 40520
rect 27252 40468 27304 40520
rect 28448 40511 28500 40520
rect 7012 40400 7064 40452
rect 8116 40400 8168 40452
rect 5080 40375 5132 40384
rect 5080 40341 5089 40375
rect 5089 40341 5123 40375
rect 5123 40341 5132 40375
rect 5080 40332 5132 40341
rect 5540 40375 5592 40384
rect 5540 40341 5549 40375
rect 5549 40341 5583 40375
rect 5583 40341 5592 40375
rect 5540 40332 5592 40341
rect 9036 40400 9088 40452
rect 10232 40400 10284 40452
rect 12532 40400 12584 40452
rect 15476 40400 15528 40452
rect 18512 40443 18564 40452
rect 18512 40409 18521 40443
rect 18521 40409 18555 40443
rect 18555 40409 18564 40443
rect 18512 40400 18564 40409
rect 18604 40400 18656 40452
rect 23480 40400 23532 40452
rect 23756 40400 23808 40452
rect 9864 40332 9916 40384
rect 10600 40332 10652 40384
rect 12440 40332 12492 40384
rect 15568 40332 15620 40384
rect 16304 40375 16356 40384
rect 16304 40341 16313 40375
rect 16313 40341 16347 40375
rect 16347 40341 16356 40375
rect 16304 40332 16356 40341
rect 18788 40332 18840 40384
rect 22652 40332 22704 40384
rect 24308 40332 24360 40384
rect 28448 40477 28457 40511
rect 28457 40477 28491 40511
rect 28491 40477 28500 40511
rect 28448 40468 28500 40477
rect 58164 40511 58216 40520
rect 58164 40477 58173 40511
rect 58173 40477 58207 40511
rect 58207 40477 58216 40511
rect 58164 40468 58216 40477
rect 29552 40400 29604 40452
rect 30288 40400 30340 40452
rect 28908 40332 28960 40384
rect 29092 40332 29144 40384
rect 30012 40332 30064 40384
rect 31852 40332 31904 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 6000 40128 6052 40180
rect 9772 40171 9824 40180
rect 9772 40137 9781 40171
rect 9781 40137 9815 40171
rect 9815 40137 9824 40171
rect 9772 40128 9824 40137
rect 5540 40060 5592 40112
rect 8576 40060 8628 40112
rect 9036 40060 9088 40112
rect 10324 40060 10376 40112
rect 2412 40035 2464 40044
rect 2412 40001 2446 40035
rect 2446 40001 2464 40035
rect 2412 39992 2464 40001
rect 4068 39924 4120 39976
rect 3240 39856 3292 39908
rect 4436 39924 4488 39976
rect 7104 39992 7156 40044
rect 8484 39992 8536 40044
rect 9220 39992 9272 40044
rect 7012 39967 7064 39976
rect 7012 39933 7021 39967
rect 7021 39933 7055 39967
rect 7055 39933 7064 39967
rect 7012 39924 7064 39933
rect 10232 39967 10284 39976
rect 10232 39933 10241 39967
rect 10241 39933 10275 39967
rect 10275 39933 10284 39967
rect 10232 39924 10284 39933
rect 4712 39856 4764 39908
rect 6644 39856 6696 39908
rect 9956 39856 10008 39908
rect 10692 40035 10744 40044
rect 10692 40001 10701 40035
rect 10701 40001 10735 40035
rect 10735 40001 10744 40035
rect 10692 39992 10744 40001
rect 11428 40060 11480 40112
rect 18788 40103 18840 40112
rect 11612 39992 11664 40044
rect 18788 40069 18797 40103
rect 18797 40069 18831 40103
rect 18831 40069 18840 40103
rect 18788 40060 18840 40069
rect 12992 40035 13044 40044
rect 2780 39788 2832 39840
rect 3976 39788 4028 39840
rect 10232 39788 10284 39840
rect 12532 39924 12584 39976
rect 12992 40001 13001 40035
rect 13001 40001 13035 40035
rect 13035 40001 13044 40035
rect 12992 39992 13044 40001
rect 18420 39992 18472 40044
rect 18972 40035 19024 40044
rect 18972 40001 18981 40035
rect 18981 40001 19015 40035
rect 19015 40001 19024 40035
rect 18972 39992 19024 40001
rect 19156 39992 19208 40044
rect 19340 39992 19392 40044
rect 20168 40035 20220 40044
rect 20168 40001 20202 40035
rect 20202 40001 20220 40035
rect 20168 39992 20220 40001
rect 22284 39992 22336 40044
rect 22560 40035 22612 40044
rect 22560 40001 22569 40035
rect 22569 40001 22603 40035
rect 22603 40001 22612 40035
rect 22560 39992 22612 40001
rect 23112 40060 23164 40112
rect 24952 40060 25004 40112
rect 12900 39924 12952 39976
rect 13360 39924 13412 39976
rect 23204 39992 23256 40044
rect 27712 40128 27764 40180
rect 29000 40128 29052 40180
rect 30288 40171 30340 40180
rect 30288 40137 30297 40171
rect 30297 40137 30331 40171
rect 30331 40137 30340 40171
rect 30288 40128 30340 40137
rect 19432 39856 19484 39908
rect 11612 39831 11664 39840
rect 11612 39797 11621 39831
rect 11621 39797 11655 39831
rect 11655 39797 11664 39831
rect 11612 39788 11664 39797
rect 16672 39831 16724 39840
rect 16672 39797 16681 39831
rect 16681 39797 16715 39831
rect 16715 39797 16724 39831
rect 16672 39788 16724 39797
rect 18512 39788 18564 39840
rect 22836 39924 22888 39976
rect 23756 39924 23808 39976
rect 25964 39924 26016 39976
rect 27712 40035 27764 40044
rect 27712 40001 27746 40035
rect 27746 40001 27764 40035
rect 27712 39992 27764 40001
rect 28448 39992 28500 40044
rect 31852 40060 31904 40112
rect 29184 39856 29236 39908
rect 30012 40035 30064 40044
rect 30012 40001 30021 40035
rect 30021 40001 30055 40035
rect 30055 40001 30064 40035
rect 30012 39992 30064 40001
rect 31208 39992 31260 40044
rect 30104 39856 30156 39908
rect 20260 39788 20312 39840
rect 21272 39831 21324 39840
rect 21272 39797 21281 39831
rect 21281 39797 21315 39831
rect 21315 39797 21324 39831
rect 21272 39788 21324 39797
rect 23664 39788 23716 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 2412 39584 2464 39636
rect 6368 39627 6420 39636
rect 6368 39593 6377 39627
rect 6377 39593 6411 39627
rect 6411 39593 6420 39627
rect 6368 39584 6420 39593
rect 9220 39627 9272 39636
rect 9220 39593 9229 39627
rect 9229 39593 9263 39627
rect 9263 39593 9272 39627
rect 9220 39584 9272 39593
rect 10692 39627 10744 39636
rect 10692 39593 10701 39627
rect 10701 39593 10735 39627
rect 10735 39593 10744 39627
rect 10692 39584 10744 39593
rect 20168 39584 20220 39636
rect 20352 39584 20404 39636
rect 22560 39584 22612 39636
rect 23204 39627 23256 39636
rect 23204 39593 23213 39627
rect 23213 39593 23247 39627
rect 23247 39593 23256 39627
rect 23204 39584 23256 39593
rect 29552 39627 29604 39636
rect 29552 39593 29561 39627
rect 29561 39593 29595 39627
rect 29595 39593 29604 39627
rect 29552 39584 29604 39593
rect 2872 39423 2924 39432
rect 2872 39389 2881 39423
rect 2881 39389 2915 39423
rect 2915 39389 2924 39423
rect 2872 39380 2924 39389
rect 4712 39448 4764 39500
rect 3240 39423 3292 39432
rect 2596 39312 2648 39364
rect 3240 39389 3249 39423
rect 3249 39389 3283 39423
rect 3283 39389 3292 39423
rect 3240 39380 3292 39389
rect 3792 39380 3844 39432
rect 5080 39380 5132 39432
rect 3976 39355 4028 39364
rect 3976 39321 3985 39355
rect 3985 39321 4019 39355
rect 4019 39321 4028 39355
rect 3976 39312 4028 39321
rect 6000 39312 6052 39364
rect 9680 39423 9732 39432
rect 9680 39389 9689 39423
rect 9689 39389 9723 39423
rect 9723 39389 9732 39423
rect 9680 39380 9732 39389
rect 10324 39423 10376 39432
rect 9956 39312 10008 39364
rect 10324 39389 10333 39423
rect 10333 39389 10367 39423
rect 10367 39389 10376 39423
rect 10324 39380 10376 39389
rect 10232 39312 10284 39364
rect 10600 39312 10652 39364
rect 19984 39516 20036 39568
rect 19524 39448 19576 39500
rect 19340 39312 19392 39364
rect 20352 39380 20404 39432
rect 22100 39380 22152 39432
rect 22284 39380 22336 39432
rect 19984 39312 20036 39364
rect 24308 39448 24360 39500
rect 22836 39423 22888 39432
rect 22836 39389 22845 39423
rect 22845 39389 22879 39423
rect 22879 39389 22888 39423
rect 22836 39380 22888 39389
rect 23112 39380 23164 39432
rect 31760 39380 31812 39432
rect 33324 39380 33376 39432
rect 23848 39312 23900 39364
rect 29276 39312 29328 39364
rect 32128 39355 32180 39364
rect 32128 39321 32162 39355
rect 32162 39321 32180 39355
rect 14372 39244 14424 39296
rect 17960 39244 18012 39296
rect 19248 39244 19300 39296
rect 25964 39244 26016 39296
rect 32128 39312 32180 39321
rect 30380 39244 30432 39296
rect 31668 39244 31720 39296
rect 33232 39287 33284 39296
rect 33232 39253 33241 39287
rect 33241 39253 33275 39287
rect 33275 39253 33284 39287
rect 33232 39244 33284 39253
rect 34520 39244 34572 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4068 39040 4120 39092
rect 12072 39040 12124 39092
rect 19340 39040 19392 39092
rect 23480 39040 23532 39092
rect 23848 39083 23900 39092
rect 23848 39049 23857 39083
rect 23857 39049 23891 39083
rect 23891 39049 23900 39083
rect 23848 39040 23900 39049
rect 27712 39083 27764 39092
rect 27712 39049 27721 39083
rect 27721 39049 27755 39083
rect 27755 39049 27764 39083
rect 27712 39040 27764 39049
rect 32128 39083 32180 39092
rect 32128 39049 32137 39083
rect 32137 39049 32171 39083
rect 32171 39049 32180 39083
rect 32128 39040 32180 39049
rect 21916 38972 21968 39024
rect 5724 38904 5776 38956
rect 16672 38904 16724 38956
rect 19156 38947 19208 38956
rect 19156 38913 19165 38947
rect 19165 38913 19199 38947
rect 19199 38913 19208 38947
rect 19156 38904 19208 38913
rect 19340 38947 19392 38956
rect 19340 38913 19349 38947
rect 19349 38913 19383 38947
rect 19383 38913 19392 38947
rect 19340 38904 19392 38913
rect 21272 38904 21324 38956
rect 22284 38904 22336 38956
rect 22560 38947 22612 38956
rect 22560 38913 22569 38947
rect 22569 38913 22603 38947
rect 22603 38913 22612 38947
rect 22560 38904 22612 38913
rect 30380 38972 30432 39024
rect 31208 38972 31260 39024
rect 13360 38879 13412 38888
rect 13360 38845 13369 38879
rect 13369 38845 13403 38879
rect 13403 38845 13412 38879
rect 13360 38836 13412 38845
rect 20352 38836 20404 38888
rect 13268 38768 13320 38820
rect 22192 38836 22244 38888
rect 22928 38904 22980 38956
rect 23664 38947 23716 38956
rect 23664 38913 23673 38947
rect 23673 38913 23707 38947
rect 23707 38913 23716 38947
rect 23664 38904 23716 38913
rect 22836 38836 22888 38888
rect 23572 38768 23624 38820
rect 2872 38700 2924 38752
rect 4712 38700 4764 38752
rect 10508 38700 10560 38752
rect 11612 38700 11664 38752
rect 16396 38700 16448 38752
rect 21916 38743 21968 38752
rect 21916 38709 21925 38743
rect 21925 38709 21959 38743
rect 21959 38709 21968 38743
rect 21916 38700 21968 38709
rect 26976 38700 27028 38752
rect 28448 38904 28500 38956
rect 29000 38947 29052 38956
rect 29000 38913 29009 38947
rect 29009 38913 29043 38947
rect 29043 38913 29052 38947
rect 29000 38904 29052 38913
rect 29920 38904 29972 38956
rect 30472 38947 30524 38956
rect 30472 38913 30506 38947
rect 30506 38913 30524 38947
rect 30472 38904 30524 38913
rect 31668 38904 31720 38956
rect 33140 38972 33192 39024
rect 32588 38947 32640 38956
rect 32588 38913 32597 38947
rect 32597 38913 32631 38947
rect 32631 38913 32640 38947
rect 32588 38904 32640 38913
rect 30104 38768 30156 38820
rect 33508 38904 33560 38956
rect 34520 38904 34572 38956
rect 35348 38904 35400 38956
rect 34796 38836 34848 38888
rect 36084 38836 36136 38888
rect 58164 38811 58216 38820
rect 58164 38777 58173 38811
rect 58173 38777 58207 38811
rect 58207 38777 58216 38811
rect 58164 38768 58216 38777
rect 28448 38700 28500 38752
rect 31116 38700 31168 38752
rect 31944 38700 31996 38752
rect 34704 38700 34756 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 9680 38496 9732 38548
rect 13268 38496 13320 38548
rect 13544 38496 13596 38548
rect 19340 38496 19392 38548
rect 22560 38496 22612 38548
rect 23572 38496 23624 38548
rect 30472 38539 30524 38548
rect 12164 38471 12216 38480
rect 6644 38360 6696 38412
rect 12164 38437 12173 38471
rect 12173 38437 12207 38471
rect 12207 38437 12216 38471
rect 12164 38428 12216 38437
rect 3792 38335 3844 38344
rect 3792 38301 3801 38335
rect 3801 38301 3835 38335
rect 3835 38301 3844 38335
rect 3792 38292 3844 38301
rect 9772 38360 9824 38412
rect 13636 38428 13688 38480
rect 3884 38224 3936 38276
rect 6000 38267 6052 38276
rect 6000 38233 6009 38267
rect 6009 38233 6043 38267
rect 6043 38233 6052 38267
rect 6000 38224 6052 38233
rect 10324 38292 10376 38344
rect 12440 38292 12492 38344
rect 12624 38335 12676 38344
rect 12624 38301 12633 38335
rect 12633 38301 12667 38335
rect 12667 38301 12676 38335
rect 12624 38292 12676 38301
rect 12992 38335 13044 38344
rect 12992 38301 13001 38335
rect 13001 38301 13035 38335
rect 13035 38301 13044 38335
rect 15384 38360 15436 38412
rect 17408 38428 17460 38480
rect 18696 38428 18748 38480
rect 30472 38505 30481 38539
rect 30481 38505 30515 38539
rect 30515 38505 30524 38539
rect 30472 38496 30524 38505
rect 32588 38496 32640 38548
rect 31668 38428 31720 38480
rect 33508 38428 33560 38480
rect 12992 38292 13044 38301
rect 12808 38267 12860 38276
rect 12808 38233 12817 38267
rect 12817 38233 12851 38267
rect 12851 38233 12860 38267
rect 12808 38224 12860 38233
rect 13820 38224 13872 38276
rect 3148 38199 3200 38208
rect 3148 38165 3157 38199
rect 3157 38165 3191 38199
rect 3191 38165 3200 38199
rect 3148 38156 3200 38165
rect 5264 38156 5316 38208
rect 5540 38156 5592 38208
rect 9864 38156 9916 38208
rect 12624 38156 12676 38208
rect 13360 38156 13412 38208
rect 18328 38360 18380 38412
rect 15108 38224 15160 38276
rect 15476 38156 15528 38208
rect 22652 38335 22704 38344
rect 15844 38224 15896 38276
rect 17408 38267 17460 38276
rect 17408 38233 17417 38267
rect 17417 38233 17451 38267
rect 17451 38233 17460 38267
rect 17408 38224 17460 38233
rect 22652 38301 22661 38335
rect 22661 38301 22695 38335
rect 22695 38301 22704 38335
rect 22652 38292 22704 38301
rect 25964 38292 26016 38344
rect 33140 38360 33192 38412
rect 36084 38403 36136 38412
rect 16488 38156 16540 38208
rect 18604 38224 18656 38276
rect 18972 38224 19024 38276
rect 22100 38224 22152 38276
rect 22836 38224 22888 38276
rect 27712 38224 27764 38276
rect 31116 38335 31168 38344
rect 30104 38224 30156 38276
rect 31116 38301 31125 38335
rect 31125 38301 31159 38335
rect 31159 38301 31168 38335
rect 31116 38292 31168 38301
rect 33232 38292 33284 38344
rect 33692 38335 33744 38344
rect 31208 38224 31260 38276
rect 31944 38224 31996 38276
rect 32680 38224 32732 38276
rect 33416 38224 33468 38276
rect 33692 38301 33701 38335
rect 33701 38301 33735 38335
rect 33735 38301 33744 38335
rect 33692 38292 33744 38301
rect 36084 38369 36093 38403
rect 36093 38369 36127 38403
rect 36127 38369 36136 38403
rect 36084 38360 36136 38369
rect 34520 38292 34572 38344
rect 33600 38224 33652 38276
rect 18512 38156 18564 38208
rect 19340 38156 19392 38208
rect 29000 38156 29052 38208
rect 29920 38199 29972 38208
rect 29920 38165 29929 38199
rect 29929 38165 29963 38199
rect 29963 38165 29972 38199
rect 29920 38156 29972 38165
rect 34060 38156 34112 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 2596 37952 2648 38004
rect 15108 37952 15160 38004
rect 6368 37884 6420 37936
rect 2872 37816 2924 37868
rect 3240 37816 3292 37868
rect 4620 37816 4672 37868
rect 5724 37816 5776 37868
rect 6828 37816 6880 37868
rect 11980 37884 12032 37936
rect 12808 37884 12860 37936
rect 8300 37859 8352 37868
rect 3148 37748 3200 37800
rect 2780 37680 2832 37732
rect 3792 37748 3844 37800
rect 8300 37825 8309 37859
rect 8309 37825 8343 37859
rect 8343 37825 8352 37859
rect 8300 37816 8352 37825
rect 8576 37859 8628 37868
rect 8576 37825 8585 37859
rect 8585 37825 8619 37859
rect 8619 37825 8628 37859
rect 8576 37816 8628 37825
rect 12992 37816 13044 37868
rect 13360 37859 13412 37868
rect 13360 37825 13369 37859
rect 13369 37825 13403 37859
rect 13403 37825 13412 37859
rect 13360 37816 13412 37825
rect 13452 37859 13504 37868
rect 13452 37825 13462 37859
rect 13462 37825 13496 37859
rect 13496 37825 13504 37859
rect 13636 37859 13688 37868
rect 13452 37816 13504 37825
rect 13636 37825 13645 37859
rect 13645 37825 13679 37859
rect 13679 37825 13688 37859
rect 13636 37816 13688 37825
rect 12808 37748 12860 37800
rect 13544 37748 13596 37800
rect 14004 37816 14056 37868
rect 15568 37884 15620 37936
rect 18788 37952 18840 38004
rect 20444 37952 20496 38004
rect 33692 37952 33744 38004
rect 34796 37952 34848 38004
rect 15476 37859 15528 37868
rect 15476 37825 15485 37859
rect 15485 37825 15519 37859
rect 15519 37825 15528 37859
rect 15476 37816 15528 37825
rect 16764 37816 16816 37868
rect 10600 37680 10652 37732
rect 13912 37680 13964 37732
rect 14096 37748 14148 37800
rect 14924 37748 14976 37800
rect 15200 37680 15252 37732
rect 16488 37680 16540 37732
rect 2320 37655 2372 37664
rect 2320 37621 2329 37655
rect 2329 37621 2363 37655
rect 2363 37621 2372 37655
rect 2320 37612 2372 37621
rect 5724 37655 5776 37664
rect 5724 37621 5733 37655
rect 5733 37621 5767 37655
rect 5767 37621 5776 37655
rect 5724 37612 5776 37621
rect 8668 37612 8720 37664
rect 8944 37612 8996 37664
rect 14464 37612 14516 37664
rect 17960 37612 18012 37664
rect 18328 37680 18380 37732
rect 18972 37859 19024 37868
rect 18972 37825 18986 37859
rect 18986 37825 19020 37859
rect 19020 37825 19024 37859
rect 18972 37816 19024 37825
rect 19340 37816 19392 37868
rect 19800 37859 19852 37868
rect 19800 37825 19809 37859
rect 19809 37825 19843 37859
rect 19843 37825 19852 37859
rect 19800 37816 19852 37825
rect 33416 37884 33468 37936
rect 24216 37816 24268 37868
rect 25136 37816 25188 37868
rect 31116 37816 31168 37868
rect 25964 37791 26016 37800
rect 25964 37757 25973 37791
rect 25973 37757 26007 37791
rect 26007 37757 26016 37791
rect 25964 37748 26016 37757
rect 19984 37680 20036 37732
rect 21180 37680 21232 37732
rect 18788 37612 18840 37664
rect 24032 37655 24084 37664
rect 24032 37621 24041 37655
rect 24041 37621 24075 37655
rect 24075 37621 24084 37655
rect 24032 37612 24084 37621
rect 24492 37612 24544 37664
rect 29828 37612 29880 37664
rect 32312 37748 32364 37800
rect 34060 37816 34112 37868
rect 34704 37816 34756 37868
rect 33600 37680 33652 37732
rect 34520 37612 34572 37664
rect 35532 37612 35584 37664
rect 58164 37655 58216 37664
rect 58164 37621 58173 37655
rect 58173 37621 58207 37655
rect 58207 37621 58216 37655
rect 58164 37612 58216 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2596 37408 2648 37460
rect 3884 37408 3936 37460
rect 15844 37408 15896 37460
rect 19800 37408 19852 37460
rect 11980 37315 12032 37324
rect 2320 37136 2372 37188
rect 2780 37136 2832 37188
rect 4436 37247 4488 37256
rect 4436 37213 4445 37247
rect 4445 37213 4479 37247
rect 4479 37213 4488 37247
rect 4436 37204 4488 37213
rect 11980 37281 11989 37315
rect 11989 37281 12023 37315
rect 12023 37281 12032 37315
rect 11980 37272 12032 37281
rect 14096 37315 14148 37324
rect 14096 37281 14105 37315
rect 14105 37281 14139 37315
rect 14139 37281 14148 37315
rect 14096 37272 14148 37281
rect 5356 37204 5408 37256
rect 4988 37179 5040 37188
rect 4988 37145 4997 37179
rect 4997 37145 5031 37179
rect 5031 37145 5040 37179
rect 4988 37136 5040 37145
rect 3056 37068 3108 37120
rect 3792 37068 3844 37120
rect 10324 37204 10376 37256
rect 12624 37204 12676 37256
rect 17960 37272 18012 37324
rect 18052 37247 18104 37256
rect 18052 37213 18061 37247
rect 18061 37213 18095 37247
rect 18095 37213 18104 37247
rect 18052 37204 18104 37213
rect 18604 37204 18656 37256
rect 18696 37204 18748 37256
rect 19156 37204 19208 37256
rect 20720 37204 20772 37256
rect 23388 37247 23440 37256
rect 10416 37179 10468 37188
rect 5632 37068 5684 37120
rect 10416 37145 10425 37179
rect 10425 37145 10459 37179
rect 10459 37145 10468 37179
rect 10416 37136 10468 37145
rect 14096 37136 14148 37188
rect 16948 37179 17000 37188
rect 16948 37145 16957 37179
rect 16957 37145 16991 37179
rect 16991 37145 17000 37179
rect 16948 37136 17000 37145
rect 18328 37179 18380 37188
rect 18328 37145 18337 37179
rect 18337 37145 18371 37179
rect 18371 37145 18380 37179
rect 18328 37136 18380 37145
rect 6184 37068 6236 37120
rect 6828 37111 6880 37120
rect 6828 37077 6837 37111
rect 6837 37077 6871 37111
rect 6871 37077 6880 37111
rect 6828 37068 6880 37077
rect 10600 37111 10652 37120
rect 10600 37077 10609 37111
rect 10609 37077 10643 37111
rect 10643 37077 10652 37111
rect 10600 37068 10652 37077
rect 16212 37068 16264 37120
rect 18604 37068 18656 37120
rect 21180 37179 21232 37188
rect 21180 37145 21198 37179
rect 21198 37145 21232 37179
rect 21180 37136 21232 37145
rect 22744 37111 22796 37120
rect 22744 37077 22753 37111
rect 22753 37077 22787 37111
rect 22787 37077 22796 37111
rect 22744 37068 22796 37077
rect 23388 37213 23397 37247
rect 23397 37213 23431 37247
rect 23431 37213 23440 37247
rect 23388 37204 23440 37213
rect 24676 37408 24728 37460
rect 32312 37451 32364 37460
rect 32312 37417 32321 37451
rect 32321 37417 32355 37451
rect 32355 37417 32364 37451
rect 32312 37408 32364 37417
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 25964 37204 26016 37256
rect 27896 37179 27948 37188
rect 27896 37145 27930 37179
rect 27930 37145 27948 37179
rect 27896 37136 27948 37145
rect 24032 37068 24084 37120
rect 25688 37068 25740 37120
rect 28632 37068 28684 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 2872 36907 2924 36916
rect 2872 36873 2881 36907
rect 2881 36873 2915 36907
rect 2915 36873 2924 36907
rect 2872 36864 2924 36873
rect 6000 36796 6052 36848
rect 10416 36864 10468 36916
rect 3056 36771 3108 36780
rect 3056 36737 3065 36771
rect 3065 36737 3099 36771
rect 3099 36737 3108 36771
rect 3056 36728 3108 36737
rect 10508 36796 10560 36848
rect 10140 36728 10192 36780
rect 11704 36864 11756 36916
rect 18052 36864 18104 36916
rect 12256 36796 12308 36848
rect 12440 36796 12492 36848
rect 12716 36796 12768 36848
rect 13452 36796 13504 36848
rect 15844 36796 15896 36848
rect 24492 36864 24544 36916
rect 24676 36864 24728 36916
rect 25136 36864 25188 36916
rect 27252 36907 27304 36916
rect 27252 36873 27261 36907
rect 27261 36873 27295 36907
rect 27295 36873 27304 36907
rect 27252 36864 27304 36873
rect 27712 36907 27764 36916
rect 27712 36873 27721 36907
rect 27721 36873 27755 36907
rect 27755 36873 27764 36907
rect 27712 36864 27764 36873
rect 12808 36728 12860 36780
rect 14832 36771 14884 36780
rect 14832 36737 14841 36771
rect 14841 36737 14875 36771
rect 14875 36737 14884 36771
rect 14832 36728 14884 36737
rect 16948 36728 17000 36780
rect 17132 36771 17184 36780
rect 17132 36737 17141 36771
rect 17141 36737 17175 36771
rect 17175 36737 17184 36771
rect 17132 36728 17184 36737
rect 17316 36771 17368 36780
rect 17316 36737 17325 36771
rect 17325 36737 17359 36771
rect 17359 36737 17368 36771
rect 17316 36728 17368 36737
rect 12624 36660 12676 36712
rect 16672 36660 16724 36712
rect 13084 36592 13136 36644
rect 22744 36728 22796 36780
rect 23296 36771 23348 36780
rect 20720 36660 20772 36712
rect 23296 36737 23305 36771
rect 23305 36737 23339 36771
rect 23339 36737 23348 36771
rect 23296 36728 23348 36737
rect 23664 36728 23716 36780
rect 24032 36728 24084 36780
rect 23388 36660 23440 36712
rect 24124 36660 24176 36712
rect 24860 36728 24912 36780
rect 25504 36771 25556 36780
rect 25504 36737 25513 36771
rect 25513 36737 25547 36771
rect 25547 36737 25556 36771
rect 25504 36728 25556 36737
rect 25688 36771 25740 36780
rect 25688 36737 25697 36771
rect 25697 36737 25731 36771
rect 25731 36737 25740 36771
rect 25688 36728 25740 36737
rect 28077 36771 28129 36780
rect 28077 36737 28104 36771
rect 28104 36737 28129 36771
rect 28077 36728 28129 36737
rect 33416 36771 33468 36780
rect 28264 36660 28316 36712
rect 33416 36737 33425 36771
rect 33425 36737 33459 36771
rect 33459 36737 33468 36771
rect 33416 36728 33468 36737
rect 34520 36728 34572 36780
rect 12256 36524 12308 36576
rect 12900 36524 12952 36576
rect 14556 36524 14608 36576
rect 18696 36524 18748 36576
rect 28172 36592 28224 36644
rect 31760 36592 31812 36644
rect 32036 36592 32088 36644
rect 36636 36592 36688 36644
rect 20812 36524 20864 36576
rect 22468 36567 22520 36576
rect 22468 36533 22477 36567
rect 22477 36533 22511 36567
rect 22511 36533 22520 36567
rect 22468 36524 22520 36533
rect 22560 36524 22612 36576
rect 23480 36524 23532 36576
rect 33784 36567 33836 36576
rect 33784 36533 33793 36567
rect 33793 36533 33827 36567
rect 33827 36533 33836 36567
rect 33784 36524 33836 36533
rect 35348 36524 35400 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 10140 36363 10192 36372
rect 10140 36329 10149 36363
rect 10149 36329 10183 36363
rect 10183 36329 10192 36363
rect 10140 36320 10192 36329
rect 13084 36320 13136 36372
rect 13452 36320 13504 36372
rect 14096 36363 14148 36372
rect 14096 36329 14105 36363
rect 14105 36329 14139 36363
rect 14139 36329 14148 36363
rect 14096 36320 14148 36329
rect 16764 36320 16816 36372
rect 17316 36363 17368 36372
rect 17316 36329 17325 36363
rect 17325 36329 17359 36363
rect 17359 36329 17368 36363
rect 17316 36320 17368 36329
rect 20812 36363 20864 36372
rect 20812 36329 20821 36363
rect 20821 36329 20855 36363
rect 20855 36329 20864 36363
rect 20812 36320 20864 36329
rect 24124 36320 24176 36372
rect 27896 36320 27948 36372
rect 33324 36363 33376 36372
rect 33324 36329 33333 36363
rect 33333 36329 33367 36363
rect 33367 36329 33376 36363
rect 33324 36320 33376 36329
rect 36636 36363 36688 36372
rect 36636 36329 36645 36363
rect 36645 36329 36679 36363
rect 36679 36329 36688 36363
rect 36636 36320 36688 36329
rect 8300 36184 8352 36236
rect 6092 36159 6144 36168
rect 6092 36125 6101 36159
rect 6101 36125 6135 36159
rect 6135 36125 6144 36159
rect 6092 36116 6144 36125
rect 28080 36252 28132 36304
rect 6920 36048 6972 36100
rect 7380 36048 7432 36100
rect 8300 36091 8352 36100
rect 8300 36057 8309 36091
rect 8309 36057 8343 36091
rect 8343 36057 8352 36091
rect 8300 36048 8352 36057
rect 9956 36048 10008 36100
rect 10600 36159 10652 36168
rect 10600 36125 10609 36159
rect 10609 36125 10643 36159
rect 10643 36125 10652 36159
rect 10600 36116 10652 36125
rect 10876 36116 10928 36168
rect 14372 36159 14424 36168
rect 4988 35980 5040 36032
rect 5540 35980 5592 36032
rect 10416 35980 10468 36032
rect 10508 35980 10560 36032
rect 14372 36125 14381 36159
rect 14381 36125 14415 36159
rect 14415 36125 14424 36159
rect 14372 36116 14424 36125
rect 14648 36184 14700 36236
rect 14556 36159 14608 36168
rect 14556 36125 14565 36159
rect 14565 36125 14599 36159
rect 14599 36125 14608 36159
rect 14556 36116 14608 36125
rect 16212 36159 16264 36168
rect 12440 36048 12492 36100
rect 13912 36048 13964 36100
rect 16212 36125 16221 36159
rect 16221 36125 16255 36159
rect 16255 36125 16264 36159
rect 16212 36116 16264 36125
rect 16672 36184 16724 36236
rect 16396 36159 16448 36168
rect 16396 36125 16405 36159
rect 16405 36125 16439 36159
rect 16439 36125 16448 36159
rect 16396 36116 16448 36125
rect 17040 36116 17092 36168
rect 17132 36048 17184 36100
rect 18696 36116 18748 36168
rect 20812 36116 20864 36168
rect 17684 36091 17736 36100
rect 17684 36057 17693 36091
rect 17693 36057 17727 36091
rect 17727 36057 17736 36091
rect 17684 36048 17736 36057
rect 21824 36159 21876 36168
rect 21824 36125 21833 36159
rect 21833 36125 21867 36159
rect 21867 36125 21876 36159
rect 21824 36116 21876 36125
rect 22284 36116 22336 36168
rect 22652 36116 22704 36168
rect 25688 36184 25740 36236
rect 23480 36159 23532 36168
rect 23480 36125 23489 36159
rect 23489 36125 23523 36159
rect 23523 36125 23532 36159
rect 23480 36116 23532 36125
rect 24492 36116 24544 36168
rect 24860 36116 24912 36168
rect 25504 36116 25556 36168
rect 27804 36116 27856 36168
rect 28448 36184 28500 36236
rect 33508 36184 33560 36236
rect 28264 36159 28316 36168
rect 22192 36048 22244 36100
rect 22468 36048 22520 36100
rect 23296 36091 23348 36100
rect 23296 36057 23305 36091
rect 23305 36057 23339 36091
rect 23339 36057 23348 36091
rect 23296 36048 23348 36057
rect 27620 36048 27672 36100
rect 14372 35980 14424 36032
rect 15568 35980 15620 36032
rect 22376 35980 22428 36032
rect 22652 36023 22704 36032
rect 22652 35989 22661 36023
rect 22661 35989 22695 36023
rect 22695 35989 22704 36023
rect 22652 35980 22704 35989
rect 23664 36023 23716 36032
rect 23664 35989 23673 36023
rect 23673 35989 23707 36023
rect 23707 35989 23716 36023
rect 23664 35980 23716 35989
rect 24492 35980 24544 36032
rect 24768 35980 24820 36032
rect 27804 35980 27856 36032
rect 28264 36125 28273 36159
rect 28273 36125 28307 36159
rect 28307 36125 28316 36159
rect 28264 36116 28316 36125
rect 33600 36116 33652 36168
rect 30104 36091 30156 36100
rect 30104 36057 30113 36091
rect 30113 36057 30147 36091
rect 30147 36057 30156 36091
rect 30104 36048 30156 36057
rect 30932 36048 30984 36100
rect 28540 35980 28592 36032
rect 30840 36023 30892 36032
rect 30840 35989 30849 36023
rect 30849 35989 30883 36023
rect 30883 35989 30892 36023
rect 30840 35980 30892 35989
rect 31116 36048 31168 36100
rect 32036 36091 32088 36100
rect 32036 36057 32045 36091
rect 32045 36057 32079 36091
rect 32079 36057 32088 36091
rect 32036 36048 32088 36057
rect 33140 36048 33192 36100
rect 35348 36116 35400 36168
rect 58164 36159 58216 36168
rect 58164 36125 58173 36159
rect 58173 36125 58207 36159
rect 58207 36125 58216 36159
rect 58164 36116 58216 36125
rect 36084 36048 36136 36100
rect 38568 36048 38620 36100
rect 32404 35980 32456 36032
rect 34612 35980 34664 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 6920 35819 6972 35828
rect 6920 35785 6929 35819
rect 6929 35785 6963 35819
rect 6963 35785 6972 35819
rect 6920 35776 6972 35785
rect 12440 35819 12492 35828
rect 12440 35785 12449 35819
rect 12449 35785 12483 35819
rect 12483 35785 12492 35819
rect 12440 35776 12492 35785
rect 10324 35708 10376 35760
rect 4068 35640 4120 35692
rect 2780 35615 2832 35624
rect 2780 35581 2789 35615
rect 2789 35581 2823 35615
rect 2823 35581 2832 35615
rect 2780 35572 2832 35581
rect 4712 35436 4764 35488
rect 6276 35436 6328 35488
rect 7380 35683 7432 35692
rect 7380 35649 7389 35683
rect 7389 35649 7423 35683
rect 7423 35649 7432 35683
rect 7380 35640 7432 35649
rect 10232 35640 10284 35692
rect 10876 35708 10928 35760
rect 10968 35708 11020 35760
rect 11888 35640 11940 35692
rect 12900 35683 12952 35692
rect 12900 35649 12909 35683
rect 12909 35649 12943 35683
rect 12943 35649 12952 35683
rect 12900 35640 12952 35649
rect 7656 35572 7708 35624
rect 7564 35504 7616 35556
rect 16580 35776 16632 35828
rect 19340 35776 19392 35828
rect 19524 35776 19576 35828
rect 21824 35819 21876 35828
rect 21824 35785 21833 35819
rect 21833 35785 21867 35819
rect 21867 35785 21876 35819
rect 21824 35776 21876 35785
rect 24952 35776 25004 35828
rect 25688 35776 25740 35828
rect 28172 35776 28224 35828
rect 33140 35776 33192 35828
rect 22100 35708 22152 35760
rect 33324 35708 33376 35760
rect 21916 35640 21968 35692
rect 22836 35640 22888 35692
rect 27436 35640 27488 35692
rect 29000 35640 29052 35692
rect 29552 35683 29604 35692
rect 29552 35649 29561 35683
rect 29561 35649 29595 35683
rect 29595 35649 29604 35683
rect 29552 35640 29604 35649
rect 31116 35640 31168 35692
rect 14648 35572 14700 35624
rect 27344 35615 27396 35624
rect 27344 35581 27353 35615
rect 27353 35581 27387 35615
rect 27387 35581 27396 35615
rect 27344 35572 27396 35581
rect 30472 35572 30524 35624
rect 31208 35572 31260 35624
rect 31576 35572 31628 35624
rect 33048 35640 33100 35692
rect 34612 35640 34664 35692
rect 36084 35708 36136 35760
rect 34796 35640 34848 35692
rect 33140 35572 33192 35624
rect 33416 35572 33468 35624
rect 19340 35504 19392 35556
rect 23664 35504 23716 35556
rect 10692 35436 10744 35488
rect 16856 35436 16908 35488
rect 23388 35436 23440 35488
rect 24492 35436 24544 35488
rect 28264 35436 28316 35488
rect 33048 35436 33100 35488
rect 34520 35436 34572 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 11888 35275 11940 35284
rect 11888 35241 11897 35275
rect 11897 35241 11931 35275
rect 11931 35241 11940 35275
rect 11888 35232 11940 35241
rect 17224 35232 17276 35284
rect 27160 35232 27212 35284
rect 27436 35275 27488 35284
rect 27436 35241 27445 35275
rect 27445 35241 27479 35275
rect 27479 35241 27488 35275
rect 27436 35232 27488 35241
rect 28540 35275 28592 35284
rect 28540 35241 28549 35275
rect 28549 35241 28583 35275
rect 28583 35241 28592 35275
rect 28540 35232 28592 35241
rect 30932 35232 30984 35284
rect 10508 35139 10560 35148
rect 6184 35071 6236 35080
rect 6184 35037 6193 35071
rect 6193 35037 6227 35071
rect 6227 35037 6236 35071
rect 6184 35028 6236 35037
rect 10508 35105 10517 35139
rect 10517 35105 10551 35139
rect 10551 35105 10560 35139
rect 10508 35096 10560 35105
rect 4712 34960 4764 35012
rect 5264 34960 5316 35012
rect 5448 34960 5500 35012
rect 4804 34892 4856 34944
rect 5080 34935 5132 34944
rect 5080 34901 5089 34935
rect 5089 34901 5123 34935
rect 5123 34901 5132 34935
rect 5080 34892 5132 34901
rect 6000 34935 6052 34944
rect 6000 34901 6009 34935
rect 6009 34901 6043 34935
rect 6043 34901 6052 34935
rect 6000 34892 6052 34901
rect 6736 34960 6788 35012
rect 8300 35028 8352 35080
rect 17316 35164 17368 35216
rect 30288 35164 30340 35216
rect 12532 35096 12584 35148
rect 12808 35028 12860 35080
rect 16856 35071 16908 35080
rect 16856 35037 16865 35071
rect 16865 35037 16899 35071
rect 16899 35037 16908 35071
rect 16856 35028 16908 35037
rect 8576 34960 8628 35012
rect 11152 34960 11204 35012
rect 12440 34960 12492 35012
rect 16672 34960 16724 35012
rect 17132 35028 17184 35080
rect 17684 35071 17736 35080
rect 17684 35037 17693 35071
rect 17693 35037 17727 35071
rect 17727 35037 17736 35071
rect 17684 35028 17736 35037
rect 19340 35071 19392 35080
rect 19340 35037 19349 35071
rect 19349 35037 19383 35071
rect 19383 35037 19392 35071
rect 19340 35028 19392 35037
rect 19432 35028 19484 35080
rect 20076 35028 20128 35080
rect 28448 35096 28500 35148
rect 29736 35096 29788 35148
rect 17868 35003 17920 35012
rect 17868 34969 17877 35003
rect 17877 34969 17911 35003
rect 17911 34969 17920 35003
rect 17868 34960 17920 34969
rect 7932 34892 7984 34944
rect 16764 34892 16816 34944
rect 19340 34892 19392 34944
rect 19524 34892 19576 34944
rect 20720 34892 20772 34944
rect 22376 34960 22428 35012
rect 27988 35028 28040 35080
rect 28080 35071 28132 35080
rect 28080 35037 28089 35071
rect 28089 35037 28123 35071
rect 28123 35037 28132 35071
rect 28080 35028 28132 35037
rect 29552 35028 29604 35080
rect 29920 35028 29972 35080
rect 28632 34960 28684 35012
rect 30564 35028 30616 35080
rect 33324 35096 33376 35148
rect 33508 35139 33560 35148
rect 33508 35105 33517 35139
rect 33517 35105 33551 35139
rect 33551 35105 33560 35139
rect 33508 35096 33560 35105
rect 58164 35071 58216 35080
rect 58164 35037 58173 35071
rect 58173 35037 58207 35071
rect 58207 35037 58216 35071
rect 58164 35028 58216 35037
rect 30840 34960 30892 35012
rect 22100 34892 22152 34944
rect 26976 34935 27028 34944
rect 26976 34901 26985 34935
rect 26985 34901 27019 34935
rect 27019 34901 27028 34935
rect 26976 34892 27028 34901
rect 32404 34892 32456 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 2780 34688 2832 34740
rect 4068 34688 4120 34740
rect 8576 34731 8628 34740
rect 8576 34697 8585 34731
rect 8585 34697 8619 34731
rect 8619 34697 8628 34731
rect 8576 34688 8628 34697
rect 12072 34688 12124 34740
rect 17224 34688 17276 34740
rect 17500 34688 17552 34740
rect 17868 34688 17920 34740
rect 20076 34731 20128 34740
rect 20076 34697 20085 34731
rect 20085 34697 20119 34731
rect 20119 34697 20128 34731
rect 20076 34688 20128 34697
rect 27988 34731 28040 34740
rect 27988 34697 27997 34731
rect 27997 34697 28031 34731
rect 28031 34697 28040 34731
rect 27988 34688 28040 34697
rect 29184 34688 29236 34740
rect 29920 34688 29972 34740
rect 33140 34731 33192 34740
rect 33140 34697 33149 34731
rect 33149 34697 33183 34731
rect 33183 34697 33192 34731
rect 33140 34688 33192 34697
rect 34796 34688 34848 34740
rect 3792 34552 3844 34604
rect 4620 34595 4672 34604
rect 4620 34561 4629 34595
rect 4629 34561 4663 34595
rect 4663 34561 4672 34595
rect 4620 34552 4672 34561
rect 4804 34595 4856 34604
rect 4804 34561 4813 34595
rect 4813 34561 4847 34595
rect 4847 34561 4856 34595
rect 4804 34552 4856 34561
rect 5080 34552 5132 34604
rect 6092 34552 6144 34604
rect 6828 34552 6880 34604
rect 7472 34595 7524 34604
rect 7472 34561 7506 34595
rect 7506 34561 7524 34595
rect 7472 34552 7524 34561
rect 10232 34552 10284 34604
rect 12072 34552 12124 34604
rect 20720 34620 20772 34672
rect 16764 34552 16816 34604
rect 19156 34595 19208 34604
rect 19156 34561 19165 34595
rect 19165 34561 19199 34595
rect 19199 34561 19208 34595
rect 19156 34552 19208 34561
rect 19432 34552 19484 34604
rect 4896 34484 4948 34536
rect 10600 34527 10652 34536
rect 10600 34493 10609 34527
rect 10609 34493 10643 34527
rect 10643 34493 10652 34527
rect 10600 34484 10652 34493
rect 13176 34484 13228 34536
rect 27620 34620 27672 34672
rect 28080 34620 28132 34672
rect 29552 34620 29604 34672
rect 33508 34620 33560 34672
rect 24124 34595 24176 34604
rect 24124 34561 24142 34595
rect 24142 34561 24176 34595
rect 24124 34552 24176 34561
rect 24860 34595 24912 34604
rect 24860 34561 24869 34595
rect 24869 34561 24903 34595
rect 24903 34561 24912 34595
rect 24860 34552 24912 34561
rect 25044 34595 25096 34604
rect 25044 34561 25053 34595
rect 25053 34561 25087 34595
rect 25087 34561 25096 34595
rect 25044 34552 25096 34561
rect 28172 34595 28224 34604
rect 28172 34561 28181 34595
rect 28181 34561 28215 34595
rect 28215 34561 28224 34595
rect 28172 34552 28224 34561
rect 31576 34552 31628 34604
rect 33600 34595 33652 34604
rect 33600 34561 33609 34595
rect 33609 34561 33643 34595
rect 33643 34561 33652 34595
rect 33600 34552 33652 34561
rect 33784 34595 33836 34604
rect 33784 34561 33793 34595
rect 33793 34561 33827 34595
rect 33827 34561 33836 34595
rect 33784 34552 33836 34561
rect 4988 34348 5040 34400
rect 5080 34348 5132 34400
rect 7104 34348 7156 34400
rect 12532 34348 12584 34400
rect 26240 34484 26292 34536
rect 27344 34484 27396 34536
rect 27528 34484 27580 34536
rect 29828 34527 29880 34536
rect 29828 34493 29837 34527
rect 29837 34493 29871 34527
rect 29871 34493 29880 34527
rect 29828 34484 29880 34493
rect 30564 34527 30616 34536
rect 30564 34493 30573 34527
rect 30573 34493 30607 34527
rect 30607 34493 30616 34527
rect 30564 34484 30616 34493
rect 33416 34484 33468 34536
rect 24492 34416 24544 34468
rect 35348 34416 35400 34468
rect 19340 34348 19392 34400
rect 23020 34391 23072 34400
rect 23020 34357 23029 34391
rect 23029 34357 23063 34391
rect 23063 34357 23072 34391
rect 23020 34348 23072 34357
rect 25228 34391 25280 34400
rect 25228 34357 25237 34391
rect 25237 34357 25271 34391
rect 25271 34357 25280 34391
rect 25228 34348 25280 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 3792 34187 3844 34196
rect 3792 34153 3801 34187
rect 3801 34153 3835 34187
rect 3835 34153 3844 34187
rect 3792 34144 3844 34153
rect 5632 34187 5684 34196
rect 5632 34153 5641 34187
rect 5641 34153 5675 34187
rect 5675 34153 5684 34187
rect 5632 34144 5684 34153
rect 7104 34144 7156 34196
rect 7472 34187 7524 34196
rect 7472 34153 7481 34187
rect 7481 34153 7515 34187
rect 7515 34153 7524 34187
rect 7472 34144 7524 34153
rect 11152 34187 11204 34196
rect 11152 34153 11161 34187
rect 11161 34153 11195 34187
rect 11195 34153 11204 34187
rect 11152 34144 11204 34153
rect 12532 34144 12584 34196
rect 29184 34144 29236 34196
rect 35348 34187 35400 34196
rect 35348 34153 35357 34187
rect 35357 34153 35391 34187
rect 35391 34153 35400 34187
rect 35348 34144 35400 34153
rect 3424 34008 3476 34060
rect 3148 33940 3200 33992
rect 4068 33983 4120 33992
rect 4068 33949 4077 33983
rect 4077 33949 4111 33983
rect 4111 33949 4120 33983
rect 4068 33940 4120 33949
rect 4252 33983 4304 33992
rect 4252 33949 4261 33983
rect 4261 33949 4295 33983
rect 4295 33949 4304 33983
rect 4252 33940 4304 33949
rect 5080 33940 5132 33992
rect 5908 33983 5960 33992
rect 5908 33949 5917 33983
rect 5917 33949 5951 33983
rect 5951 33949 5960 33983
rect 5908 33940 5960 33949
rect 7656 34008 7708 34060
rect 8208 34008 8260 34060
rect 6092 33983 6144 33992
rect 6092 33949 6101 33983
rect 6101 33949 6135 33983
rect 6135 33949 6144 33983
rect 6092 33940 6144 33949
rect 4896 33872 4948 33924
rect 7104 33940 7156 33992
rect 7932 33983 7984 33992
rect 7932 33949 7946 33983
rect 7946 33949 7980 33983
rect 7980 33949 7984 33983
rect 7932 33940 7984 33949
rect 8944 33983 8996 33992
rect 8024 33872 8076 33924
rect 3332 33804 3384 33856
rect 6184 33804 6236 33856
rect 8944 33949 8953 33983
rect 8953 33949 8987 33983
rect 8987 33949 8996 33983
rect 8944 33940 8996 33949
rect 13728 34076 13780 34128
rect 9864 34008 9916 34060
rect 10416 34008 10468 34060
rect 10140 33940 10192 33992
rect 10232 33940 10284 33992
rect 10692 33983 10744 33992
rect 10692 33949 10701 33983
rect 10701 33949 10735 33983
rect 10735 33949 10744 33983
rect 10692 33940 10744 33949
rect 16856 34076 16908 34128
rect 14648 34008 14700 34060
rect 13728 33940 13780 33992
rect 8576 33872 8628 33924
rect 8300 33804 8352 33856
rect 9588 33847 9640 33856
rect 9588 33813 9597 33847
rect 9597 33813 9631 33847
rect 9631 33813 9640 33847
rect 9588 33804 9640 33813
rect 10600 33872 10652 33924
rect 13912 33872 13964 33924
rect 14188 33940 14240 33992
rect 17316 33983 17368 33992
rect 17316 33949 17325 33983
rect 17325 33949 17359 33983
rect 17359 33949 17368 33983
rect 17316 33940 17368 33949
rect 17500 33983 17552 33992
rect 17500 33949 17507 33983
rect 17507 33949 17552 33983
rect 17500 33940 17552 33949
rect 17776 33983 17828 33992
rect 17776 33949 17790 33983
rect 17790 33949 17824 33983
rect 17824 33949 17828 33983
rect 20720 34051 20772 34060
rect 20720 34017 20729 34051
rect 20729 34017 20763 34051
rect 20763 34017 20772 34051
rect 20720 34008 20772 34017
rect 22376 34008 22428 34060
rect 22652 34008 22704 34060
rect 17776 33940 17828 33949
rect 20168 33940 20220 33992
rect 23388 33983 23440 33992
rect 16580 33872 16632 33924
rect 19248 33804 19300 33856
rect 19432 33872 19484 33924
rect 19984 33872 20036 33924
rect 23388 33949 23397 33983
rect 23397 33949 23431 33983
rect 23431 33949 23440 33983
rect 23388 33940 23440 33949
rect 24308 33940 24360 33992
rect 23020 33872 23072 33924
rect 24216 33872 24268 33924
rect 24952 34008 25004 34060
rect 24584 33940 24636 33992
rect 25207 33983 25259 33992
rect 25207 33949 25216 33983
rect 25216 33949 25250 33983
rect 25250 33949 25259 33983
rect 25207 33940 25259 33949
rect 27528 34051 27580 34060
rect 27528 34017 27537 34051
rect 27537 34017 27571 34051
rect 27571 34017 27580 34051
rect 27528 34008 27580 34017
rect 30288 34051 30340 34060
rect 30288 34017 30297 34051
rect 30297 34017 30331 34051
rect 30331 34017 30340 34051
rect 30288 34008 30340 34017
rect 35900 33983 35952 33992
rect 35900 33949 35909 33983
rect 35909 33949 35943 33983
rect 35943 33949 35952 33983
rect 35900 33940 35952 33949
rect 36084 33983 36136 33992
rect 36084 33949 36093 33983
rect 36093 33949 36127 33983
rect 36127 33949 36136 33983
rect 36084 33940 36136 33949
rect 29644 33872 29696 33924
rect 31116 33872 31168 33924
rect 22376 33804 22428 33856
rect 22744 33847 22796 33856
rect 22744 33813 22753 33847
rect 22753 33813 22787 33847
rect 22787 33813 22796 33847
rect 22744 33804 22796 33813
rect 23204 33847 23256 33856
rect 23204 33813 23213 33847
rect 23213 33813 23247 33847
rect 23247 33813 23256 33847
rect 23204 33804 23256 33813
rect 23572 33804 23624 33856
rect 24860 33804 24912 33856
rect 25044 33804 25096 33856
rect 31484 33804 31536 33856
rect 36452 33872 36504 33924
rect 32496 33847 32548 33856
rect 32496 33813 32505 33847
rect 32505 33813 32539 33847
rect 32539 33813 32548 33847
rect 32496 33804 32548 33813
rect 33416 33847 33468 33856
rect 33416 33813 33425 33847
rect 33425 33813 33459 33847
rect 33459 33813 33468 33847
rect 33416 33804 33468 33813
rect 38200 33804 38252 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4252 33600 4304 33652
rect 4896 33600 4948 33652
rect 6644 33600 6696 33652
rect 8300 33643 8352 33652
rect 8300 33609 8309 33643
rect 8309 33609 8343 33643
rect 8343 33609 8352 33643
rect 8300 33600 8352 33609
rect 10324 33600 10376 33652
rect 14832 33600 14884 33652
rect 19340 33600 19392 33652
rect 19984 33600 20036 33652
rect 24124 33600 24176 33652
rect 24400 33600 24452 33652
rect 24768 33600 24820 33652
rect 24952 33600 25004 33652
rect 29092 33643 29144 33652
rect 29092 33609 29101 33643
rect 29101 33609 29135 33643
rect 29135 33609 29144 33643
rect 29092 33600 29144 33609
rect 29644 33643 29696 33652
rect 29644 33609 29653 33643
rect 29653 33609 29687 33643
rect 29687 33609 29696 33643
rect 29644 33600 29696 33609
rect 29736 33600 29788 33652
rect 4712 33532 4764 33584
rect 4988 33575 5040 33584
rect 4988 33541 4997 33575
rect 4997 33541 5031 33575
rect 5031 33541 5040 33575
rect 4988 33532 5040 33541
rect 6736 33532 6788 33584
rect 8024 33532 8076 33584
rect 10140 33532 10192 33584
rect 15200 33532 15252 33584
rect 16948 33532 17000 33584
rect 17776 33532 17828 33584
rect 9128 33507 9180 33516
rect 9128 33473 9137 33507
rect 9137 33473 9171 33507
rect 9171 33473 9180 33507
rect 9128 33464 9180 33473
rect 10600 33507 10652 33516
rect 4988 33396 5040 33448
rect 10600 33473 10609 33507
rect 10609 33473 10643 33507
rect 10643 33473 10652 33507
rect 10600 33464 10652 33473
rect 15016 33464 15068 33516
rect 19064 33507 19116 33516
rect 19064 33473 19073 33507
rect 19073 33473 19107 33507
rect 19107 33473 19116 33507
rect 19064 33464 19116 33473
rect 23020 33532 23072 33584
rect 23572 33575 23624 33584
rect 23572 33541 23581 33575
rect 23581 33541 23615 33575
rect 23615 33541 23624 33575
rect 23572 33532 23624 33541
rect 23940 33532 23992 33584
rect 17132 33396 17184 33448
rect 20260 33464 20312 33516
rect 22928 33464 22980 33516
rect 24584 33532 24636 33584
rect 24387 33507 24439 33519
rect 24387 33473 24409 33507
rect 24409 33473 24439 33507
rect 24387 33467 24439 33473
rect 20076 33396 20128 33448
rect 6184 33328 6236 33380
rect 10692 33328 10744 33380
rect 25136 33507 25188 33516
rect 25136 33473 25145 33507
rect 25145 33473 25179 33507
rect 25179 33473 25188 33507
rect 25136 33464 25188 33473
rect 31208 33600 31260 33652
rect 33416 33600 33468 33652
rect 32496 33532 32548 33584
rect 30564 33464 30616 33516
rect 35900 33532 35952 33584
rect 35992 33507 36044 33516
rect 35992 33473 36001 33507
rect 36001 33473 36035 33507
rect 36035 33473 36044 33507
rect 35992 33464 36044 33473
rect 38568 33464 38620 33516
rect 25228 33328 25280 33380
rect 36452 33396 36504 33448
rect 31852 33328 31904 33380
rect 58164 33371 58216 33380
rect 58164 33337 58173 33371
rect 58173 33337 58207 33371
rect 58207 33337 58216 33371
rect 58164 33328 58216 33337
rect 4620 33260 4672 33312
rect 4896 33260 4948 33312
rect 24492 33260 24544 33312
rect 25136 33260 25188 33312
rect 31208 33260 31260 33312
rect 37280 33303 37332 33312
rect 37280 33269 37289 33303
rect 37289 33269 37323 33303
rect 37323 33269 37332 33303
rect 37280 33260 37332 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 6736 33056 6788 33108
rect 7472 33056 7524 33108
rect 9036 33056 9088 33108
rect 17408 33056 17460 33108
rect 19156 33056 19208 33108
rect 4804 32988 4856 33040
rect 7656 32988 7708 33040
rect 4620 32920 4672 32972
rect 5080 32920 5132 32972
rect 7012 32920 7064 32972
rect 6736 32852 6788 32904
rect 7380 32895 7432 32904
rect 7380 32861 7389 32895
rect 7389 32861 7423 32895
rect 7423 32861 7432 32895
rect 7380 32852 7432 32861
rect 10048 32920 10100 32972
rect 9864 32895 9916 32904
rect 9864 32861 9873 32895
rect 9873 32861 9907 32895
rect 9907 32861 9916 32895
rect 9864 32852 9916 32861
rect 9956 32852 10008 32904
rect 12808 32920 12860 32972
rect 16856 32988 16908 33040
rect 20352 33056 20404 33108
rect 22008 33056 22060 33108
rect 23664 33056 23716 33108
rect 23940 33056 23992 33108
rect 25136 33056 25188 33108
rect 27344 33056 27396 33108
rect 32036 33056 32088 33108
rect 35992 33056 36044 33108
rect 31116 33031 31168 33040
rect 31116 32997 31125 33031
rect 31125 32997 31159 33031
rect 31159 32997 31168 33031
rect 31116 32988 31168 32997
rect 35348 32988 35400 33040
rect 35808 32988 35860 33040
rect 25228 32920 25280 32972
rect 34796 32920 34848 32972
rect 12992 32852 13044 32904
rect 16120 32852 16172 32904
rect 17592 32895 17644 32904
rect 17592 32861 17601 32895
rect 17601 32861 17635 32895
rect 17635 32861 17644 32895
rect 17592 32852 17644 32861
rect 20812 32852 20864 32904
rect 24492 32852 24544 32904
rect 30472 32852 30524 32904
rect 30564 32852 30616 32904
rect 32588 32852 32640 32904
rect 33048 32895 33100 32904
rect 33048 32861 33057 32895
rect 33057 32861 33091 32895
rect 33091 32861 33100 32895
rect 33048 32852 33100 32861
rect 33140 32852 33192 32904
rect 37280 32920 37332 32972
rect 38568 32920 38620 32972
rect 35900 32895 35952 32904
rect 35900 32861 35909 32895
rect 35909 32861 35943 32895
rect 35943 32861 35952 32895
rect 36084 32895 36136 32904
rect 35900 32852 35952 32861
rect 36084 32861 36093 32895
rect 36093 32861 36127 32895
rect 36127 32861 36136 32895
rect 36084 32852 36136 32861
rect 5172 32784 5224 32836
rect 7104 32784 7156 32836
rect 3792 32759 3844 32768
rect 3792 32725 3801 32759
rect 3801 32725 3835 32759
rect 3835 32725 3844 32759
rect 3792 32716 3844 32725
rect 6920 32716 6972 32768
rect 11980 32827 12032 32836
rect 11980 32793 11989 32827
rect 11989 32793 12023 32827
rect 12023 32793 12032 32827
rect 11980 32784 12032 32793
rect 12532 32784 12584 32836
rect 12624 32784 12676 32836
rect 13084 32759 13136 32768
rect 13084 32725 13093 32759
rect 13093 32725 13127 32759
rect 13127 32725 13136 32759
rect 13084 32716 13136 32725
rect 14556 32784 14608 32836
rect 21824 32784 21876 32836
rect 28540 32784 28592 32836
rect 15108 32716 15160 32768
rect 15476 32759 15528 32768
rect 15476 32725 15485 32759
rect 15485 32725 15519 32759
rect 15519 32725 15528 32759
rect 15476 32716 15528 32725
rect 15568 32716 15620 32768
rect 17776 32716 17828 32768
rect 21088 32716 21140 32768
rect 23572 32716 23624 32768
rect 27712 32716 27764 32768
rect 28724 32716 28776 32768
rect 31668 32716 31720 32768
rect 31944 32716 31996 32768
rect 32128 32716 32180 32768
rect 32864 32827 32916 32836
rect 32864 32793 32873 32827
rect 32873 32793 32907 32827
rect 32907 32793 32916 32827
rect 35072 32827 35124 32836
rect 32864 32784 32916 32793
rect 35072 32793 35081 32827
rect 35081 32793 35115 32827
rect 35115 32793 35124 32827
rect 35072 32784 35124 32793
rect 36268 32895 36320 32904
rect 36268 32861 36277 32895
rect 36277 32861 36311 32895
rect 36311 32861 36320 32895
rect 36268 32852 36320 32861
rect 38200 32895 38252 32904
rect 38200 32861 38218 32895
rect 38218 32861 38252 32895
rect 38200 32852 38252 32861
rect 36452 32784 36504 32836
rect 35808 32716 35860 32768
rect 36544 32759 36596 32768
rect 36544 32725 36553 32759
rect 36553 32725 36587 32759
rect 36587 32725 36596 32759
rect 36544 32716 36596 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 5172 32512 5224 32564
rect 6092 32512 6144 32564
rect 6460 32512 6512 32564
rect 7288 32512 7340 32564
rect 2136 32308 2188 32360
rect 6184 32444 6236 32496
rect 3792 32376 3844 32428
rect 5540 32376 5592 32428
rect 7472 32444 7524 32496
rect 5448 32308 5500 32360
rect 6460 32308 6512 32360
rect 4712 32240 4764 32292
rect 6552 32240 6604 32292
rect 6460 32172 6512 32224
rect 6644 32172 6696 32224
rect 6920 32376 6972 32428
rect 7012 32419 7064 32428
rect 7012 32385 7021 32419
rect 7021 32385 7055 32419
rect 7055 32385 7064 32419
rect 9956 32487 10008 32496
rect 9956 32453 9965 32487
rect 9965 32453 9999 32487
rect 9999 32453 10008 32487
rect 9956 32444 10008 32453
rect 11980 32512 12032 32564
rect 14556 32487 14608 32496
rect 14556 32453 14565 32487
rect 14565 32453 14599 32487
rect 14599 32453 14608 32487
rect 14556 32444 14608 32453
rect 15016 32487 15068 32496
rect 15016 32453 15025 32487
rect 15025 32453 15059 32487
rect 15059 32453 15068 32487
rect 15016 32444 15068 32453
rect 15476 32444 15528 32496
rect 7012 32376 7064 32385
rect 9128 32376 9180 32428
rect 9404 32376 9456 32428
rect 12716 32419 12768 32428
rect 12716 32385 12734 32419
rect 12734 32385 12768 32419
rect 12716 32376 12768 32385
rect 12992 32419 13044 32428
rect 12992 32385 13001 32419
rect 13001 32385 13035 32419
rect 13035 32385 13044 32419
rect 12992 32376 13044 32385
rect 13912 32419 13964 32428
rect 13912 32385 13921 32419
rect 13921 32385 13955 32419
rect 13955 32385 13964 32419
rect 13912 32376 13964 32385
rect 7288 32308 7340 32360
rect 14188 32419 14240 32428
rect 14188 32385 14200 32419
rect 14200 32385 14234 32419
rect 14234 32385 14240 32419
rect 14188 32376 14240 32385
rect 14372 32376 14424 32428
rect 15108 32376 15160 32428
rect 17500 32444 17552 32496
rect 21088 32487 21140 32496
rect 21088 32453 21097 32487
rect 21097 32453 21131 32487
rect 21131 32453 21140 32487
rect 21088 32444 21140 32453
rect 21640 32444 21692 32496
rect 21824 32487 21876 32496
rect 21824 32453 21833 32487
rect 21833 32453 21867 32487
rect 21867 32453 21876 32487
rect 21824 32444 21876 32453
rect 20904 32419 20956 32428
rect 16580 32308 16632 32360
rect 16948 32240 17000 32292
rect 20904 32385 20913 32419
rect 20913 32385 20947 32419
rect 20947 32385 20956 32419
rect 20904 32376 20956 32385
rect 22008 32376 22060 32428
rect 22192 32419 22244 32428
rect 22192 32385 22201 32419
rect 22201 32385 22235 32419
rect 22235 32385 22244 32419
rect 22192 32376 22244 32385
rect 22468 32419 22520 32428
rect 22468 32385 22477 32419
rect 22477 32385 22511 32419
rect 22511 32385 22520 32419
rect 22468 32376 22520 32385
rect 22928 32419 22980 32428
rect 22928 32385 22937 32419
rect 22937 32385 22971 32419
rect 22971 32385 22980 32419
rect 22928 32376 22980 32385
rect 17408 32240 17460 32292
rect 23572 32308 23624 32360
rect 23112 32283 23164 32292
rect 23112 32249 23121 32283
rect 23121 32249 23155 32283
rect 23155 32249 23164 32283
rect 23112 32240 23164 32249
rect 24492 32512 24544 32564
rect 28540 32512 28592 32564
rect 28816 32512 28868 32564
rect 31944 32512 31996 32564
rect 24676 32444 24728 32496
rect 24860 32444 24912 32496
rect 27344 32487 27396 32496
rect 27344 32453 27353 32487
rect 27353 32453 27387 32487
rect 27387 32453 27396 32487
rect 27344 32444 27396 32453
rect 33140 32444 33192 32496
rect 35072 32444 35124 32496
rect 35348 32444 35400 32496
rect 36084 32512 36136 32564
rect 36268 32444 36320 32496
rect 23848 32308 23900 32360
rect 25228 32419 25280 32428
rect 25228 32385 25237 32419
rect 25237 32385 25271 32419
rect 25271 32385 25280 32419
rect 25228 32376 25280 32385
rect 28264 32376 28316 32428
rect 31760 32376 31812 32428
rect 31944 32376 31996 32428
rect 32588 32419 32640 32428
rect 32588 32385 32597 32419
rect 32597 32385 32631 32419
rect 32631 32385 32640 32419
rect 32588 32376 32640 32385
rect 32772 32419 32824 32428
rect 32772 32385 32781 32419
rect 32781 32385 32815 32419
rect 32815 32385 32824 32419
rect 32772 32376 32824 32385
rect 34520 32376 34572 32428
rect 36084 32376 36136 32428
rect 24860 32308 24912 32360
rect 28540 32240 28592 32292
rect 10140 32215 10192 32224
rect 10140 32181 10149 32215
rect 10149 32181 10183 32215
rect 10183 32181 10192 32215
rect 10140 32172 10192 32181
rect 17684 32172 17736 32224
rect 17776 32172 17828 32224
rect 23940 32172 23992 32224
rect 24768 32215 24820 32224
rect 24768 32181 24777 32215
rect 24777 32181 24811 32215
rect 24811 32181 24820 32215
rect 24768 32172 24820 32181
rect 26792 32172 26844 32224
rect 32220 32172 32272 32224
rect 58164 32215 58216 32224
rect 58164 32181 58173 32215
rect 58173 32181 58207 32215
rect 58207 32181 58216 32215
rect 58164 32172 58216 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 6828 31968 6880 32020
rect 7380 31968 7432 32020
rect 9956 31968 10008 32020
rect 12716 31968 12768 32020
rect 16764 31968 16816 32020
rect 17500 32011 17552 32020
rect 17500 31977 17509 32011
rect 17509 31977 17543 32011
rect 17543 31977 17552 32011
rect 17500 31968 17552 31977
rect 20904 31968 20956 32020
rect 8944 31875 8996 31884
rect 8944 31841 8953 31875
rect 8953 31841 8987 31875
rect 8987 31841 8996 31875
rect 8944 31832 8996 31841
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 1952 31764 2004 31816
rect 5724 31807 5776 31816
rect 5724 31773 5733 31807
rect 5733 31773 5767 31807
rect 5767 31773 5776 31807
rect 5724 31764 5776 31773
rect 11060 31764 11112 31816
rect 12716 31764 12768 31816
rect 12992 31807 13044 31816
rect 12992 31773 13001 31807
rect 13001 31773 13035 31807
rect 13035 31773 13044 31807
rect 12992 31764 13044 31773
rect 13176 31807 13228 31816
rect 13176 31773 13185 31807
rect 13185 31773 13219 31807
rect 13219 31773 13228 31807
rect 13176 31764 13228 31773
rect 16672 31764 16724 31816
rect 16764 31764 16816 31816
rect 22928 31968 22980 32020
rect 27160 31968 27212 32020
rect 27712 32011 27764 32020
rect 27712 31977 27721 32011
rect 27721 31977 27755 32011
rect 27755 31977 27764 32011
rect 27712 31968 27764 31977
rect 28264 32011 28316 32020
rect 28264 31977 28273 32011
rect 28273 31977 28307 32011
rect 28307 31977 28316 32011
rect 28264 31968 28316 31977
rect 28540 31968 28592 32020
rect 30380 31968 30432 32020
rect 31668 31968 31720 32020
rect 35992 32011 36044 32020
rect 35992 31977 36001 32011
rect 36001 31977 36035 32011
rect 36035 31977 36044 32011
rect 35992 31968 36044 31977
rect 36084 31968 36136 32020
rect 31300 31900 31352 31952
rect 31760 31900 31812 31952
rect 22836 31832 22888 31884
rect 26240 31832 26292 31884
rect 26792 31832 26844 31884
rect 2596 31696 2648 31748
rect 9680 31696 9732 31748
rect 3884 31628 3936 31680
rect 16580 31696 16632 31748
rect 16856 31696 16908 31748
rect 19432 31764 19484 31816
rect 24768 31764 24820 31816
rect 26516 31807 26568 31816
rect 26516 31773 26525 31807
rect 26525 31773 26559 31807
rect 26559 31773 26568 31807
rect 26516 31764 26568 31773
rect 27712 31764 27764 31816
rect 30104 31832 30156 31884
rect 28724 31807 28776 31816
rect 28724 31773 28733 31807
rect 28733 31773 28767 31807
rect 28767 31773 28776 31807
rect 28724 31764 28776 31773
rect 17592 31696 17644 31748
rect 22928 31696 22980 31748
rect 28448 31696 28500 31748
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 31484 31764 31536 31773
rect 31944 31764 31996 31816
rect 32312 31764 32364 31816
rect 32588 31832 32640 31884
rect 32680 31832 32732 31884
rect 32496 31807 32548 31816
rect 32496 31773 32505 31807
rect 32505 31773 32539 31807
rect 32539 31773 32548 31807
rect 32496 31764 32548 31773
rect 35808 31807 35860 31816
rect 35808 31773 35817 31807
rect 35817 31773 35851 31807
rect 35851 31773 35860 31807
rect 35808 31764 35860 31773
rect 36544 31764 36596 31816
rect 38568 31764 38620 31816
rect 29828 31696 29880 31748
rect 32680 31696 32732 31748
rect 35348 31696 35400 31748
rect 13268 31628 13320 31680
rect 14372 31628 14424 31680
rect 17316 31628 17368 31680
rect 18328 31671 18380 31680
rect 18328 31637 18337 31671
rect 18337 31637 18371 31671
rect 18371 31637 18380 31671
rect 18328 31628 18380 31637
rect 24400 31671 24452 31680
rect 24400 31637 24409 31671
rect 24409 31637 24443 31671
rect 24443 31637 24452 31671
rect 24400 31628 24452 31637
rect 26516 31628 26568 31680
rect 31116 31628 31168 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 2964 31424 3016 31476
rect 3424 31424 3476 31476
rect 3792 31424 3844 31476
rect 4068 31424 4120 31476
rect 9680 31467 9732 31476
rect 9680 31433 9689 31467
rect 9689 31433 9723 31467
rect 9723 31433 9732 31467
rect 9680 31424 9732 31433
rect 13176 31424 13228 31476
rect 16672 31467 16724 31476
rect 16672 31433 16681 31467
rect 16681 31433 16715 31467
rect 16715 31433 16724 31467
rect 16672 31424 16724 31433
rect 6460 31356 6512 31408
rect 12716 31356 12768 31408
rect 2136 31331 2188 31340
rect 2136 31297 2145 31331
rect 2145 31297 2179 31331
rect 2179 31297 2188 31331
rect 2136 31288 2188 31297
rect 2688 31288 2740 31340
rect 9864 31288 9916 31340
rect 10029 31331 10081 31340
rect 10029 31297 10054 31331
rect 10054 31297 10081 31331
rect 10029 31288 10081 31297
rect 10140 31331 10192 31340
rect 10140 31297 10154 31331
rect 10154 31297 10188 31331
rect 10188 31297 10192 31331
rect 10140 31288 10192 31297
rect 6184 31220 6236 31272
rect 10232 31220 10284 31272
rect 10508 31288 10560 31340
rect 14372 31288 14424 31340
rect 17132 31424 17184 31476
rect 21916 31424 21968 31476
rect 23848 31424 23900 31476
rect 18328 31356 18380 31408
rect 17960 31288 18012 31340
rect 19064 31288 19116 31340
rect 22192 31356 22244 31408
rect 25504 31424 25556 31476
rect 26516 31424 26568 31476
rect 29000 31424 29052 31476
rect 30380 31424 30432 31476
rect 9864 31152 9916 31204
rect 10508 31152 10560 31204
rect 11704 31152 11756 31204
rect 14188 31152 14240 31204
rect 22928 31288 22980 31340
rect 24676 31356 24728 31408
rect 36084 31356 36136 31408
rect 24400 31331 24452 31340
rect 24400 31297 24409 31331
rect 24409 31297 24443 31331
rect 24443 31297 24452 31331
rect 24400 31288 24452 31297
rect 28540 31288 28592 31340
rect 24952 31220 25004 31272
rect 26056 31220 26108 31272
rect 28724 31220 28776 31272
rect 29276 31288 29328 31340
rect 32312 31288 32364 31340
rect 32680 31331 32732 31340
rect 32680 31297 32689 31331
rect 32689 31297 32723 31331
rect 32723 31297 32732 31331
rect 32680 31288 32732 31297
rect 33232 31288 33284 31340
rect 25136 31152 25188 31204
rect 25688 31152 25740 31204
rect 3516 31127 3568 31136
rect 3516 31093 3525 31127
rect 3525 31093 3559 31127
rect 3559 31093 3568 31127
rect 3516 31084 3568 31093
rect 4068 31127 4120 31136
rect 4068 31093 4077 31127
rect 4077 31093 4111 31127
rect 4111 31093 4120 31127
rect 4068 31084 4120 31093
rect 7104 31084 7156 31136
rect 7748 31127 7800 31136
rect 7748 31093 7757 31127
rect 7757 31093 7791 31127
rect 7791 31093 7800 31127
rect 7748 31084 7800 31093
rect 12256 31127 12308 31136
rect 12256 31093 12265 31127
rect 12265 31093 12299 31127
rect 12299 31093 12308 31127
rect 12256 31084 12308 31093
rect 12440 31084 12492 31136
rect 17408 31084 17460 31136
rect 19340 31127 19392 31136
rect 19340 31093 19349 31127
rect 19349 31093 19383 31127
rect 19383 31093 19392 31127
rect 19340 31084 19392 31093
rect 23848 31084 23900 31136
rect 24032 31084 24084 31136
rect 29000 31084 29052 31136
rect 29828 31084 29880 31136
rect 32864 31084 32916 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2596 30923 2648 30932
rect 2596 30889 2605 30923
rect 2605 30889 2639 30923
rect 2639 30889 2648 30923
rect 2596 30880 2648 30889
rect 7104 30880 7156 30932
rect 8208 30880 8260 30932
rect 24676 30880 24728 30932
rect 26056 30880 26108 30932
rect 33692 30880 33744 30932
rect 4068 30812 4120 30864
rect 16120 30744 16172 30796
rect 17776 30744 17828 30796
rect 24400 30812 24452 30864
rect 3332 30676 3384 30728
rect 3884 30676 3936 30728
rect 4620 30676 4672 30728
rect 5448 30676 5500 30728
rect 6184 30719 6236 30728
rect 6184 30685 6193 30719
rect 6193 30685 6227 30719
rect 6227 30685 6236 30719
rect 6184 30676 6236 30685
rect 6828 30676 6880 30728
rect 9680 30719 9732 30728
rect 9680 30685 9689 30719
rect 9689 30685 9723 30719
rect 9723 30685 9732 30719
rect 9680 30676 9732 30685
rect 10784 30676 10836 30728
rect 6460 30651 6512 30660
rect 6460 30617 6494 30651
rect 6494 30617 6512 30651
rect 6460 30608 6512 30617
rect 12256 30608 12308 30660
rect 12716 30608 12768 30660
rect 13360 30651 13412 30660
rect 13360 30617 13369 30651
rect 13369 30617 13403 30651
rect 13403 30617 13412 30651
rect 15200 30651 15252 30660
rect 13360 30608 13412 30617
rect 2964 30540 3016 30592
rect 9404 30540 9456 30592
rect 11060 30540 11112 30592
rect 12992 30540 13044 30592
rect 13728 30540 13780 30592
rect 15200 30617 15218 30651
rect 15218 30617 15252 30651
rect 15200 30608 15252 30617
rect 20904 30676 20956 30728
rect 21640 30719 21692 30728
rect 21640 30685 21649 30719
rect 21649 30685 21683 30719
rect 21683 30685 21692 30719
rect 21640 30676 21692 30685
rect 21824 30676 21876 30728
rect 24952 30744 25004 30796
rect 30932 30744 30984 30796
rect 22560 30676 22612 30728
rect 23664 30719 23716 30728
rect 23664 30685 23673 30719
rect 23673 30685 23707 30719
rect 23707 30685 23716 30719
rect 23664 30676 23716 30685
rect 24492 30719 24544 30728
rect 24492 30685 24501 30719
rect 24501 30685 24535 30719
rect 24535 30685 24544 30719
rect 24492 30676 24544 30685
rect 24676 30719 24728 30728
rect 24676 30685 24685 30719
rect 24685 30685 24719 30719
rect 24719 30685 24728 30719
rect 24676 30676 24728 30685
rect 15844 30608 15896 30660
rect 19984 30608 20036 30660
rect 22008 30608 22060 30660
rect 25228 30676 25280 30728
rect 20628 30583 20680 30592
rect 20628 30549 20637 30583
rect 20637 30549 20671 30583
rect 20671 30549 20680 30583
rect 20628 30540 20680 30549
rect 20996 30540 21048 30592
rect 24584 30540 24636 30592
rect 25596 30583 25648 30592
rect 25596 30549 25605 30583
rect 25605 30549 25639 30583
rect 25639 30549 25648 30583
rect 25596 30540 25648 30549
rect 26884 30676 26936 30728
rect 28540 30719 28592 30728
rect 28540 30685 28549 30719
rect 28549 30685 28583 30719
rect 28583 30685 28592 30719
rect 28540 30676 28592 30685
rect 28908 30719 28960 30728
rect 28908 30685 28917 30719
rect 28917 30685 28951 30719
rect 28951 30685 28960 30719
rect 28908 30676 28960 30685
rect 30380 30676 30432 30728
rect 31208 30719 31260 30728
rect 31208 30685 31217 30719
rect 31217 30685 31251 30719
rect 31251 30685 31260 30719
rect 31208 30676 31260 30685
rect 32312 30744 32364 30796
rect 28172 30608 28224 30660
rect 28724 30651 28776 30660
rect 28724 30617 28733 30651
rect 28733 30617 28767 30651
rect 28767 30617 28776 30651
rect 28724 30608 28776 30617
rect 31484 30676 31536 30728
rect 32496 30676 32548 30728
rect 34520 30676 34572 30728
rect 38568 30676 38620 30728
rect 58164 30719 58216 30728
rect 58164 30685 58173 30719
rect 58173 30685 58207 30719
rect 58207 30685 58216 30719
rect 58164 30676 58216 30685
rect 31576 30608 31628 30660
rect 33968 30651 34020 30660
rect 33968 30617 33977 30651
rect 33977 30617 34011 30651
rect 34011 30617 34020 30651
rect 33968 30608 34020 30617
rect 31852 30540 31904 30592
rect 34336 30540 34388 30592
rect 35348 30540 35400 30592
rect 35900 30608 35952 30660
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 2688 30379 2740 30388
rect 2688 30345 2697 30379
rect 2697 30345 2731 30379
rect 2731 30345 2740 30379
rect 2688 30336 2740 30345
rect 2964 30336 3016 30388
rect 3240 30336 3292 30388
rect 6460 30336 6512 30388
rect 10784 30379 10836 30388
rect 10784 30345 10793 30379
rect 10793 30345 10827 30379
rect 10827 30345 10836 30379
rect 10784 30336 10836 30345
rect 13268 30336 13320 30388
rect 15844 30379 15896 30388
rect 15844 30345 15853 30379
rect 15853 30345 15887 30379
rect 15887 30345 15896 30379
rect 15844 30336 15896 30345
rect 3976 30268 4028 30320
rect 12624 30268 12676 30320
rect 3332 30243 3384 30252
rect 3332 30209 3341 30243
rect 3341 30209 3375 30243
rect 3375 30209 3384 30243
rect 3332 30200 3384 30209
rect 3884 30200 3936 30252
rect 5080 30200 5132 30252
rect 5632 30200 5684 30252
rect 6368 30200 6420 30252
rect 4988 30132 5040 30184
rect 6920 30200 6972 30252
rect 7564 30200 7616 30252
rect 7472 30132 7524 30184
rect 3424 30064 3476 30116
rect 10140 30243 10192 30252
rect 10140 30209 10154 30243
rect 10154 30209 10188 30243
rect 10188 30209 10192 30243
rect 10140 30200 10192 30209
rect 12164 30243 12216 30252
rect 10232 30132 10284 30184
rect 12164 30209 12173 30243
rect 12173 30209 12207 30243
rect 12207 30209 12216 30243
rect 12164 30200 12216 30209
rect 12992 30243 13044 30252
rect 12992 30209 13001 30243
rect 13001 30209 13035 30243
rect 13035 30209 13044 30243
rect 12992 30200 13044 30209
rect 13176 30200 13228 30252
rect 13728 30243 13780 30252
rect 13728 30209 13737 30243
rect 13737 30209 13771 30243
rect 13771 30209 13780 30243
rect 13728 30200 13780 30209
rect 15200 30268 15252 30320
rect 16764 30311 16816 30320
rect 16764 30277 16773 30311
rect 16773 30277 16807 30311
rect 16807 30277 16816 30311
rect 16764 30268 16816 30277
rect 20628 30268 20680 30320
rect 22008 30268 22060 30320
rect 25044 30268 25096 30320
rect 26056 30268 26108 30320
rect 30932 30336 30984 30388
rect 31208 30379 31260 30388
rect 31208 30345 31217 30379
rect 31217 30345 31251 30379
rect 31251 30345 31260 30379
rect 31208 30336 31260 30345
rect 28632 30311 28684 30320
rect 28632 30277 28641 30311
rect 28641 30277 28675 30311
rect 28675 30277 28684 30311
rect 28632 30268 28684 30277
rect 28724 30311 28776 30320
rect 28724 30277 28733 30311
rect 28733 30277 28767 30311
rect 28767 30277 28776 30311
rect 28724 30268 28776 30277
rect 30380 30268 30432 30320
rect 12440 30132 12492 30184
rect 13452 30132 13504 30184
rect 4804 29996 4856 30048
rect 7564 30039 7616 30048
rect 7564 30005 7573 30039
rect 7573 30005 7607 30039
rect 7607 30005 7616 30039
rect 7564 29996 7616 30005
rect 9496 29996 9548 30048
rect 10048 30064 10100 30116
rect 10784 30064 10836 30116
rect 14372 30064 14424 30116
rect 12900 29996 12952 30048
rect 15292 30200 15344 30252
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 19432 30200 19484 30252
rect 19892 30243 19944 30252
rect 19892 30209 19901 30243
rect 19901 30209 19935 30243
rect 19935 30209 19944 30243
rect 19892 30200 19944 30209
rect 22100 30243 22152 30252
rect 22100 30209 22109 30243
rect 22109 30209 22143 30243
rect 22143 30209 22152 30243
rect 22100 30200 22152 30209
rect 16672 30132 16724 30184
rect 20904 30132 20956 30184
rect 23112 30200 23164 30252
rect 24860 30200 24912 30252
rect 28540 30243 28592 30252
rect 28540 30209 28549 30243
rect 28549 30209 28583 30243
rect 28583 30209 28592 30243
rect 28540 30200 28592 30209
rect 24584 30132 24636 30184
rect 28816 30200 28868 30252
rect 29920 30243 29972 30252
rect 29920 30209 29929 30243
rect 29929 30209 29963 30243
rect 29963 30209 29972 30243
rect 32956 30268 33008 30320
rect 33692 30311 33744 30320
rect 33692 30277 33701 30311
rect 33701 30277 33735 30311
rect 33735 30277 33744 30311
rect 33692 30268 33744 30277
rect 34244 30268 34296 30320
rect 29920 30200 29972 30209
rect 31576 30243 31628 30252
rect 31576 30209 31585 30243
rect 31585 30209 31619 30243
rect 31619 30209 31628 30243
rect 31576 30200 31628 30209
rect 32680 30243 32732 30252
rect 32680 30209 32689 30243
rect 32689 30209 32723 30243
rect 32723 30209 32732 30243
rect 32680 30200 32732 30209
rect 33600 30200 33652 30252
rect 34336 30243 34388 30252
rect 34336 30209 34345 30243
rect 34345 30209 34379 30243
rect 34379 30209 34388 30243
rect 34336 30200 34388 30209
rect 35900 30268 35952 30320
rect 14832 29996 14884 30048
rect 19432 29996 19484 30048
rect 22652 30039 22704 30048
rect 22652 30005 22661 30039
rect 22661 30005 22695 30039
rect 22695 30005 22704 30039
rect 22652 29996 22704 30005
rect 29828 30064 29880 30116
rect 29552 29996 29604 30048
rect 33048 30132 33100 30184
rect 30932 30064 30984 30116
rect 35992 30200 36044 30252
rect 36452 30200 36504 30252
rect 37464 30243 37516 30252
rect 31760 29996 31812 30048
rect 35348 30132 35400 30184
rect 37464 30209 37473 30243
rect 37473 30209 37507 30243
rect 37507 30209 37516 30243
rect 37464 30200 37516 30209
rect 35716 29996 35768 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3240 29835 3292 29844
rect 3240 29801 3249 29835
rect 3249 29801 3283 29835
rect 3283 29801 3292 29835
rect 3240 29792 3292 29801
rect 6920 29835 6972 29844
rect 6920 29801 6929 29835
rect 6929 29801 6963 29835
rect 6963 29801 6972 29835
rect 6920 29792 6972 29801
rect 2780 29588 2832 29640
rect 4620 29724 4672 29776
rect 3148 29656 3200 29708
rect 3516 29588 3568 29640
rect 5080 29588 5132 29640
rect 7104 29588 7156 29640
rect 13176 29792 13228 29844
rect 19984 29792 20036 29844
rect 29552 29835 29604 29844
rect 15016 29724 15068 29776
rect 15752 29724 15804 29776
rect 21180 29724 21232 29776
rect 21824 29724 21876 29776
rect 8944 29656 8996 29708
rect 12532 29656 12584 29708
rect 12900 29656 12952 29708
rect 9496 29631 9548 29640
rect 9496 29597 9530 29631
rect 9530 29597 9548 29631
rect 9496 29588 9548 29597
rect 11152 29588 11204 29640
rect 12808 29631 12860 29640
rect 4988 29520 5040 29572
rect 7012 29520 7064 29572
rect 4712 29452 4764 29504
rect 9956 29452 10008 29504
rect 12808 29597 12817 29631
rect 12817 29597 12851 29631
rect 12851 29597 12860 29631
rect 12808 29588 12860 29597
rect 16764 29588 16816 29640
rect 17592 29588 17644 29640
rect 19432 29631 19484 29640
rect 19432 29597 19441 29631
rect 19441 29597 19475 29631
rect 19475 29597 19484 29631
rect 19432 29588 19484 29597
rect 20628 29656 20680 29708
rect 13360 29520 13412 29572
rect 15936 29563 15988 29572
rect 15936 29529 15945 29563
rect 15945 29529 15979 29563
rect 15979 29529 15988 29563
rect 15936 29520 15988 29529
rect 14740 29452 14792 29504
rect 16028 29452 16080 29504
rect 16672 29495 16724 29504
rect 16672 29461 16681 29495
rect 16681 29461 16715 29495
rect 16715 29461 16724 29495
rect 16672 29452 16724 29461
rect 18420 29452 18472 29504
rect 19340 29520 19392 29572
rect 20904 29588 20956 29640
rect 29552 29801 29561 29835
rect 29561 29801 29595 29835
rect 29595 29801 29604 29835
rect 29552 29792 29604 29801
rect 32956 29835 33008 29844
rect 32956 29801 32965 29835
rect 32965 29801 32999 29835
rect 32999 29801 33008 29835
rect 32956 29792 33008 29801
rect 31484 29724 31536 29776
rect 21456 29588 21508 29640
rect 21088 29563 21140 29572
rect 21088 29529 21097 29563
rect 21097 29529 21131 29563
rect 21131 29529 21140 29563
rect 21088 29520 21140 29529
rect 20720 29452 20772 29504
rect 22008 29520 22060 29572
rect 24492 29588 24544 29640
rect 24952 29631 25004 29640
rect 24952 29597 24961 29631
rect 24961 29597 24995 29631
rect 24995 29597 25004 29631
rect 24952 29588 25004 29597
rect 24584 29520 24636 29572
rect 31576 29631 31628 29640
rect 31576 29597 31585 29631
rect 31585 29597 31619 29631
rect 31619 29597 31628 29631
rect 31576 29588 31628 29597
rect 31852 29631 31904 29640
rect 31852 29597 31886 29631
rect 31886 29597 31904 29631
rect 31852 29588 31904 29597
rect 35440 29588 35492 29640
rect 35716 29631 35768 29640
rect 35716 29597 35725 29631
rect 35725 29597 35759 29631
rect 35759 29597 35768 29631
rect 35716 29588 35768 29597
rect 35992 29656 36044 29708
rect 35900 29631 35952 29640
rect 35900 29597 35909 29631
rect 35909 29597 35943 29631
rect 35943 29597 35952 29631
rect 35900 29588 35952 29597
rect 38568 29588 38620 29640
rect 58164 29631 58216 29640
rect 58164 29597 58173 29631
rect 58173 29597 58207 29631
rect 58207 29597 58216 29631
rect 58164 29588 58216 29597
rect 22468 29452 22520 29504
rect 25872 29495 25924 29504
rect 25872 29461 25881 29495
rect 25881 29461 25915 29495
rect 25915 29461 25924 29495
rect 25872 29452 25924 29461
rect 26792 29520 26844 29572
rect 33876 29520 33928 29572
rect 30380 29495 30432 29504
rect 30380 29461 30389 29495
rect 30389 29461 30423 29495
rect 30423 29461 30432 29495
rect 30380 29452 30432 29461
rect 34612 29452 34664 29504
rect 35532 29452 35584 29504
rect 35808 29452 35860 29504
rect 37464 29452 37516 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 11704 29112 11756 29164
rect 12808 29112 12860 29164
rect 14648 29112 14700 29164
rect 14832 29112 14884 29164
rect 15752 29155 15804 29164
rect 15752 29121 15761 29155
rect 15761 29121 15795 29155
rect 15795 29121 15804 29155
rect 15752 29112 15804 29121
rect 17132 29180 17184 29232
rect 17316 29223 17368 29232
rect 17316 29189 17325 29223
rect 17325 29189 17359 29223
rect 17359 29189 17368 29223
rect 17316 29180 17368 29189
rect 18144 29180 18196 29232
rect 24952 29248 25004 29300
rect 31760 29248 31812 29300
rect 34796 29248 34848 29300
rect 20628 29223 20680 29232
rect 7472 29044 7524 29096
rect 9680 29044 9732 29096
rect 11428 29044 11480 29096
rect 15108 29044 15160 29096
rect 16028 29112 16080 29164
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 17776 29155 17828 29164
rect 16120 29112 16172 29121
rect 17776 29121 17785 29155
rect 17785 29121 17819 29155
rect 17819 29121 17828 29155
rect 17776 29112 17828 29121
rect 17868 29112 17920 29164
rect 19984 29155 20036 29164
rect 19984 29121 19993 29155
rect 19993 29121 20027 29155
rect 20027 29121 20036 29155
rect 19984 29112 20036 29121
rect 20628 29189 20637 29223
rect 20637 29189 20671 29223
rect 20671 29189 20680 29223
rect 20628 29180 20680 29189
rect 21088 29180 21140 29232
rect 11152 28976 11204 29028
rect 11888 28976 11940 29028
rect 12440 28976 12492 29028
rect 17132 28976 17184 29028
rect 20904 29112 20956 29164
rect 23664 29112 23716 29164
rect 24768 29155 24820 29164
rect 24768 29121 24777 29155
rect 24777 29121 24811 29155
rect 24811 29121 24820 29155
rect 24768 29112 24820 29121
rect 25872 29180 25924 29232
rect 33876 29223 33928 29232
rect 33876 29189 33885 29223
rect 33885 29189 33919 29223
rect 33919 29189 33928 29223
rect 33876 29180 33928 29189
rect 25504 29112 25556 29164
rect 29828 29155 29880 29164
rect 29828 29121 29837 29155
rect 29837 29121 29871 29155
rect 29871 29121 29880 29155
rect 29828 29112 29880 29121
rect 23388 29044 23440 29096
rect 30380 29112 30432 29164
rect 32496 29112 32548 29164
rect 33048 29044 33100 29096
rect 34060 29112 34112 29164
rect 34980 29112 35032 29164
rect 35440 29155 35492 29164
rect 35440 29121 35449 29155
rect 35449 29121 35483 29155
rect 35483 29121 35492 29155
rect 35440 29112 35492 29121
rect 35624 29155 35676 29164
rect 35624 29121 35633 29155
rect 35633 29121 35667 29155
rect 35667 29121 35676 29155
rect 35624 29112 35676 29121
rect 35992 29180 36044 29232
rect 38568 29112 38620 29164
rect 25596 28976 25648 29028
rect 25780 29019 25832 29028
rect 25780 28985 25789 29019
rect 25789 28985 25823 29019
rect 25823 28985 25832 29019
rect 25780 28976 25832 28985
rect 33784 28976 33836 29028
rect 34244 28976 34296 29028
rect 35440 28976 35492 29028
rect 35900 28976 35952 29028
rect 14372 28951 14424 28960
rect 14372 28917 14381 28951
rect 14381 28917 14415 28951
rect 14415 28917 14424 28951
rect 14372 28908 14424 28917
rect 15476 28951 15528 28960
rect 15476 28917 15485 28951
rect 15485 28917 15519 28951
rect 15519 28917 15528 28951
rect 15476 28908 15528 28917
rect 19616 28951 19668 28960
rect 19616 28917 19625 28951
rect 19625 28917 19659 28951
rect 19659 28917 19668 28951
rect 19616 28908 19668 28917
rect 20536 28908 20588 28960
rect 30104 28908 30156 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 10140 28747 10192 28756
rect 10140 28713 10149 28747
rect 10149 28713 10183 28747
rect 10183 28713 10192 28747
rect 10140 28704 10192 28713
rect 12900 28704 12952 28756
rect 13820 28704 13872 28756
rect 15016 28704 15068 28756
rect 17868 28747 17920 28756
rect 17868 28713 17877 28747
rect 17877 28713 17911 28747
rect 17911 28713 17920 28747
rect 17868 28704 17920 28713
rect 10048 28636 10100 28688
rect 16212 28636 16264 28688
rect 23388 28704 23440 28756
rect 24676 28747 24728 28756
rect 24676 28713 24685 28747
rect 24685 28713 24719 28747
rect 24719 28713 24728 28747
rect 24676 28704 24728 28713
rect 25504 28747 25556 28756
rect 25504 28713 25513 28747
rect 25513 28713 25547 28747
rect 25547 28713 25556 28747
rect 25504 28704 25556 28713
rect 29552 28704 29604 28756
rect 30564 28704 30616 28756
rect 2780 28543 2832 28552
rect 2780 28509 2789 28543
rect 2789 28509 2823 28543
rect 2823 28509 2832 28543
rect 2780 28500 2832 28509
rect 3700 28500 3752 28552
rect 4988 28568 5040 28620
rect 5080 28543 5132 28552
rect 5080 28509 5089 28543
rect 5089 28509 5123 28543
rect 5123 28509 5132 28543
rect 9680 28568 9732 28620
rect 5080 28500 5132 28509
rect 5356 28432 5408 28484
rect 6000 28432 6052 28484
rect 7012 28432 7064 28484
rect 8208 28432 8260 28484
rect 9312 28543 9364 28552
rect 9312 28509 9321 28543
rect 9321 28509 9355 28543
rect 9355 28509 9364 28543
rect 9312 28500 9364 28509
rect 9404 28500 9456 28552
rect 9956 28543 10008 28552
rect 9956 28509 9965 28543
rect 9965 28509 9999 28543
rect 9999 28509 10008 28543
rect 9956 28500 10008 28509
rect 11428 28543 11480 28552
rect 11428 28509 11437 28543
rect 11437 28509 11471 28543
rect 11471 28509 11480 28543
rect 11428 28500 11480 28509
rect 12164 28568 12216 28620
rect 14372 28568 14424 28620
rect 14924 28568 14976 28620
rect 18420 28636 18472 28688
rect 20812 28636 20864 28688
rect 21088 28636 21140 28688
rect 23940 28636 23992 28688
rect 25228 28636 25280 28688
rect 29276 28636 29328 28688
rect 13728 28432 13780 28484
rect 14832 28500 14884 28552
rect 15476 28543 15528 28552
rect 15476 28509 15510 28543
rect 15510 28509 15528 28543
rect 15476 28500 15528 28509
rect 17040 28500 17092 28552
rect 17592 28500 17644 28552
rect 18144 28543 18196 28552
rect 15016 28432 15068 28484
rect 17132 28475 17184 28484
rect 17132 28441 17141 28475
rect 17141 28441 17175 28475
rect 17175 28441 17184 28475
rect 17132 28432 17184 28441
rect 18144 28509 18153 28543
rect 18153 28509 18187 28543
rect 18187 28509 18196 28543
rect 18144 28500 18196 28509
rect 19616 28568 19668 28620
rect 22192 28568 22244 28620
rect 22836 28568 22888 28620
rect 23112 28543 23164 28552
rect 23112 28509 23121 28543
rect 23121 28509 23155 28543
rect 23155 28509 23164 28543
rect 23112 28500 23164 28509
rect 26516 28568 26568 28620
rect 32036 28704 32088 28756
rect 32588 28704 32640 28756
rect 33416 28636 33468 28688
rect 34612 28704 34664 28756
rect 35624 28704 35676 28756
rect 33692 28636 33744 28688
rect 34520 28636 34572 28688
rect 25596 28500 25648 28552
rect 29828 28500 29880 28552
rect 24676 28432 24728 28484
rect 3148 28407 3200 28416
rect 3148 28373 3157 28407
rect 3157 28373 3191 28407
rect 3191 28373 3200 28407
rect 3148 28364 3200 28373
rect 6736 28364 6788 28416
rect 7380 28364 7432 28416
rect 9312 28364 9364 28416
rect 9772 28364 9824 28416
rect 13452 28364 13504 28416
rect 14188 28364 14240 28416
rect 15200 28364 15252 28416
rect 15936 28364 15988 28416
rect 24216 28364 24268 28416
rect 32496 28500 32548 28552
rect 34704 28500 34756 28552
rect 35348 28543 35400 28552
rect 35348 28509 35357 28543
rect 35357 28509 35391 28543
rect 35391 28509 35400 28543
rect 35348 28500 35400 28509
rect 35900 28500 35952 28552
rect 30748 28475 30800 28484
rect 30748 28441 30757 28475
rect 30757 28441 30791 28475
rect 30791 28441 30800 28475
rect 30748 28432 30800 28441
rect 33784 28475 33836 28484
rect 33784 28441 33793 28475
rect 33793 28441 33827 28475
rect 33827 28441 33836 28475
rect 33784 28432 33836 28441
rect 33692 28364 33744 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 3700 28203 3752 28212
rect 3700 28169 3709 28203
rect 3709 28169 3743 28203
rect 3743 28169 3752 28203
rect 3700 28160 3752 28169
rect 8208 28203 8260 28212
rect 8208 28169 8217 28203
rect 8217 28169 8251 28203
rect 8251 28169 8260 28203
rect 8208 28160 8260 28169
rect 6552 28092 6604 28144
rect 2596 28067 2648 28076
rect 2596 28033 2630 28067
rect 2630 28033 2648 28067
rect 6828 28067 6880 28076
rect 2596 28024 2648 28033
rect 6828 28033 6837 28067
rect 6837 28033 6871 28067
rect 6871 28033 6880 28067
rect 6828 28024 6880 28033
rect 6920 28024 6972 28076
rect 2320 27999 2372 28008
rect 2320 27965 2329 27999
rect 2329 27965 2363 27999
rect 2363 27965 2372 27999
rect 2320 27956 2372 27965
rect 8668 28067 8720 28076
rect 8668 28033 8677 28067
rect 8677 28033 8711 28067
rect 8711 28033 8720 28067
rect 8668 28024 8720 28033
rect 8944 28067 8996 28076
rect 8944 28033 8953 28067
rect 8953 28033 8987 28067
rect 8987 28033 8996 28067
rect 8944 28024 8996 28033
rect 9128 28067 9180 28076
rect 9128 28033 9142 28067
rect 9142 28033 9176 28067
rect 9176 28033 9180 28067
rect 12532 28160 12584 28212
rect 9128 28024 9180 28033
rect 10692 28024 10744 28076
rect 13820 28160 13872 28212
rect 14188 28203 14240 28212
rect 14188 28169 14197 28203
rect 14197 28169 14231 28203
rect 14231 28169 14240 28203
rect 14188 28160 14240 28169
rect 16212 28160 16264 28212
rect 16948 28203 17000 28212
rect 16948 28169 16957 28203
rect 16957 28169 16991 28203
rect 16991 28169 17000 28203
rect 16948 28160 17000 28169
rect 17132 28160 17184 28212
rect 13084 28092 13136 28144
rect 15200 28135 15252 28144
rect 11704 27888 11756 27940
rect 13452 28067 13504 28076
rect 13452 28033 13461 28067
rect 13461 28033 13495 28067
rect 13495 28033 13504 28067
rect 13452 28024 13504 28033
rect 12532 27956 12584 28008
rect 14740 28024 14792 28076
rect 15200 28101 15209 28135
rect 15209 28101 15243 28135
rect 15243 28101 15252 28135
rect 15200 28092 15252 28101
rect 16120 28092 16172 28144
rect 17960 28092 18012 28144
rect 23848 28160 23900 28212
rect 15016 28024 15068 28076
rect 14372 27956 14424 28008
rect 15292 28067 15344 28076
rect 15292 28033 15306 28067
rect 15306 28033 15340 28067
rect 15340 28033 15344 28067
rect 15292 28024 15344 28033
rect 16304 28024 16356 28076
rect 19340 28024 19392 28076
rect 20720 28067 20772 28076
rect 20720 28033 20729 28067
rect 20729 28033 20763 28067
rect 20763 28033 20772 28067
rect 20720 28024 20772 28033
rect 16856 27956 16908 28008
rect 20444 27999 20496 28008
rect 20444 27965 20453 27999
rect 20453 27965 20487 27999
rect 20487 27965 20496 27999
rect 20444 27956 20496 27965
rect 12900 27888 12952 27940
rect 15108 27888 15160 27940
rect 18328 27888 18380 27940
rect 4620 27820 4672 27872
rect 9220 27820 9272 27872
rect 9772 27863 9824 27872
rect 9772 27829 9781 27863
rect 9781 27829 9815 27863
rect 9815 27829 9824 27863
rect 9772 27820 9824 27829
rect 11980 27820 12032 27872
rect 15384 27820 15436 27872
rect 18420 27820 18472 27872
rect 19984 27820 20036 27872
rect 22008 27863 22060 27872
rect 22008 27829 22017 27863
rect 22017 27829 22051 27863
rect 22051 27829 22060 27863
rect 22008 27820 22060 27829
rect 23020 27820 23072 27872
rect 23572 28024 23624 28076
rect 29920 28024 29972 28076
rect 32496 28024 32548 28076
rect 33416 28092 33468 28144
rect 32956 28067 33008 28076
rect 24308 27820 24360 27872
rect 30564 27999 30616 28008
rect 30564 27965 30573 27999
rect 30573 27965 30607 27999
rect 30607 27965 30616 27999
rect 30564 27956 30616 27965
rect 32956 28033 32965 28067
rect 32965 28033 32999 28067
rect 32999 28033 33008 28067
rect 32956 28024 33008 28033
rect 33784 28067 33836 28076
rect 33784 28033 33793 28067
rect 33793 28033 33827 28067
rect 33827 28033 33836 28067
rect 33784 28024 33836 28033
rect 34060 28024 34112 28076
rect 34520 28067 34572 28076
rect 34520 28033 34529 28067
rect 34529 28033 34563 28067
rect 34563 28033 34572 28067
rect 34520 28024 34572 28033
rect 37280 28024 37332 28076
rect 32588 27888 32640 27940
rect 38660 28024 38712 28076
rect 58164 27931 58216 27940
rect 58164 27897 58173 27931
rect 58173 27897 58207 27931
rect 58207 27897 58216 27931
rect 58164 27888 58216 27897
rect 32404 27863 32456 27872
rect 32404 27829 32413 27863
rect 32413 27829 32447 27863
rect 32447 27829 32456 27863
rect 32404 27820 32456 27829
rect 33508 27820 33560 27872
rect 34796 27820 34848 27872
rect 40224 27863 40276 27872
rect 40224 27829 40233 27863
rect 40233 27829 40267 27863
rect 40267 27829 40276 27863
rect 40224 27820 40276 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2596 27659 2648 27668
rect 2596 27625 2605 27659
rect 2605 27625 2639 27659
rect 2639 27625 2648 27659
rect 2596 27616 2648 27625
rect 6920 27659 6972 27668
rect 6920 27625 6929 27659
rect 6929 27625 6963 27659
rect 6963 27625 6972 27659
rect 6920 27616 6972 27625
rect 4896 27548 4948 27600
rect 10968 27616 11020 27668
rect 13084 27659 13136 27668
rect 4620 27480 4672 27532
rect 3332 27412 3384 27464
rect 3884 27412 3936 27464
rect 4712 27455 4764 27464
rect 4712 27421 4721 27455
rect 4721 27421 4755 27455
rect 4755 27421 4764 27455
rect 4712 27412 4764 27421
rect 4988 27455 5040 27464
rect 3148 27344 3200 27396
rect 3976 27387 4028 27396
rect 3976 27353 3985 27387
rect 3985 27353 4019 27387
rect 4019 27353 4028 27387
rect 3976 27344 4028 27353
rect 2964 27276 3016 27328
rect 3608 27276 3660 27328
rect 4988 27421 4997 27455
rect 4997 27421 5031 27455
rect 5031 27421 5040 27455
rect 4988 27412 5040 27421
rect 11704 27548 11756 27600
rect 13084 27625 13093 27659
rect 13093 27625 13127 27659
rect 13127 27625 13136 27659
rect 13084 27616 13136 27625
rect 16120 27616 16172 27668
rect 19340 27591 19392 27600
rect 19340 27557 19349 27591
rect 19349 27557 19383 27591
rect 19383 27557 19392 27591
rect 23112 27616 23164 27668
rect 25228 27616 25280 27668
rect 32404 27616 32456 27668
rect 37280 27659 37332 27668
rect 37280 27625 37289 27659
rect 37289 27625 37323 27659
rect 37323 27625 37332 27659
rect 37280 27616 37332 27625
rect 19340 27548 19392 27557
rect 28448 27548 28500 27600
rect 5448 27412 5500 27464
rect 5908 27412 5960 27464
rect 7104 27412 7156 27464
rect 7472 27480 7524 27532
rect 8944 27480 8996 27532
rect 15292 27480 15344 27532
rect 21272 27480 21324 27532
rect 7380 27455 7432 27464
rect 7380 27421 7389 27455
rect 7389 27421 7423 27455
rect 7423 27421 7432 27455
rect 7380 27412 7432 27421
rect 7564 27455 7616 27464
rect 7564 27421 7573 27455
rect 7573 27421 7607 27455
rect 7607 27421 7616 27455
rect 9772 27455 9824 27464
rect 7564 27412 7616 27421
rect 4896 27276 4948 27328
rect 5080 27276 5132 27328
rect 9772 27421 9781 27455
rect 9781 27421 9815 27455
rect 9815 27421 9824 27455
rect 9772 27412 9824 27421
rect 9956 27455 10008 27464
rect 9956 27421 9965 27455
rect 9965 27421 9999 27455
rect 9999 27421 10008 27455
rect 9956 27412 10008 27421
rect 13452 27412 13504 27464
rect 20812 27412 20864 27464
rect 22008 27480 22060 27532
rect 26792 27523 26844 27532
rect 26792 27489 26801 27523
rect 26801 27489 26835 27523
rect 26835 27489 26844 27523
rect 26792 27480 26844 27489
rect 11980 27387 12032 27396
rect 11980 27353 12014 27387
rect 12014 27353 12032 27387
rect 11980 27344 12032 27353
rect 12164 27344 12216 27396
rect 14832 27344 14884 27396
rect 17040 27387 17092 27396
rect 8116 27319 8168 27328
rect 8116 27285 8125 27319
rect 8125 27285 8159 27319
rect 8159 27285 8168 27319
rect 8116 27276 8168 27285
rect 10416 27319 10468 27328
rect 10416 27285 10425 27319
rect 10425 27285 10459 27319
rect 10459 27285 10468 27319
rect 10416 27276 10468 27285
rect 15016 27276 15068 27328
rect 17040 27353 17049 27387
rect 17049 27353 17083 27387
rect 17083 27353 17092 27387
rect 17040 27344 17092 27353
rect 21640 27412 21692 27464
rect 31760 27548 31812 27600
rect 31576 27480 31628 27532
rect 32496 27480 32548 27532
rect 32772 27480 32824 27532
rect 31392 27455 31444 27464
rect 21548 27276 21600 27328
rect 21824 27319 21876 27328
rect 21824 27285 21833 27319
rect 21833 27285 21867 27319
rect 21867 27285 21876 27319
rect 21824 27276 21876 27285
rect 22560 27344 22612 27396
rect 23204 27344 23256 27396
rect 23756 27344 23808 27396
rect 24860 27344 24912 27396
rect 25964 27344 26016 27396
rect 29000 27344 29052 27396
rect 30380 27344 30432 27396
rect 31392 27421 31401 27455
rect 31401 27421 31435 27455
rect 31435 27421 31444 27455
rect 31392 27412 31444 27421
rect 33232 27480 33284 27532
rect 33140 27412 33192 27464
rect 33416 27412 33468 27464
rect 33968 27455 34020 27464
rect 33968 27421 33977 27455
rect 33977 27421 34011 27455
rect 34011 27421 34020 27455
rect 33968 27412 34020 27421
rect 34520 27412 34572 27464
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 34796 27412 34848 27464
rect 35072 27455 35124 27464
rect 35072 27421 35081 27455
rect 35081 27421 35115 27455
rect 35115 27421 35124 27455
rect 35072 27412 35124 27421
rect 35440 27412 35492 27464
rect 38568 27412 38620 27464
rect 40224 27412 40276 27464
rect 33784 27387 33836 27396
rect 23388 27276 23440 27328
rect 23848 27319 23900 27328
rect 23848 27285 23857 27319
rect 23857 27285 23891 27319
rect 23891 27285 23900 27319
rect 23848 27276 23900 27285
rect 24124 27276 24176 27328
rect 26332 27319 26384 27328
rect 26332 27285 26341 27319
rect 26341 27285 26375 27319
rect 26375 27285 26384 27319
rect 26332 27276 26384 27285
rect 29368 27276 29420 27328
rect 29552 27319 29604 27328
rect 29552 27285 29561 27319
rect 29561 27285 29595 27319
rect 29595 27285 29604 27319
rect 29552 27276 29604 27285
rect 33784 27353 33793 27387
rect 33793 27353 33827 27387
rect 33827 27353 33836 27387
rect 33784 27344 33836 27353
rect 33232 27276 33284 27328
rect 33416 27276 33468 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 3516 27072 3568 27124
rect 2688 26936 2740 26988
rect 3424 26979 3476 26988
rect 3424 26945 3433 26979
rect 3433 26945 3467 26979
rect 3467 26945 3476 26979
rect 3424 26936 3476 26945
rect 3608 26982 3660 26988
rect 3608 26948 3617 26982
rect 3617 26948 3651 26982
rect 3651 26948 3660 26982
rect 3608 26936 3660 26948
rect 4896 27072 4948 27124
rect 4988 27072 5040 27124
rect 4804 26979 4856 26988
rect 4804 26945 4813 26979
rect 4813 26945 4847 26979
rect 4847 26945 4856 26979
rect 4804 26936 4856 26945
rect 8944 27072 8996 27124
rect 16120 27072 16172 27124
rect 17132 27072 17184 27124
rect 24676 27072 24728 27124
rect 24860 27115 24912 27124
rect 24860 27081 24869 27115
rect 24869 27081 24903 27115
rect 24903 27081 24912 27115
rect 24860 27072 24912 27081
rect 25964 27115 26016 27124
rect 25964 27081 25973 27115
rect 25973 27081 26007 27115
rect 26007 27081 26016 27115
rect 25964 27072 26016 27081
rect 30564 27072 30616 27124
rect 31484 27072 31536 27124
rect 33140 27072 33192 27124
rect 33968 27072 34020 27124
rect 35072 27115 35124 27124
rect 35072 27081 35081 27115
rect 35081 27081 35115 27115
rect 35115 27081 35124 27115
rect 35072 27072 35124 27081
rect 3700 26868 3752 26920
rect 7748 27004 7800 27056
rect 12348 27004 12400 27056
rect 14832 27047 14884 27056
rect 14832 27013 14841 27047
rect 14841 27013 14875 27047
rect 14875 27013 14884 27047
rect 14832 27004 14884 27013
rect 21824 27004 21876 27056
rect 24124 27004 24176 27056
rect 6736 26979 6788 26988
rect 6736 26945 6745 26979
rect 6745 26945 6779 26979
rect 6779 26945 6788 26979
rect 6736 26936 6788 26945
rect 6828 26979 6880 26988
rect 6828 26945 6838 26979
rect 6838 26945 6872 26979
rect 6872 26945 6880 26979
rect 6828 26936 6880 26945
rect 5448 26868 5500 26920
rect 9128 26936 9180 26988
rect 9956 26936 10008 26988
rect 13728 26936 13780 26988
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16120 26936 16172 26945
rect 10876 26868 10928 26920
rect 18972 26979 19024 26988
rect 18972 26945 18981 26979
rect 18981 26945 19015 26979
rect 19015 26945 19024 26979
rect 18972 26936 19024 26945
rect 19156 26979 19208 26988
rect 19156 26945 19165 26979
rect 19165 26945 19199 26979
rect 19199 26945 19208 26979
rect 19156 26936 19208 26945
rect 20904 26936 20956 26988
rect 24216 26979 24268 26988
rect 24216 26945 24225 26979
rect 24225 26945 24259 26979
rect 24259 26945 24268 26979
rect 24216 26936 24268 26945
rect 24400 26979 24452 26988
rect 24400 26945 24409 26979
rect 24409 26945 24443 26979
rect 24443 26945 24452 26979
rect 24400 26936 24452 26945
rect 31576 27004 31628 27056
rect 16580 26868 16632 26920
rect 18696 26868 18748 26920
rect 21640 26868 21692 26920
rect 24768 26936 24820 26988
rect 25504 26979 25556 26988
rect 25504 26945 25513 26979
rect 25513 26945 25547 26979
rect 25547 26945 25556 26979
rect 25504 26936 25556 26945
rect 25044 26868 25096 26920
rect 25780 26936 25832 26988
rect 5264 26800 5316 26852
rect 21456 26800 21508 26852
rect 2688 26775 2740 26784
rect 2688 26741 2697 26775
rect 2697 26741 2731 26775
rect 2731 26741 2740 26775
rect 2688 26732 2740 26741
rect 3148 26775 3200 26784
rect 3148 26741 3157 26775
rect 3157 26741 3191 26775
rect 3191 26741 3200 26775
rect 3148 26732 3200 26741
rect 5448 26775 5500 26784
rect 5448 26741 5457 26775
rect 5457 26741 5491 26775
rect 5491 26741 5500 26775
rect 5448 26732 5500 26741
rect 7380 26775 7432 26784
rect 7380 26741 7389 26775
rect 7389 26741 7423 26775
rect 7423 26741 7432 26775
rect 7380 26732 7432 26741
rect 16396 26732 16448 26784
rect 19708 26732 19760 26784
rect 22928 26732 22980 26784
rect 23664 26732 23716 26784
rect 29000 26936 29052 26988
rect 29828 26936 29880 26988
rect 33416 26979 33468 26988
rect 33416 26945 33450 26979
rect 33450 26945 33468 26979
rect 33416 26936 33468 26945
rect 28724 26732 28776 26784
rect 31392 26868 31444 26920
rect 58164 26775 58216 26784
rect 58164 26741 58173 26775
rect 58173 26741 58207 26775
rect 58207 26741 58216 26775
rect 58164 26732 58216 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3884 26528 3936 26580
rect 2596 26324 2648 26376
rect 3700 26392 3752 26444
rect 3884 26324 3936 26376
rect 4068 26367 4120 26376
rect 4068 26333 4077 26367
rect 4077 26333 4111 26367
rect 4111 26333 4120 26367
rect 4068 26324 4120 26333
rect 4896 26324 4948 26376
rect 7564 26528 7616 26580
rect 8116 26528 8168 26580
rect 11060 26528 11112 26580
rect 12348 26528 12400 26580
rect 6552 26392 6604 26444
rect 6000 26324 6052 26376
rect 6368 26324 6420 26376
rect 6828 26324 6880 26376
rect 7472 26460 7524 26512
rect 21824 26528 21876 26580
rect 24216 26528 24268 26580
rect 25504 26528 25556 26580
rect 31576 26528 31628 26580
rect 32588 26571 32640 26580
rect 32588 26537 32597 26571
rect 32597 26537 32631 26571
rect 32631 26537 32640 26571
rect 32588 26528 32640 26537
rect 15936 26460 15988 26512
rect 20352 26503 20404 26512
rect 14372 26435 14424 26444
rect 14372 26401 14381 26435
rect 14381 26401 14415 26435
rect 14415 26401 14424 26435
rect 14372 26392 14424 26401
rect 16396 26435 16448 26444
rect 16396 26401 16405 26435
rect 16405 26401 16439 26435
rect 16439 26401 16448 26435
rect 16396 26392 16448 26401
rect 20352 26469 20361 26503
rect 20361 26469 20395 26503
rect 20395 26469 20404 26503
rect 20352 26460 20404 26469
rect 23204 26460 23256 26512
rect 19064 26392 19116 26444
rect 3700 26256 3752 26308
rect 3516 26188 3568 26240
rect 10600 26324 10652 26376
rect 11704 26367 11756 26376
rect 11704 26333 11713 26367
rect 11713 26333 11747 26367
rect 11747 26333 11756 26367
rect 11704 26324 11756 26333
rect 13452 26324 13504 26376
rect 16120 26367 16172 26376
rect 16120 26333 16129 26367
rect 16129 26333 16163 26367
rect 16163 26333 16172 26367
rect 16120 26324 16172 26333
rect 4620 26256 4672 26308
rect 4988 26256 5040 26308
rect 6552 26256 6604 26308
rect 6736 26299 6788 26308
rect 6736 26265 6745 26299
rect 6745 26265 6779 26299
rect 6779 26265 6788 26299
rect 6736 26256 6788 26265
rect 7564 26256 7616 26308
rect 10416 26256 10468 26308
rect 15108 26256 15160 26308
rect 18696 26324 18748 26376
rect 21272 26392 21324 26444
rect 22008 26392 22060 26444
rect 25780 26392 25832 26444
rect 38568 26392 38620 26444
rect 16948 26299 17000 26308
rect 16948 26265 16957 26299
rect 16957 26265 16991 26299
rect 16991 26265 17000 26299
rect 16948 26256 17000 26265
rect 19708 26367 19760 26376
rect 19708 26333 19717 26367
rect 19717 26333 19751 26367
rect 19751 26333 19760 26367
rect 19708 26324 19760 26333
rect 20812 26324 20864 26376
rect 32588 26324 32640 26376
rect 38936 26324 38988 26376
rect 20352 26256 20404 26308
rect 21640 26299 21692 26308
rect 21640 26265 21649 26299
rect 21649 26265 21683 26299
rect 21683 26265 21692 26299
rect 21640 26256 21692 26265
rect 23664 26256 23716 26308
rect 24216 26256 24268 26308
rect 24400 26299 24452 26308
rect 24400 26265 24409 26299
rect 24409 26265 24443 26299
rect 24443 26265 24452 26299
rect 24400 26256 24452 26265
rect 7472 26188 7524 26240
rect 18420 26188 18472 26240
rect 18604 26188 18656 26240
rect 19248 26231 19300 26240
rect 19248 26197 19257 26231
rect 19257 26197 19291 26231
rect 19291 26197 19300 26231
rect 19248 26188 19300 26197
rect 23480 26188 23532 26240
rect 23848 26188 23900 26240
rect 26148 26256 26200 26308
rect 29368 26256 29420 26308
rect 37280 26256 37332 26308
rect 39028 26256 39080 26308
rect 29644 26231 29696 26240
rect 29644 26197 29653 26231
rect 29653 26197 29687 26231
rect 29687 26197 29696 26231
rect 29644 26188 29696 26197
rect 36636 26188 36688 26240
rect 38016 26188 38068 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 3976 26027 4028 26036
rect 3976 25993 3985 26027
rect 3985 25993 4019 26027
rect 4019 25993 4028 26027
rect 3976 25984 4028 25993
rect 4068 25984 4120 26036
rect 6368 26027 6420 26036
rect 6368 25993 6377 26027
rect 6377 25993 6411 26027
rect 6411 25993 6420 26027
rect 6368 25984 6420 25993
rect 14372 25984 14424 26036
rect 19156 25984 19208 26036
rect 20720 25984 20772 26036
rect 21088 25984 21140 26036
rect 21272 25984 21324 26036
rect 3148 25916 3200 25968
rect 4896 25916 4948 25968
rect 6736 25916 6788 25968
rect 13912 25916 13964 25968
rect 14648 25959 14700 25968
rect 14648 25925 14657 25959
rect 14657 25925 14691 25959
rect 14691 25925 14700 25959
rect 14648 25916 14700 25925
rect 15016 25916 15068 25968
rect 19248 25959 19300 25968
rect 19248 25925 19266 25959
rect 19266 25925 19300 25959
rect 19248 25916 19300 25925
rect 20812 25916 20864 25968
rect 2320 25848 2372 25900
rect 9680 25891 9732 25900
rect 9680 25857 9689 25891
rect 9689 25857 9723 25891
rect 9723 25857 9732 25891
rect 9680 25848 9732 25857
rect 11704 25848 11756 25900
rect 6828 25644 6880 25696
rect 9772 25780 9824 25832
rect 12992 25780 13044 25832
rect 14280 25848 14332 25900
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 17224 25848 17276 25900
rect 22560 25984 22612 26036
rect 23388 25984 23440 26036
rect 30380 25984 30432 26036
rect 37280 26027 37332 26036
rect 37280 25993 37289 26027
rect 37289 25993 37323 26027
rect 37323 25993 37332 26027
rect 37280 25984 37332 25993
rect 23572 25959 23624 25968
rect 23572 25925 23581 25959
rect 23581 25925 23615 25959
rect 23615 25925 23624 25959
rect 23572 25916 23624 25925
rect 10784 25644 10836 25696
rect 13084 25644 13136 25696
rect 15568 25687 15620 25696
rect 15568 25653 15577 25687
rect 15577 25653 15611 25687
rect 15611 25653 15620 25687
rect 15568 25644 15620 25653
rect 15660 25644 15712 25696
rect 19248 25644 19300 25696
rect 21640 25780 21692 25832
rect 22192 25891 22244 25900
rect 22192 25857 22201 25891
rect 22201 25857 22235 25891
rect 22235 25857 22244 25891
rect 22192 25848 22244 25857
rect 23112 25848 23164 25900
rect 24216 25916 24268 25968
rect 26332 25916 26384 25968
rect 27436 25916 27488 25968
rect 23204 25780 23256 25832
rect 23388 25712 23440 25764
rect 23848 25891 23900 25900
rect 23848 25857 23857 25891
rect 23857 25857 23891 25891
rect 23891 25857 23900 25891
rect 23848 25848 23900 25857
rect 24400 25848 24452 25900
rect 26056 25848 26108 25900
rect 27620 25848 27672 25900
rect 31576 25916 31628 25968
rect 38752 25916 38804 25968
rect 29644 25891 29696 25900
rect 29644 25857 29653 25891
rect 29653 25857 29687 25891
rect 29687 25857 29696 25891
rect 29644 25848 29696 25857
rect 29828 25891 29880 25900
rect 29828 25857 29837 25891
rect 29837 25857 29871 25891
rect 29871 25857 29880 25891
rect 29828 25848 29880 25857
rect 24492 25780 24544 25832
rect 28816 25823 28868 25832
rect 28816 25789 28825 25823
rect 28825 25789 28859 25823
rect 28859 25789 28868 25823
rect 28816 25780 28868 25789
rect 30196 25848 30248 25900
rect 27804 25712 27856 25764
rect 29920 25712 29972 25764
rect 30380 25712 30432 25764
rect 37188 25848 37240 25900
rect 37556 25712 37608 25764
rect 37832 25848 37884 25900
rect 37924 25891 37976 25900
rect 37924 25857 37933 25891
rect 37933 25857 37967 25891
rect 37967 25857 37976 25891
rect 37924 25848 37976 25857
rect 38568 25848 38620 25900
rect 40224 25848 40276 25900
rect 22192 25644 22244 25696
rect 23296 25644 23348 25696
rect 27896 25644 27948 25696
rect 30196 25644 30248 25696
rect 37464 25644 37516 25696
rect 38936 25644 38988 25696
rect 39856 25644 39908 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 9036 25483 9088 25492
rect 9036 25449 9045 25483
rect 9045 25449 9079 25483
rect 9079 25449 9088 25483
rect 9036 25440 9088 25449
rect 3792 25372 3844 25424
rect 10140 25372 10192 25424
rect 17224 25440 17276 25492
rect 18420 25440 18472 25492
rect 16948 25372 17000 25424
rect 11060 25304 11112 25356
rect 12164 25347 12216 25356
rect 12164 25313 12173 25347
rect 12173 25313 12207 25347
rect 12207 25313 12216 25347
rect 12164 25304 12216 25313
rect 22376 25440 22428 25492
rect 23388 25440 23440 25492
rect 26976 25440 27028 25492
rect 29828 25440 29880 25492
rect 37832 25440 37884 25492
rect 38568 25483 38620 25492
rect 38568 25449 38577 25483
rect 38577 25449 38611 25483
rect 38611 25449 38620 25483
rect 38568 25440 38620 25449
rect 19248 25347 19300 25356
rect 19248 25313 19257 25347
rect 19257 25313 19291 25347
rect 19291 25313 19300 25347
rect 19248 25304 19300 25313
rect 22652 25304 22704 25356
rect 9036 25236 9088 25288
rect 10048 25279 10100 25288
rect 10048 25245 10062 25279
rect 10062 25245 10096 25279
rect 10096 25245 10100 25279
rect 10048 25236 10100 25245
rect 10968 25236 11020 25288
rect 13820 25236 13872 25288
rect 23112 25279 23164 25288
rect 5540 25211 5592 25220
rect 5540 25177 5549 25211
rect 5549 25177 5583 25211
rect 5583 25177 5592 25211
rect 5540 25168 5592 25177
rect 9588 25143 9640 25152
rect 9588 25109 9597 25143
rect 9597 25109 9631 25143
rect 9631 25109 9640 25143
rect 9588 25100 9640 25109
rect 12624 25168 12676 25220
rect 14740 25168 14792 25220
rect 11060 25100 11112 25152
rect 12164 25100 12216 25152
rect 12716 25100 12768 25152
rect 13912 25100 13964 25152
rect 14280 25143 14332 25152
rect 14280 25109 14289 25143
rect 14289 25109 14323 25143
rect 14323 25109 14332 25143
rect 14280 25100 14332 25109
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 18328 25143 18380 25152
rect 18328 25109 18337 25143
rect 18337 25109 18371 25143
rect 18371 25109 18380 25143
rect 18328 25100 18380 25109
rect 19432 25100 19484 25152
rect 20628 25143 20680 25152
rect 20628 25109 20637 25143
rect 20637 25109 20671 25143
rect 20671 25109 20680 25143
rect 20628 25100 20680 25109
rect 23112 25245 23116 25279
rect 23116 25245 23150 25279
rect 23150 25245 23164 25279
rect 23112 25236 23164 25245
rect 23204 25279 23256 25288
rect 23204 25245 23213 25279
rect 23213 25245 23247 25279
rect 23247 25245 23256 25279
rect 23480 25279 23532 25288
rect 23204 25236 23256 25245
rect 23480 25245 23488 25279
rect 23488 25245 23522 25279
rect 23522 25245 23532 25279
rect 23480 25236 23532 25245
rect 28816 25304 28868 25356
rect 29920 25304 29972 25356
rect 24768 25279 24820 25288
rect 24768 25245 24777 25279
rect 24777 25245 24811 25279
rect 24811 25245 24820 25279
rect 24768 25236 24820 25245
rect 24952 25279 25004 25288
rect 24952 25245 24961 25279
rect 24961 25245 24995 25279
rect 24995 25245 25004 25279
rect 24952 25236 25004 25245
rect 25044 25279 25096 25288
rect 25044 25245 25053 25279
rect 25053 25245 25087 25279
rect 25087 25245 25096 25279
rect 25044 25236 25096 25245
rect 23204 25100 23256 25152
rect 24032 25168 24084 25220
rect 24584 25168 24636 25220
rect 28908 25236 28960 25288
rect 29736 25236 29788 25288
rect 30012 25279 30064 25288
rect 30012 25245 30021 25279
rect 30021 25245 30055 25279
rect 30055 25245 30064 25279
rect 30012 25236 30064 25245
rect 38016 25304 38068 25356
rect 27804 25168 27856 25220
rect 29552 25168 29604 25220
rect 23572 25100 23624 25152
rect 25780 25100 25832 25152
rect 28540 25100 28592 25152
rect 30380 25236 30432 25288
rect 31576 25236 31628 25288
rect 36728 25236 36780 25288
rect 37464 25279 37516 25288
rect 37464 25245 37473 25279
rect 37473 25245 37507 25279
rect 37507 25245 37516 25279
rect 37464 25236 37516 25245
rect 37740 25236 37792 25288
rect 37924 25279 37976 25288
rect 37924 25245 37933 25279
rect 37933 25245 37967 25279
rect 37967 25245 37976 25279
rect 37924 25236 37976 25245
rect 58164 25279 58216 25288
rect 36636 25211 36688 25220
rect 36636 25177 36645 25211
rect 36645 25177 36679 25211
rect 36679 25177 36688 25211
rect 36636 25168 36688 25177
rect 30564 25100 30616 25152
rect 37556 25100 37608 25152
rect 58164 25245 58173 25279
rect 58173 25245 58207 25279
rect 58207 25245 58216 25279
rect 58164 25236 58216 25245
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 2596 24939 2648 24948
rect 2596 24905 2605 24939
rect 2605 24905 2639 24939
rect 2639 24905 2648 24939
rect 2596 24896 2648 24905
rect 12624 24939 12676 24948
rect 12624 24905 12633 24939
rect 12633 24905 12667 24939
rect 12667 24905 12676 24939
rect 12624 24896 12676 24905
rect 14740 24939 14792 24948
rect 14740 24905 14749 24939
rect 14749 24905 14783 24939
rect 14783 24905 14792 24939
rect 14740 24896 14792 24905
rect 15568 24896 15620 24948
rect 16028 24896 16080 24948
rect 2320 24828 2372 24880
rect 3700 24803 3752 24812
rect 9588 24828 9640 24880
rect 10140 24828 10192 24880
rect 3700 24769 3718 24803
rect 3718 24769 3752 24803
rect 3700 24760 3752 24769
rect 5540 24760 5592 24812
rect 6092 24760 6144 24812
rect 11060 24828 11112 24880
rect 12716 24828 12768 24880
rect 6828 24692 6880 24744
rect 10784 24803 10836 24812
rect 10784 24769 10798 24803
rect 10798 24769 10832 24803
rect 10832 24769 10836 24803
rect 10784 24760 10836 24769
rect 10968 24803 11020 24812
rect 10968 24769 10977 24803
rect 10977 24769 11011 24803
rect 11011 24769 11020 24803
rect 12900 24803 12952 24812
rect 10968 24760 11020 24769
rect 12900 24769 12909 24803
rect 12909 24769 12943 24803
rect 12943 24769 12952 24803
rect 12900 24760 12952 24769
rect 13084 24803 13136 24812
rect 13084 24769 13093 24803
rect 13093 24769 13127 24803
rect 13127 24769 13136 24803
rect 13084 24760 13136 24769
rect 13268 24803 13320 24812
rect 13268 24769 13277 24803
rect 13277 24769 13311 24803
rect 13311 24769 13320 24803
rect 13268 24760 13320 24769
rect 14188 24760 14240 24812
rect 16120 24828 16172 24880
rect 19432 24896 19484 24948
rect 24768 24896 24820 24948
rect 24952 24896 25004 24948
rect 27620 24939 27672 24948
rect 27620 24905 27629 24939
rect 27629 24905 27663 24939
rect 27663 24905 27672 24939
rect 27620 24896 27672 24905
rect 20628 24828 20680 24880
rect 22928 24828 22980 24880
rect 23204 24828 23256 24880
rect 25780 24828 25832 24880
rect 30012 24896 30064 24948
rect 38844 24828 38896 24880
rect 15200 24803 15252 24812
rect 15200 24769 15209 24803
rect 15209 24769 15243 24803
rect 15243 24769 15252 24803
rect 15200 24760 15252 24769
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 18880 24803 18932 24812
rect 12900 24624 12952 24676
rect 18880 24769 18889 24803
rect 18889 24769 18923 24803
rect 18923 24769 18932 24803
rect 18880 24760 18932 24769
rect 6460 24556 6512 24608
rect 8024 24556 8076 24608
rect 9864 24599 9916 24608
rect 9864 24565 9873 24599
rect 9873 24565 9907 24599
rect 9907 24565 9916 24599
rect 9864 24556 9916 24565
rect 10324 24599 10376 24608
rect 10324 24565 10333 24599
rect 10333 24565 10367 24599
rect 10367 24565 10376 24599
rect 10324 24556 10376 24565
rect 11060 24556 11112 24608
rect 14188 24599 14240 24608
rect 14188 24565 14197 24599
rect 14197 24565 14231 24599
rect 14231 24565 14240 24599
rect 14188 24556 14240 24565
rect 16120 24599 16172 24608
rect 16120 24565 16129 24599
rect 16129 24565 16163 24599
rect 16163 24565 16172 24599
rect 16120 24556 16172 24565
rect 17408 24556 17460 24608
rect 19340 24760 19392 24812
rect 20260 24760 20312 24812
rect 22652 24760 22704 24812
rect 23112 24760 23164 24812
rect 23572 24803 23624 24812
rect 23572 24769 23617 24803
rect 23617 24769 23624 24803
rect 23572 24760 23624 24769
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 24584 24803 24636 24812
rect 23756 24760 23808 24769
rect 24584 24769 24593 24803
rect 24593 24769 24627 24803
rect 24627 24769 24636 24803
rect 24584 24760 24636 24769
rect 26056 24760 26108 24812
rect 27804 24760 27856 24812
rect 19156 24624 19208 24676
rect 23112 24599 23164 24608
rect 23112 24565 23121 24599
rect 23121 24565 23155 24599
rect 23155 24565 23164 24599
rect 23112 24556 23164 24565
rect 27252 24556 27304 24608
rect 27804 24624 27856 24676
rect 28080 24803 28132 24812
rect 28080 24769 28094 24803
rect 28094 24769 28128 24803
rect 28128 24769 28132 24803
rect 28264 24803 28316 24812
rect 28080 24760 28132 24769
rect 28264 24769 28273 24803
rect 28273 24769 28307 24803
rect 28307 24769 28316 24803
rect 28264 24760 28316 24769
rect 28908 24760 28960 24812
rect 30564 24760 30616 24812
rect 30840 24760 30892 24812
rect 31576 24803 31628 24812
rect 31576 24769 31585 24803
rect 31585 24769 31619 24803
rect 31619 24769 31628 24803
rect 31576 24760 31628 24769
rect 33600 24760 33652 24812
rect 37372 24760 37424 24812
rect 37924 24803 37976 24812
rect 37924 24769 37933 24803
rect 37933 24769 37967 24803
rect 37967 24769 37976 24803
rect 37924 24760 37976 24769
rect 39028 24803 39080 24812
rect 37464 24692 37516 24744
rect 33048 24624 33100 24676
rect 28632 24556 28684 24608
rect 29828 24556 29880 24608
rect 33876 24599 33928 24608
rect 33876 24565 33885 24599
rect 33885 24565 33919 24599
rect 33919 24565 33928 24599
rect 33876 24556 33928 24565
rect 37556 24624 37608 24676
rect 39028 24769 39037 24803
rect 39037 24769 39071 24803
rect 39071 24769 39080 24803
rect 39028 24760 39080 24769
rect 39856 24828 39908 24880
rect 38752 24624 38804 24676
rect 40132 24556 40184 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 5816 24395 5868 24404
rect 5816 24361 5825 24395
rect 5825 24361 5859 24395
rect 5859 24361 5868 24395
rect 5816 24352 5868 24361
rect 12532 24352 12584 24404
rect 8024 24284 8076 24336
rect 15016 24352 15068 24404
rect 15200 24395 15252 24404
rect 15200 24361 15209 24395
rect 15209 24361 15243 24395
rect 15243 24361 15252 24395
rect 15200 24352 15252 24361
rect 15384 24352 15436 24404
rect 16304 24352 16356 24404
rect 17408 24352 17460 24404
rect 19984 24352 20036 24404
rect 21456 24395 21508 24404
rect 21456 24361 21465 24395
rect 21465 24361 21499 24395
rect 21499 24361 21508 24395
rect 21456 24352 21508 24361
rect 21916 24352 21968 24404
rect 5540 24216 5592 24268
rect 6828 24216 6880 24268
rect 10048 24259 10100 24268
rect 10048 24225 10057 24259
rect 10057 24225 10091 24259
rect 10091 24225 10100 24259
rect 10048 24216 10100 24225
rect 6460 24191 6512 24200
rect 6460 24157 6469 24191
rect 6469 24157 6503 24191
rect 6503 24157 6512 24191
rect 6460 24148 6512 24157
rect 10324 24148 10376 24200
rect 11060 24148 11112 24200
rect 12348 24148 12400 24200
rect 12624 24148 12676 24200
rect 13268 24284 13320 24336
rect 19340 24284 19392 24336
rect 24584 24352 24636 24404
rect 28080 24395 28132 24404
rect 28080 24361 28089 24395
rect 28089 24361 28123 24395
rect 28123 24361 28132 24395
rect 28080 24352 28132 24361
rect 28632 24352 28684 24404
rect 29736 24352 29788 24404
rect 30104 24352 30156 24404
rect 30840 24352 30892 24404
rect 31760 24352 31812 24404
rect 33600 24395 33652 24404
rect 33600 24361 33609 24395
rect 33609 24361 33643 24395
rect 33643 24361 33652 24395
rect 33600 24352 33652 24361
rect 38660 24352 38712 24404
rect 22744 24284 22796 24336
rect 18328 24216 18380 24268
rect 18972 24216 19024 24268
rect 20260 24216 20312 24268
rect 20628 24216 20680 24268
rect 6092 24080 6144 24132
rect 6828 24080 6880 24132
rect 9864 24123 9916 24132
rect 6276 24055 6328 24064
rect 6276 24021 6285 24055
rect 6285 24021 6319 24055
rect 6319 24021 6328 24055
rect 6276 24012 6328 24021
rect 9588 24012 9640 24064
rect 9864 24089 9873 24123
rect 9873 24089 9907 24123
rect 9907 24089 9916 24123
rect 9864 24080 9916 24089
rect 11152 24123 11204 24132
rect 9772 24012 9824 24064
rect 11152 24089 11161 24123
rect 11161 24089 11195 24123
rect 11195 24089 11204 24123
rect 11152 24080 11204 24089
rect 11336 24123 11388 24132
rect 11336 24089 11345 24123
rect 11345 24089 11379 24123
rect 11379 24089 11388 24123
rect 11336 24080 11388 24089
rect 12992 24080 13044 24132
rect 11796 24055 11848 24064
rect 11796 24021 11805 24055
rect 11805 24021 11839 24055
rect 11839 24021 11848 24055
rect 11796 24012 11848 24021
rect 12164 24012 12216 24064
rect 12532 24012 12584 24064
rect 14372 24148 14424 24200
rect 15476 24148 15528 24200
rect 16212 24148 16264 24200
rect 17408 24191 17460 24200
rect 14096 24080 14148 24132
rect 15292 24080 15344 24132
rect 15660 24080 15712 24132
rect 13912 24012 13964 24064
rect 14372 24012 14424 24064
rect 14740 24055 14792 24064
rect 14740 24021 14749 24055
rect 14749 24021 14783 24055
rect 14783 24021 14792 24055
rect 14740 24012 14792 24021
rect 15016 24012 15068 24064
rect 17408 24157 17417 24191
rect 17417 24157 17451 24191
rect 17451 24157 17460 24191
rect 17408 24148 17460 24157
rect 17592 24191 17644 24200
rect 17592 24157 17601 24191
rect 17601 24157 17635 24191
rect 17635 24157 17644 24191
rect 17592 24148 17644 24157
rect 19984 24148 20036 24200
rect 22652 24148 22704 24200
rect 27252 24259 27304 24268
rect 27252 24225 27261 24259
rect 27261 24225 27295 24259
rect 27295 24225 27304 24259
rect 27252 24216 27304 24225
rect 27712 24216 27764 24268
rect 32772 24216 32824 24268
rect 27896 24191 27948 24200
rect 27896 24157 27905 24191
rect 27905 24157 27939 24191
rect 27939 24157 27948 24191
rect 27896 24148 27948 24157
rect 30104 24191 30156 24200
rect 30104 24157 30113 24191
rect 30113 24157 30147 24191
rect 30147 24157 30156 24191
rect 30104 24148 30156 24157
rect 30288 24191 30340 24200
rect 30288 24157 30297 24191
rect 30297 24157 30331 24191
rect 30331 24157 30340 24191
rect 30288 24148 30340 24157
rect 17132 24012 17184 24064
rect 17500 24012 17552 24064
rect 22284 24080 22336 24132
rect 19432 24012 19484 24064
rect 22928 24123 22980 24132
rect 22928 24089 22937 24123
rect 22937 24089 22971 24123
rect 22971 24089 22980 24123
rect 26516 24123 26568 24132
rect 22928 24080 22980 24089
rect 26516 24089 26525 24123
rect 26525 24089 26559 24123
rect 26559 24089 26568 24123
rect 27068 24123 27120 24132
rect 26516 24080 26568 24089
rect 27068 24089 27077 24123
rect 27077 24089 27111 24123
rect 27111 24089 27120 24123
rect 27068 24080 27120 24089
rect 27620 24080 27672 24132
rect 27804 24080 27856 24132
rect 28540 24080 28592 24132
rect 31760 24148 31812 24200
rect 31944 24148 31996 24200
rect 33140 24191 33192 24200
rect 33140 24157 33149 24191
rect 33149 24157 33183 24191
rect 33183 24157 33192 24191
rect 33140 24148 33192 24157
rect 36728 24216 36780 24268
rect 39028 24216 39080 24268
rect 33048 24080 33100 24132
rect 38660 24148 38712 24200
rect 58164 24191 58216 24200
rect 58164 24157 58173 24191
rect 58173 24157 58207 24191
rect 58207 24157 58216 24191
rect 58164 24148 58216 24157
rect 33508 24080 33560 24132
rect 29828 24012 29880 24064
rect 37464 24055 37516 24064
rect 37464 24021 37473 24055
rect 37473 24021 37507 24055
rect 37507 24021 37516 24055
rect 37464 24012 37516 24021
rect 37924 24012 37976 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 11152 23808 11204 23860
rect 11612 23808 11664 23860
rect 3792 23740 3844 23792
rect 6276 23740 6328 23792
rect 1860 23672 1912 23724
rect 3424 23672 3476 23724
rect 5816 23715 5868 23724
rect 5816 23681 5825 23715
rect 5825 23681 5859 23715
rect 5859 23681 5868 23715
rect 5816 23672 5868 23681
rect 14096 23808 14148 23860
rect 11796 23740 11848 23792
rect 12992 23740 13044 23792
rect 6368 23604 6420 23656
rect 6920 23647 6972 23656
rect 6920 23613 6929 23647
rect 6929 23613 6963 23647
rect 6963 23613 6972 23647
rect 6920 23604 6972 23613
rect 10324 23715 10376 23724
rect 10324 23681 10333 23715
rect 10333 23681 10367 23715
rect 10367 23681 10376 23715
rect 10324 23672 10376 23681
rect 11704 23672 11756 23724
rect 13820 23672 13872 23724
rect 14740 23808 14792 23860
rect 14372 23783 14424 23792
rect 14372 23749 14381 23783
rect 14381 23749 14415 23783
rect 14415 23749 14424 23783
rect 15476 23783 15528 23792
rect 14372 23740 14424 23749
rect 10416 23604 10468 23656
rect 15476 23749 15485 23783
rect 15485 23749 15519 23783
rect 15519 23749 15528 23783
rect 15476 23740 15528 23749
rect 15200 23715 15252 23724
rect 15200 23681 15209 23715
rect 15209 23681 15243 23715
rect 15243 23681 15252 23715
rect 15200 23672 15252 23681
rect 17500 23808 17552 23860
rect 17592 23808 17644 23860
rect 20260 23808 20312 23860
rect 21548 23808 21600 23860
rect 21732 23808 21784 23860
rect 15660 23740 15712 23792
rect 16120 23740 16172 23792
rect 19064 23740 19116 23792
rect 20168 23740 20220 23792
rect 20444 23740 20496 23792
rect 3332 23536 3384 23588
rect 7472 23536 7524 23588
rect 3148 23511 3200 23520
rect 3148 23477 3157 23511
rect 3157 23477 3191 23511
rect 3191 23477 3200 23511
rect 3148 23468 3200 23477
rect 15016 23604 15068 23656
rect 18972 23672 19024 23724
rect 23388 23740 23440 23792
rect 30288 23808 30340 23860
rect 27344 23740 27396 23792
rect 29828 23783 29880 23792
rect 29828 23749 29837 23783
rect 29837 23749 29871 23783
rect 29871 23749 29880 23783
rect 29828 23740 29880 23749
rect 35716 23740 35768 23792
rect 18880 23604 18932 23656
rect 14096 23511 14148 23520
rect 14096 23477 14105 23511
rect 14105 23477 14139 23511
rect 14139 23477 14148 23511
rect 14096 23468 14148 23477
rect 15476 23468 15528 23520
rect 18328 23511 18380 23520
rect 18328 23477 18337 23511
rect 18337 23477 18371 23511
rect 18371 23477 18380 23511
rect 18328 23468 18380 23477
rect 19156 23536 19208 23588
rect 21456 23672 21508 23724
rect 21548 23672 21600 23724
rect 24400 23672 24452 23724
rect 27620 23672 27672 23724
rect 28908 23672 28960 23724
rect 33232 23672 33284 23724
rect 36728 23672 36780 23724
rect 38200 23715 38252 23724
rect 38200 23681 38234 23715
rect 38234 23681 38252 23715
rect 38200 23672 38252 23681
rect 24492 23604 24544 23656
rect 37924 23647 37976 23656
rect 37924 23613 37933 23647
rect 37933 23613 37967 23647
rect 37967 23613 37976 23647
rect 37924 23604 37976 23613
rect 22100 23536 22152 23588
rect 26516 23536 26568 23588
rect 31944 23536 31996 23588
rect 22468 23468 22520 23520
rect 28172 23468 28224 23520
rect 32312 23468 32364 23520
rect 37648 23468 37700 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2688 23196 2740 23248
rect 4712 23196 4764 23248
rect 3608 23128 3660 23180
rect 6920 23264 6972 23316
rect 12624 23307 12676 23316
rect 12624 23273 12633 23307
rect 12633 23273 12667 23307
rect 12667 23273 12676 23307
rect 12624 23264 12676 23273
rect 15016 23307 15068 23316
rect 15016 23273 15025 23307
rect 15025 23273 15059 23307
rect 15059 23273 15068 23307
rect 15016 23264 15068 23273
rect 7288 23196 7340 23248
rect 12164 23196 12216 23248
rect 3516 23060 3568 23112
rect 5448 23128 5500 23180
rect 5540 23128 5592 23180
rect 15200 23196 15252 23248
rect 3148 22992 3200 23044
rect 2688 22924 2740 22976
rect 6276 22992 6328 23044
rect 9772 23060 9824 23112
rect 6368 22924 6420 22976
rect 11244 22924 11296 22976
rect 11612 23103 11664 23112
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 11796 23060 11848 23112
rect 15936 23196 15988 23248
rect 22928 23264 22980 23316
rect 24492 23307 24544 23316
rect 24492 23273 24501 23307
rect 24501 23273 24535 23307
rect 24535 23273 24544 23307
rect 24492 23264 24544 23273
rect 25044 23264 25096 23316
rect 21272 23196 21324 23248
rect 23112 23196 23164 23248
rect 11704 23035 11756 23044
rect 11704 23001 11713 23035
rect 11713 23001 11747 23035
rect 11747 23001 11756 23035
rect 11704 22992 11756 23001
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15660 23103 15712 23112
rect 15476 23060 15528 23069
rect 15660 23069 15667 23103
rect 15667 23069 15712 23103
rect 15660 23060 15712 23069
rect 19156 23128 19208 23180
rect 20260 23128 20312 23180
rect 29552 23264 29604 23316
rect 33140 23264 33192 23316
rect 38200 23264 38252 23316
rect 33232 23196 33284 23248
rect 17408 23103 17460 23112
rect 12164 22992 12216 23044
rect 14188 22992 14240 23044
rect 15844 23035 15896 23044
rect 15844 23001 15853 23035
rect 15853 23001 15887 23035
rect 15887 23001 15896 23035
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 17776 23060 17828 23112
rect 28816 23128 28868 23180
rect 32772 23128 32824 23180
rect 15844 22992 15896 23001
rect 19984 22992 20036 23044
rect 20260 22992 20312 23044
rect 20444 22992 20496 23044
rect 20536 22992 20588 23044
rect 20904 22992 20956 23044
rect 16120 22967 16172 22976
rect 16120 22933 16129 22967
rect 16129 22933 16163 22967
rect 16163 22933 16172 22967
rect 16120 22924 16172 22933
rect 17224 22924 17276 22976
rect 22376 22924 22428 22976
rect 30748 23060 30800 23112
rect 31944 23060 31996 23112
rect 32128 23060 32180 23112
rect 33324 23103 33376 23112
rect 27712 22992 27764 23044
rect 31668 22992 31720 23044
rect 27344 22967 27396 22976
rect 27344 22933 27353 22967
rect 27353 22933 27387 22967
rect 27387 22933 27396 22967
rect 27344 22924 27396 22933
rect 30288 22924 30340 22976
rect 33324 23069 33333 23103
rect 33333 23069 33367 23103
rect 33367 23069 33376 23103
rect 33324 23060 33376 23069
rect 33876 23060 33928 23112
rect 37924 23128 37976 23180
rect 32496 22992 32548 23044
rect 33692 22992 33744 23044
rect 34704 22967 34756 22976
rect 34704 22933 34713 22967
rect 34713 22933 34747 22967
rect 34747 22933 34756 22967
rect 34704 22924 34756 22933
rect 37372 23060 37424 23112
rect 37648 23103 37700 23112
rect 37648 23069 37657 23103
rect 37657 23069 37691 23103
rect 37691 23069 37700 23103
rect 37648 23060 37700 23069
rect 37556 22992 37608 23044
rect 39672 23060 39724 23112
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 3608 22652 3660 22704
rect 3332 22627 3384 22636
rect 3332 22593 3341 22627
rect 3341 22593 3375 22627
rect 3375 22593 3384 22627
rect 3332 22584 3384 22593
rect 3516 22627 3568 22636
rect 3516 22593 3525 22627
rect 3525 22593 3559 22627
rect 3559 22593 3568 22627
rect 3516 22584 3568 22593
rect 3700 22516 3752 22568
rect 3884 22516 3936 22568
rect 4712 22584 4764 22636
rect 4988 22584 5040 22636
rect 6276 22720 6328 22772
rect 9312 22652 9364 22704
rect 10324 22720 10376 22772
rect 15200 22720 15252 22772
rect 17408 22720 17460 22772
rect 9864 22652 9916 22704
rect 6368 22627 6420 22636
rect 4068 22448 4120 22500
rect 6368 22593 6377 22627
rect 6377 22593 6411 22627
rect 6411 22593 6420 22627
rect 6368 22584 6420 22593
rect 7104 22584 7156 22636
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 11520 22584 11572 22636
rect 16120 22584 16172 22636
rect 6920 22516 6972 22568
rect 7472 22516 7524 22568
rect 12256 22516 12308 22568
rect 17224 22516 17276 22568
rect 13912 22448 13964 22500
rect 27344 22720 27396 22772
rect 27712 22763 27764 22772
rect 27712 22729 27721 22763
rect 27721 22729 27755 22763
rect 27755 22729 27764 22763
rect 27712 22720 27764 22729
rect 29276 22720 29328 22772
rect 32128 22763 32180 22772
rect 22100 22695 22152 22704
rect 22100 22661 22134 22695
rect 22134 22661 22152 22695
rect 22100 22652 22152 22661
rect 20444 22627 20496 22636
rect 20444 22593 20448 22627
rect 20448 22593 20482 22627
rect 20482 22593 20496 22627
rect 20444 22584 20496 22593
rect 20536 22516 20588 22568
rect 20720 22627 20772 22636
rect 20720 22593 20765 22627
rect 20765 22593 20772 22627
rect 20720 22584 20772 22593
rect 20996 22584 21048 22636
rect 21640 22584 21692 22636
rect 23848 22627 23900 22636
rect 23848 22593 23857 22627
rect 23857 22593 23891 22627
rect 23891 22593 23900 22627
rect 23848 22584 23900 22593
rect 24768 22652 24820 22704
rect 26332 22652 26384 22704
rect 32128 22729 32137 22763
rect 32137 22729 32171 22763
rect 32171 22729 32180 22763
rect 32128 22720 32180 22729
rect 33692 22763 33744 22772
rect 33692 22729 33701 22763
rect 33701 22729 33735 22763
rect 33735 22729 33744 22763
rect 33692 22720 33744 22729
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 25044 22627 25096 22636
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 26056 22584 26108 22636
rect 2964 22380 3016 22432
rect 4620 22423 4672 22432
rect 4620 22389 4629 22423
rect 4629 22389 4663 22423
rect 4663 22389 4672 22423
rect 4620 22380 4672 22389
rect 7012 22423 7064 22432
rect 7012 22389 7021 22423
rect 7021 22389 7055 22423
rect 7055 22389 7064 22423
rect 7012 22380 7064 22389
rect 7104 22380 7156 22432
rect 7564 22423 7616 22432
rect 7564 22389 7573 22423
rect 7573 22389 7607 22423
rect 7607 22389 7616 22423
rect 7564 22380 7616 22389
rect 9956 22423 10008 22432
rect 9956 22389 9965 22423
rect 9965 22389 9999 22423
rect 9999 22389 10008 22423
rect 9956 22380 10008 22389
rect 16120 22380 16172 22432
rect 18880 22380 18932 22432
rect 19248 22423 19300 22432
rect 19248 22389 19257 22423
rect 19257 22389 19291 22423
rect 19291 22389 19300 22423
rect 19248 22380 19300 22389
rect 20076 22380 20128 22432
rect 20352 22380 20404 22432
rect 23388 22380 23440 22432
rect 24952 22448 25004 22500
rect 25044 22448 25096 22500
rect 27068 22448 27120 22500
rect 27528 22448 27580 22500
rect 25136 22380 25188 22432
rect 25320 22423 25372 22432
rect 25320 22389 25329 22423
rect 25329 22389 25363 22423
rect 25363 22389 25372 22423
rect 25320 22380 25372 22389
rect 27344 22380 27396 22432
rect 27804 22516 27856 22568
rect 28172 22627 28224 22636
rect 28172 22593 28181 22627
rect 28181 22593 28215 22627
rect 28215 22593 28224 22627
rect 28172 22584 28224 22593
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 32036 22652 32088 22704
rect 32312 22695 32364 22704
rect 32312 22661 32321 22695
rect 32321 22661 32355 22695
rect 32355 22661 32364 22695
rect 32312 22652 32364 22661
rect 32496 22695 32548 22704
rect 32496 22661 32505 22695
rect 32505 22661 32539 22695
rect 32539 22661 32548 22695
rect 32496 22652 32548 22661
rect 33140 22652 33192 22704
rect 31944 22584 31996 22636
rect 33232 22627 33284 22636
rect 33232 22593 33241 22627
rect 33241 22593 33275 22627
rect 33275 22593 33284 22627
rect 33232 22584 33284 22593
rect 33508 22652 33560 22704
rect 29276 22448 29328 22500
rect 30288 22491 30340 22500
rect 30288 22457 30297 22491
rect 30297 22457 30331 22491
rect 30331 22457 30340 22491
rect 30288 22448 30340 22457
rect 31668 22448 31720 22500
rect 33140 22448 33192 22500
rect 37924 22584 37976 22636
rect 39856 22584 39908 22636
rect 33508 22448 33560 22500
rect 40132 22448 40184 22500
rect 58164 22491 58216 22500
rect 58164 22457 58173 22491
rect 58173 22457 58207 22491
rect 58207 22457 58216 22491
rect 58164 22448 58216 22457
rect 38660 22380 38712 22432
rect 40224 22380 40276 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 4068 22176 4120 22228
rect 5540 22176 5592 22228
rect 6736 22176 6788 22228
rect 7288 22176 7340 22228
rect 7472 22219 7524 22228
rect 7472 22185 7481 22219
rect 7481 22185 7515 22219
rect 7515 22185 7524 22219
rect 7472 22176 7524 22185
rect 14648 22176 14700 22228
rect 15660 22219 15712 22228
rect 15660 22185 15669 22219
rect 15669 22185 15703 22219
rect 15703 22185 15712 22219
rect 15660 22176 15712 22185
rect 16948 22176 17000 22228
rect 17132 22176 17184 22228
rect 18512 22219 18564 22228
rect 18512 22185 18521 22219
rect 18521 22185 18555 22219
rect 18555 22185 18564 22219
rect 18512 22176 18564 22185
rect 18788 22176 18840 22228
rect 22468 22176 22520 22228
rect 21272 22108 21324 22160
rect 26332 22151 26384 22160
rect 26332 22117 26341 22151
rect 26341 22117 26375 22151
rect 26375 22117 26384 22151
rect 26332 22108 26384 22117
rect 27068 22108 27120 22160
rect 28356 22176 28408 22228
rect 39856 22219 39908 22228
rect 39856 22185 39865 22219
rect 39865 22185 39899 22219
rect 39899 22185 39908 22219
rect 39856 22176 39908 22185
rect 29368 22108 29420 22160
rect 29552 22151 29604 22160
rect 29552 22117 29561 22151
rect 29561 22117 29595 22151
rect 29595 22117 29604 22151
rect 29552 22108 29604 22117
rect 13820 22040 13872 22092
rect 2964 22015 3016 22024
rect 2964 21981 2982 22015
rect 2982 21981 3016 22015
rect 2964 21972 3016 21981
rect 4252 21972 4304 22024
rect 7748 21972 7800 22024
rect 3792 21947 3844 21956
rect 3792 21913 3801 21947
rect 3801 21913 3835 21947
rect 3835 21913 3844 21947
rect 3792 21904 3844 21913
rect 3976 21947 4028 21956
rect 3976 21913 3985 21947
rect 3985 21913 4019 21947
rect 4019 21913 4028 21947
rect 3976 21904 4028 21913
rect 1860 21879 1912 21888
rect 1860 21845 1869 21879
rect 1869 21845 1903 21879
rect 1903 21845 1912 21879
rect 1860 21836 1912 21845
rect 3424 21836 3476 21888
rect 3884 21836 3936 21888
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 7012 21904 7064 21956
rect 9312 21972 9364 22024
rect 9772 21972 9824 22024
rect 20536 22040 20588 22092
rect 22008 22040 22060 22092
rect 18144 21972 18196 22024
rect 18604 22015 18656 22024
rect 18604 21981 18613 22015
rect 18613 21981 18647 22015
rect 18647 21981 18656 22015
rect 18604 21972 18656 21981
rect 9680 21904 9732 21956
rect 14556 21947 14608 21956
rect 14556 21913 14590 21947
rect 14590 21913 14608 21947
rect 16120 21947 16172 21956
rect 14556 21904 14608 21913
rect 16120 21913 16129 21947
rect 16129 21913 16163 21947
rect 16163 21913 16172 21947
rect 16120 21904 16172 21913
rect 22192 21972 22244 22024
rect 26240 21972 26292 22024
rect 29920 22040 29972 22092
rect 33600 22108 33652 22160
rect 30380 22040 30432 22092
rect 31024 22040 31076 22092
rect 33232 22040 33284 22092
rect 19432 21904 19484 21956
rect 9772 21879 9824 21888
rect 9772 21845 9781 21879
rect 9781 21845 9815 21879
rect 9815 21845 9824 21879
rect 9772 21836 9824 21845
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 18328 21836 18380 21845
rect 18788 21836 18840 21888
rect 19984 21836 20036 21888
rect 20904 21879 20956 21888
rect 20904 21845 20913 21879
rect 20913 21845 20947 21879
rect 20947 21845 20956 21879
rect 20904 21836 20956 21845
rect 23388 21836 23440 21888
rect 25504 21904 25556 21956
rect 26700 21904 26752 21956
rect 28264 21904 28316 21956
rect 29184 21904 29236 21956
rect 30656 21972 30708 22024
rect 31116 21972 31168 22024
rect 34704 21972 34756 22024
rect 35900 22040 35952 22092
rect 37740 22040 37792 22092
rect 38844 21972 38896 22024
rect 39120 22108 39172 22160
rect 39856 21972 39908 22024
rect 40132 22015 40184 22024
rect 40132 21981 40141 22015
rect 40141 21981 40175 22015
rect 40175 21981 40184 22015
rect 40132 21972 40184 21981
rect 32588 21947 32640 21956
rect 23848 21836 23900 21888
rect 26608 21836 26660 21888
rect 28080 21836 28132 21888
rect 32588 21913 32597 21947
rect 32597 21913 32631 21947
rect 32631 21913 32640 21947
rect 32588 21904 32640 21913
rect 31944 21836 31996 21888
rect 33324 21836 33376 21888
rect 33508 21879 33560 21888
rect 33508 21845 33517 21879
rect 33517 21845 33551 21879
rect 33551 21845 33560 21879
rect 33508 21836 33560 21845
rect 35624 21879 35676 21888
rect 35624 21845 35633 21879
rect 35633 21845 35667 21879
rect 35667 21845 35676 21879
rect 35624 21836 35676 21845
rect 35992 21947 36044 21956
rect 35992 21913 36001 21947
rect 36001 21913 36035 21947
rect 36035 21913 36044 21947
rect 35992 21904 36044 21913
rect 38752 21904 38804 21956
rect 40316 22015 40368 22024
rect 40316 21981 40325 22015
rect 40325 21981 40359 22015
rect 40359 21981 40368 22015
rect 40316 21972 40368 21981
rect 40500 22015 40552 22024
rect 40500 21981 40509 22015
rect 40509 21981 40543 22015
rect 40543 21981 40552 22015
rect 40500 21972 40552 21981
rect 40684 21904 40736 21956
rect 40960 21947 41012 21956
rect 40960 21913 40969 21947
rect 40969 21913 41003 21947
rect 41003 21913 41012 21947
rect 40960 21904 41012 21913
rect 41144 21947 41196 21956
rect 41144 21913 41153 21947
rect 41153 21913 41187 21947
rect 41187 21913 41196 21947
rect 41144 21904 41196 21913
rect 37188 21879 37240 21888
rect 37188 21845 37197 21879
rect 37197 21845 37231 21879
rect 37231 21845 37240 21879
rect 37188 21836 37240 21845
rect 38660 21879 38712 21888
rect 38660 21845 38669 21879
rect 38669 21845 38703 21879
rect 38703 21845 38712 21879
rect 38660 21836 38712 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 3884 21632 3936 21684
rect 3976 21632 4028 21684
rect 9404 21632 9456 21684
rect 4620 21564 4672 21616
rect 6736 21607 6788 21616
rect 6736 21573 6745 21607
rect 6745 21573 6779 21607
rect 6779 21573 6788 21607
rect 6736 21564 6788 21573
rect 7932 21564 7984 21616
rect 12164 21564 12216 21616
rect 14280 21632 14332 21684
rect 14556 21675 14608 21684
rect 14556 21641 14565 21675
rect 14565 21641 14599 21675
rect 14599 21641 14608 21675
rect 14556 21632 14608 21641
rect 12808 21564 12860 21616
rect 18236 21632 18288 21684
rect 2688 21539 2740 21548
rect 2688 21505 2722 21539
rect 2722 21505 2740 21539
rect 2688 21496 2740 21505
rect 4252 21539 4304 21548
rect 4252 21505 4261 21539
rect 4261 21505 4295 21539
rect 4295 21505 4304 21539
rect 4252 21496 4304 21505
rect 10140 21496 10192 21548
rect 13912 21539 13964 21548
rect 13912 21505 13921 21539
rect 13921 21505 13955 21539
rect 13955 21505 13964 21539
rect 13912 21496 13964 21505
rect 14096 21539 14148 21548
rect 14096 21505 14105 21539
rect 14105 21505 14139 21539
rect 14139 21505 14148 21539
rect 14096 21496 14148 21505
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 15200 21539 15252 21548
rect 7748 21428 7800 21480
rect 15200 21505 15209 21539
rect 15209 21505 15243 21539
rect 15243 21505 15252 21539
rect 15200 21496 15252 21505
rect 16948 21496 17000 21548
rect 17868 21539 17920 21548
rect 17868 21505 17877 21539
rect 17877 21505 17911 21539
rect 17911 21505 17920 21539
rect 17868 21496 17920 21505
rect 18032 21539 18084 21548
rect 18032 21505 18040 21539
rect 18040 21505 18074 21539
rect 18074 21505 18084 21539
rect 18032 21496 18084 21505
rect 11612 21403 11664 21412
rect 11612 21369 11621 21403
rect 11621 21369 11655 21403
rect 11655 21369 11664 21403
rect 11612 21360 11664 21369
rect 12808 21360 12860 21412
rect 14924 21428 14976 21480
rect 11336 21292 11388 21344
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 13360 21335 13412 21344
rect 13360 21301 13369 21335
rect 13369 21301 13403 21335
rect 13403 21301 13412 21335
rect 13360 21292 13412 21301
rect 15752 21292 15804 21344
rect 17776 21428 17828 21480
rect 18236 21539 18288 21548
rect 18236 21505 18245 21539
rect 18245 21505 18279 21539
rect 18279 21505 18288 21539
rect 18972 21539 19024 21548
rect 18236 21496 18288 21505
rect 18972 21505 18981 21539
rect 18981 21505 19015 21539
rect 19015 21505 19024 21539
rect 18972 21496 19024 21505
rect 20536 21496 20588 21548
rect 18604 21428 18656 21480
rect 19984 21428 20036 21480
rect 21272 21564 21324 21616
rect 22008 21564 22060 21616
rect 24860 21632 24912 21684
rect 25504 21675 25556 21684
rect 25504 21641 25513 21675
rect 25513 21641 25547 21675
rect 25547 21641 25556 21675
rect 25504 21632 25556 21641
rect 27344 21675 27396 21684
rect 27344 21641 27353 21675
rect 27353 21641 27387 21675
rect 27387 21641 27396 21675
rect 27344 21632 27396 21641
rect 26056 21564 26108 21616
rect 29000 21632 29052 21684
rect 29368 21675 29420 21684
rect 29368 21641 29377 21675
rect 29377 21641 29411 21675
rect 29411 21641 29420 21675
rect 29368 21632 29420 21641
rect 31944 21632 31996 21684
rect 32128 21675 32180 21684
rect 32128 21641 32137 21675
rect 32137 21641 32171 21675
rect 32171 21641 32180 21675
rect 32128 21632 32180 21641
rect 33508 21632 33560 21684
rect 36452 21632 36504 21684
rect 30196 21564 30248 21616
rect 30288 21564 30340 21616
rect 32036 21564 32088 21616
rect 32220 21564 32272 21616
rect 25044 21539 25096 21548
rect 20812 21428 20864 21480
rect 21732 21428 21784 21480
rect 25044 21505 25053 21539
rect 25053 21505 25087 21539
rect 25087 21505 25096 21539
rect 25044 21496 25096 21505
rect 18236 21360 18288 21412
rect 23480 21428 23532 21480
rect 24952 21428 25004 21480
rect 25228 21539 25280 21548
rect 25228 21505 25237 21539
rect 25237 21505 25271 21539
rect 25271 21505 25280 21539
rect 25228 21496 25280 21505
rect 25596 21496 25648 21548
rect 26608 21496 26660 21548
rect 27436 21496 27488 21548
rect 26976 21428 27028 21480
rect 28172 21428 28224 21480
rect 25780 21360 25832 21412
rect 28540 21360 28592 21412
rect 29736 21496 29788 21548
rect 31116 21496 31168 21548
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 37188 21496 37240 21548
rect 39120 21632 39172 21684
rect 40684 21632 40736 21684
rect 38660 21564 38712 21616
rect 39764 21564 39816 21616
rect 40960 21564 41012 21616
rect 37740 21539 37792 21548
rect 37740 21505 37749 21539
rect 37749 21505 37783 21539
rect 37783 21505 37792 21539
rect 37740 21496 37792 21505
rect 30012 21428 30064 21480
rect 32036 21428 32088 21480
rect 35348 21471 35400 21480
rect 35348 21437 35357 21471
rect 35357 21437 35391 21471
rect 35391 21437 35400 21471
rect 35348 21428 35400 21437
rect 36544 21428 36596 21480
rect 40040 21496 40092 21548
rect 40408 21496 40460 21548
rect 40592 21496 40644 21548
rect 17960 21292 18012 21344
rect 18512 21335 18564 21344
rect 18512 21301 18521 21335
rect 18521 21301 18555 21335
rect 18555 21301 18564 21335
rect 18512 21292 18564 21301
rect 22468 21292 22520 21344
rect 32220 21292 32272 21344
rect 36912 21292 36964 21344
rect 40040 21292 40092 21344
rect 40132 21335 40184 21344
rect 40132 21301 40141 21335
rect 40141 21301 40175 21335
rect 40175 21301 40184 21335
rect 40132 21292 40184 21301
rect 41144 21292 41196 21344
rect 58164 21335 58216 21344
rect 58164 21301 58173 21335
rect 58173 21301 58207 21335
rect 58207 21301 58216 21335
rect 58164 21292 58216 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 10140 21131 10192 21140
rect 10140 21097 10149 21131
rect 10149 21097 10183 21131
rect 10183 21097 10192 21131
rect 10140 21088 10192 21097
rect 1860 21020 1912 21072
rect 11796 21088 11848 21140
rect 14096 21088 14148 21140
rect 18052 21088 18104 21140
rect 18144 21088 18196 21140
rect 25136 21131 25188 21140
rect 10508 21020 10560 21072
rect 16948 21020 17000 21072
rect 18972 21020 19024 21072
rect 10232 20952 10284 21004
rect 13176 20952 13228 21004
rect 14188 20952 14240 21004
rect 9680 20927 9732 20936
rect 9680 20893 9689 20927
rect 9689 20893 9723 20927
rect 9723 20893 9732 20927
rect 9680 20884 9732 20893
rect 10508 20927 10560 20936
rect 10508 20893 10517 20927
rect 10517 20893 10551 20927
rect 10551 20893 10560 20927
rect 10508 20884 10560 20893
rect 6920 20816 6972 20868
rect 7748 20816 7800 20868
rect 10784 20927 10836 20936
rect 10784 20893 10793 20927
rect 10793 20893 10827 20927
rect 10827 20893 10836 20927
rect 10784 20884 10836 20893
rect 11612 20884 11664 20936
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 15660 20884 15712 20936
rect 15752 20927 15804 20936
rect 15752 20893 15761 20927
rect 15761 20893 15795 20927
rect 15795 20893 15804 20927
rect 17776 20952 17828 21004
rect 25136 21097 25145 21131
rect 25145 21097 25179 21131
rect 25179 21097 25188 21131
rect 25136 21088 25188 21097
rect 28356 21131 28408 21140
rect 28356 21097 28365 21131
rect 28365 21097 28399 21131
rect 28399 21097 28408 21131
rect 28356 21088 28408 21097
rect 28540 21088 28592 21140
rect 30196 21088 30248 21140
rect 32312 21088 32364 21140
rect 37740 21088 37792 21140
rect 40500 21088 40552 21140
rect 15752 20884 15804 20893
rect 11152 20816 11204 20868
rect 15292 20816 15344 20868
rect 16948 20816 17000 20868
rect 17868 20884 17920 20936
rect 18236 20927 18288 20936
rect 18236 20893 18245 20927
rect 18245 20893 18279 20927
rect 18279 20893 18288 20927
rect 18236 20884 18288 20893
rect 21088 20884 21140 20936
rect 21272 20927 21324 20936
rect 21272 20893 21281 20927
rect 21281 20893 21315 20927
rect 21315 20893 21324 20927
rect 21272 20884 21324 20893
rect 22284 21020 22336 21072
rect 25596 21020 25648 21072
rect 26976 21063 27028 21072
rect 26976 21029 26985 21063
rect 26985 21029 27019 21063
rect 27019 21029 27028 21063
rect 26976 21020 27028 21029
rect 21732 20952 21784 21004
rect 22100 20884 22152 20936
rect 22468 20884 22520 20936
rect 24124 20884 24176 20936
rect 26240 20884 26292 20936
rect 27068 20884 27120 20936
rect 28080 20927 28132 20936
rect 28080 20893 28089 20927
rect 28089 20893 28123 20927
rect 28123 20893 28132 20927
rect 28080 20884 28132 20893
rect 28172 20927 28224 20936
rect 28172 20893 28181 20927
rect 28181 20893 28215 20927
rect 28215 20893 28224 20927
rect 30104 21020 30156 21072
rect 31116 21020 31168 21072
rect 31944 21063 31996 21072
rect 31944 21029 31953 21063
rect 31953 21029 31987 21063
rect 31987 21029 31996 21063
rect 31944 21020 31996 21029
rect 32220 21020 32272 21072
rect 34796 21020 34848 21072
rect 28172 20884 28224 20893
rect 25872 20859 25924 20868
rect 25872 20825 25884 20859
rect 25884 20825 25924 20859
rect 7932 20791 7984 20800
rect 7932 20757 7941 20791
rect 7941 20757 7975 20791
rect 7975 20757 7984 20791
rect 7932 20748 7984 20757
rect 10416 20748 10468 20800
rect 17316 20748 17368 20800
rect 25872 20816 25924 20825
rect 29000 20816 29052 20868
rect 30288 20952 30340 21004
rect 30104 20927 30156 20936
rect 30104 20893 30113 20927
rect 30113 20893 30147 20927
rect 30147 20893 30156 20927
rect 30104 20884 30156 20893
rect 30196 20884 30248 20936
rect 31116 20927 31168 20936
rect 31116 20893 31125 20927
rect 31125 20893 31159 20927
rect 31159 20893 31168 20927
rect 31116 20884 31168 20893
rect 35624 20952 35676 21004
rect 32220 20927 32272 20936
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 35900 21020 35952 21072
rect 40132 20952 40184 21004
rect 32220 20884 32272 20893
rect 35992 20927 36044 20936
rect 35992 20893 36001 20927
rect 36001 20893 36035 20927
rect 36035 20893 36044 20927
rect 35992 20884 36044 20893
rect 38936 20884 38988 20936
rect 40224 20884 40276 20936
rect 30840 20816 30892 20868
rect 31760 20816 31812 20868
rect 31852 20816 31904 20868
rect 36912 20859 36964 20868
rect 36912 20825 36921 20859
rect 36921 20825 36955 20859
rect 36955 20825 36964 20859
rect 36912 20816 36964 20825
rect 39764 20816 39816 20868
rect 19340 20748 19392 20800
rect 20536 20748 20588 20800
rect 22192 20748 22244 20800
rect 23940 20748 23992 20800
rect 29736 20748 29788 20800
rect 32312 20748 32364 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 6920 20544 6972 20596
rect 10508 20544 10560 20596
rect 11152 20544 11204 20596
rect 14096 20544 14148 20596
rect 17316 20544 17368 20596
rect 19340 20544 19392 20596
rect 21272 20544 21324 20596
rect 6644 20476 6696 20528
rect 7104 20451 7156 20460
rect 7104 20417 7113 20451
rect 7113 20417 7147 20451
rect 7147 20417 7156 20451
rect 7104 20408 7156 20417
rect 10324 20408 10376 20460
rect 11336 20476 11388 20528
rect 12808 20519 12860 20528
rect 12808 20485 12817 20519
rect 12817 20485 12851 20519
rect 12851 20485 12860 20519
rect 12808 20476 12860 20485
rect 13084 20476 13136 20528
rect 13912 20476 13964 20528
rect 18512 20476 18564 20528
rect 21088 20519 21140 20528
rect 21088 20485 21097 20519
rect 21097 20485 21131 20519
rect 21131 20485 21140 20519
rect 21088 20476 21140 20485
rect 7748 20340 7800 20392
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 10600 20272 10652 20324
rect 13268 20408 13320 20460
rect 14188 20408 14240 20460
rect 14740 20451 14792 20460
rect 14740 20417 14749 20451
rect 14749 20417 14783 20451
rect 14783 20417 14792 20451
rect 14740 20408 14792 20417
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 22192 20519 22244 20528
rect 22192 20485 22226 20519
rect 22226 20485 22244 20519
rect 22192 20476 22244 20485
rect 23480 20476 23532 20528
rect 23940 20451 23992 20460
rect 23940 20417 23949 20451
rect 23949 20417 23983 20451
rect 23983 20417 23992 20451
rect 23940 20408 23992 20417
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 29552 20476 29604 20528
rect 30104 20476 30156 20528
rect 31576 20476 31628 20528
rect 29736 20408 29788 20460
rect 32864 20476 32916 20528
rect 36912 20476 36964 20528
rect 35900 20451 35952 20460
rect 12808 20272 12860 20324
rect 15752 20272 15804 20324
rect 10140 20204 10192 20256
rect 14280 20204 14332 20256
rect 14464 20204 14516 20256
rect 28172 20340 28224 20392
rect 29000 20340 29052 20392
rect 35900 20417 35909 20451
rect 35909 20417 35943 20451
rect 35943 20417 35952 20451
rect 35900 20408 35952 20417
rect 36084 20451 36136 20460
rect 36084 20417 36093 20451
rect 36093 20417 36127 20451
rect 36127 20417 36136 20451
rect 36084 20408 36136 20417
rect 36636 20408 36688 20460
rect 36452 20272 36504 20324
rect 36636 20272 36688 20324
rect 22100 20204 22152 20256
rect 23756 20204 23808 20256
rect 32312 20247 32364 20256
rect 32312 20213 32321 20247
rect 32321 20213 32355 20247
rect 32355 20213 32364 20247
rect 32312 20204 32364 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 10600 20000 10652 20052
rect 11152 20000 11204 20052
rect 11612 20000 11664 20052
rect 12164 20000 12216 20052
rect 13084 20000 13136 20052
rect 14188 20043 14240 20052
rect 14188 20009 14197 20043
rect 14197 20009 14231 20043
rect 14231 20009 14240 20043
rect 14188 20000 14240 20009
rect 15108 20000 15160 20052
rect 18236 20000 18288 20052
rect 21272 20000 21324 20052
rect 22284 20000 22336 20052
rect 34796 20000 34848 20052
rect 39672 20000 39724 20052
rect 40868 20000 40920 20052
rect 5724 19932 5776 19984
rect 13360 19932 13412 19984
rect 7564 19864 7616 19916
rect 2412 19796 2464 19848
rect 4712 19796 4764 19848
rect 4896 19796 4948 19848
rect 10324 19796 10376 19848
rect 12256 19864 12308 19916
rect 13176 19864 13228 19916
rect 3884 19728 3936 19780
rect 5724 19728 5776 19780
rect 6184 19771 6236 19780
rect 6184 19737 6193 19771
rect 6193 19737 6227 19771
rect 6227 19737 6236 19771
rect 6184 19728 6236 19737
rect 10140 19728 10192 19780
rect 10416 19771 10468 19780
rect 10416 19737 10425 19771
rect 10425 19737 10459 19771
rect 10459 19737 10468 19771
rect 10416 19728 10468 19737
rect 12900 19839 12952 19848
rect 12900 19805 12909 19839
rect 12909 19805 12943 19839
rect 12943 19805 12952 19839
rect 12900 19796 12952 19805
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 26240 19864 26292 19916
rect 13084 19796 13136 19805
rect 15568 19839 15620 19848
rect 15568 19805 15577 19839
rect 15577 19805 15611 19839
rect 15611 19805 15620 19839
rect 15568 19796 15620 19805
rect 2136 19660 2188 19712
rect 7104 19660 7156 19712
rect 12440 19703 12492 19712
rect 12440 19669 12449 19703
rect 12449 19669 12483 19703
rect 12483 19669 12492 19703
rect 13820 19728 13872 19780
rect 15292 19728 15344 19780
rect 16028 19796 16080 19848
rect 23756 19796 23808 19848
rect 30840 19796 30892 19848
rect 31760 19796 31812 19848
rect 32680 19796 32732 19848
rect 36360 19932 36412 19984
rect 36268 19864 36320 19916
rect 35716 19796 35768 19848
rect 58164 19839 58216 19848
rect 58164 19805 58173 19839
rect 58173 19805 58207 19839
rect 58207 19805 58216 19839
rect 58164 19796 58216 19805
rect 16672 19728 16724 19780
rect 20076 19728 20128 19780
rect 24124 19728 24176 19780
rect 27620 19728 27672 19780
rect 31116 19771 31168 19780
rect 31116 19737 31125 19771
rect 31125 19737 31159 19771
rect 31159 19737 31168 19771
rect 32588 19771 32640 19780
rect 31116 19728 31168 19737
rect 32588 19737 32597 19771
rect 32597 19737 32631 19771
rect 32631 19737 32640 19771
rect 32588 19728 32640 19737
rect 12440 19660 12492 19669
rect 17408 19660 17460 19712
rect 30840 19660 30892 19712
rect 32864 19660 32916 19712
rect 38660 19660 38712 19712
rect 39856 19660 39908 19712
rect 41052 19660 41104 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 2412 19499 2464 19508
rect 2412 19465 2421 19499
rect 2421 19465 2455 19499
rect 2455 19465 2464 19499
rect 2412 19456 2464 19465
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 10416 19456 10468 19508
rect 10968 19388 11020 19440
rect 3792 19320 3844 19372
rect 7932 19320 7984 19372
rect 11520 19320 11572 19372
rect 11796 19363 11848 19372
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 12256 19388 12308 19440
rect 12164 19363 12216 19372
rect 2872 19252 2924 19304
rect 3884 19184 3936 19236
rect 4068 19295 4120 19304
rect 4068 19261 4077 19295
rect 4077 19261 4111 19295
rect 4111 19261 4120 19295
rect 4068 19252 4120 19261
rect 2596 19116 2648 19168
rect 4712 19116 4764 19168
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 6184 19116 6236 19168
rect 12164 19329 12173 19363
rect 12173 19329 12207 19363
rect 12207 19329 12216 19363
rect 12164 19320 12216 19329
rect 12900 19456 12952 19508
rect 15568 19456 15620 19508
rect 17776 19456 17828 19508
rect 21732 19456 21784 19508
rect 27712 19456 27764 19508
rect 32680 19456 32732 19508
rect 38660 19456 38712 19508
rect 40500 19456 40552 19508
rect 41052 19499 41104 19508
rect 41052 19465 41061 19499
rect 41061 19465 41095 19499
rect 41095 19465 41104 19499
rect 41052 19456 41104 19465
rect 12808 19320 12860 19372
rect 13084 19320 13136 19372
rect 13820 19320 13872 19372
rect 16764 19388 16816 19440
rect 15568 19363 15620 19372
rect 15568 19329 15577 19363
rect 15577 19329 15611 19363
rect 15611 19329 15620 19363
rect 15568 19320 15620 19329
rect 16028 19320 16080 19372
rect 17592 19388 17644 19440
rect 9496 19184 9548 19236
rect 16488 19252 16540 19304
rect 18052 19320 18104 19372
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18512 19320 18564 19372
rect 20352 19320 20404 19372
rect 29736 19388 29788 19440
rect 29460 19363 29512 19372
rect 29460 19329 29469 19363
rect 29469 19329 29503 19363
rect 29503 19329 29512 19363
rect 29460 19320 29512 19329
rect 29552 19363 29604 19372
rect 29552 19329 29561 19363
rect 29561 19329 29595 19363
rect 29595 19329 29604 19363
rect 29552 19320 29604 19329
rect 30840 19363 30892 19372
rect 30840 19329 30849 19363
rect 30849 19329 30883 19363
rect 30883 19329 30892 19363
rect 30840 19320 30892 19329
rect 17776 19295 17828 19304
rect 17776 19261 17785 19295
rect 17785 19261 17819 19295
rect 17819 19261 17828 19295
rect 17776 19252 17828 19261
rect 8484 19116 8536 19168
rect 8576 19116 8628 19168
rect 10232 19184 10284 19236
rect 30288 19184 30340 19236
rect 31024 19363 31076 19372
rect 31024 19329 31033 19363
rect 31033 19329 31067 19363
rect 31067 19329 31076 19363
rect 31944 19388 31996 19440
rect 39856 19388 39908 19440
rect 31024 19320 31076 19329
rect 32312 19320 32364 19372
rect 33324 19320 33376 19372
rect 35348 19320 35400 19372
rect 35992 19320 36044 19372
rect 40040 19320 40092 19372
rect 40408 19363 40460 19372
rect 40408 19329 40417 19363
rect 40417 19329 40451 19363
rect 40451 19329 40460 19363
rect 40408 19320 40460 19329
rect 32128 19295 32180 19304
rect 32128 19261 32137 19295
rect 32137 19261 32171 19295
rect 32171 19261 32180 19295
rect 32128 19252 32180 19261
rect 36268 19252 36320 19304
rect 40868 19320 40920 19372
rect 31668 19184 31720 19236
rect 40684 19184 40736 19236
rect 11520 19159 11572 19168
rect 11520 19125 11529 19159
rect 11529 19125 11563 19159
rect 11563 19125 11572 19159
rect 11520 19116 11572 19125
rect 15384 19116 15436 19168
rect 17224 19116 17276 19168
rect 18880 19116 18932 19168
rect 19156 19116 19208 19168
rect 25780 19116 25832 19168
rect 29644 19116 29696 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 3792 18955 3844 18964
rect 3792 18921 3801 18955
rect 3801 18921 3835 18955
rect 3835 18921 3844 18955
rect 3792 18912 3844 18921
rect 4068 18912 4120 18964
rect 4252 18819 4304 18828
rect 4252 18785 4261 18819
rect 4261 18785 4295 18819
rect 4295 18785 4304 18819
rect 4252 18776 4304 18785
rect 9036 18912 9088 18964
rect 10232 18955 10284 18964
rect 10232 18921 10241 18955
rect 10241 18921 10275 18955
rect 10275 18921 10284 18955
rect 10232 18912 10284 18921
rect 13084 18912 13136 18964
rect 13360 18912 13412 18964
rect 16948 18912 17000 18964
rect 17500 18912 17552 18964
rect 17776 18912 17828 18964
rect 24308 18912 24360 18964
rect 30932 18912 30984 18964
rect 33324 18955 33376 18964
rect 33324 18921 33333 18955
rect 33333 18921 33367 18955
rect 33367 18921 33376 18955
rect 33324 18912 33376 18921
rect 40500 18912 40552 18964
rect 19984 18844 20036 18896
rect 20444 18844 20496 18896
rect 7748 18819 7800 18828
rect 7748 18785 7757 18819
rect 7757 18785 7791 18819
rect 7791 18785 7800 18819
rect 7748 18776 7800 18785
rect 18880 18776 18932 18828
rect 19248 18819 19300 18828
rect 19248 18785 19257 18819
rect 19257 18785 19291 18819
rect 19291 18785 19300 18819
rect 19248 18776 19300 18785
rect 19340 18776 19392 18828
rect 1860 18751 1912 18760
rect 1860 18717 1869 18751
rect 1869 18717 1903 18751
rect 1903 18717 1912 18751
rect 1860 18708 1912 18717
rect 2136 18751 2188 18760
rect 2136 18717 2170 18751
rect 2170 18717 2188 18751
rect 2136 18708 2188 18717
rect 9588 18708 9640 18760
rect 13544 18708 13596 18760
rect 15384 18708 15436 18760
rect 16488 18708 16540 18760
rect 17408 18751 17460 18760
rect 17408 18717 17442 18751
rect 17442 18717 17460 18751
rect 17408 18708 17460 18717
rect 19984 18751 20036 18760
rect 19984 18717 19988 18751
rect 19988 18717 20022 18751
rect 20022 18717 20036 18751
rect 19984 18708 20036 18717
rect 4712 18640 4764 18692
rect 6828 18640 6880 18692
rect 12440 18683 12492 18692
rect 12440 18649 12474 18683
rect 12474 18649 12492 18683
rect 12440 18640 12492 18649
rect 17592 18640 17644 18692
rect 19340 18640 19392 18692
rect 19892 18640 19944 18692
rect 20996 18708 21048 18760
rect 23940 18708 23992 18760
rect 20260 18640 20312 18692
rect 29000 18844 29052 18896
rect 29552 18844 29604 18896
rect 28172 18776 28224 18828
rect 24768 18751 24820 18760
rect 24768 18717 24777 18751
rect 24777 18717 24811 18751
rect 24811 18717 24820 18751
rect 24768 18708 24820 18717
rect 25780 18708 25832 18760
rect 29736 18751 29788 18760
rect 29736 18717 29745 18751
rect 29745 18717 29779 18751
rect 29779 18717 29788 18751
rect 29736 18708 29788 18717
rect 32772 18776 32824 18828
rect 35348 18776 35400 18828
rect 35900 18776 35952 18828
rect 31944 18751 31996 18760
rect 31944 18717 31962 18751
rect 31962 18717 31996 18751
rect 31944 18708 31996 18717
rect 32312 18708 32364 18760
rect 32864 18751 32916 18760
rect 32864 18717 32873 18751
rect 32873 18717 32907 18751
rect 32907 18717 32916 18751
rect 32864 18708 32916 18717
rect 25044 18640 25096 18692
rect 4160 18615 4212 18624
rect 4160 18581 4169 18615
rect 4169 18581 4203 18615
rect 4203 18581 4212 18615
rect 4160 18572 4212 18581
rect 6184 18572 6236 18624
rect 8392 18572 8444 18624
rect 11060 18572 11112 18624
rect 11796 18572 11848 18624
rect 18236 18572 18288 18624
rect 19156 18572 19208 18624
rect 19432 18572 19484 18624
rect 20996 18572 21048 18624
rect 23664 18615 23716 18624
rect 23664 18581 23673 18615
rect 23673 18581 23707 18615
rect 23707 18581 23716 18615
rect 23664 18572 23716 18581
rect 23940 18572 23992 18624
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 26056 18572 26108 18624
rect 26792 18615 26844 18624
rect 26792 18581 26801 18615
rect 26801 18581 26835 18615
rect 26835 18581 26844 18615
rect 26792 18572 26844 18581
rect 26976 18683 27028 18692
rect 26976 18649 26985 18683
rect 26985 18649 27019 18683
rect 27019 18649 27028 18683
rect 26976 18640 27028 18649
rect 27436 18640 27488 18692
rect 29828 18683 29880 18692
rect 29828 18649 29837 18683
rect 29837 18649 29871 18683
rect 29871 18649 29880 18683
rect 29828 18640 29880 18649
rect 31668 18640 31720 18692
rect 33048 18751 33100 18760
rect 33048 18717 33057 18751
rect 33057 18717 33091 18751
rect 33091 18717 33100 18751
rect 36360 18751 36412 18760
rect 33048 18708 33100 18717
rect 36360 18717 36369 18751
rect 36369 18717 36403 18751
rect 36403 18717 36412 18751
rect 36360 18708 36412 18717
rect 37648 18708 37700 18760
rect 38660 18708 38712 18760
rect 58164 18751 58216 18760
rect 58164 18717 58173 18751
rect 58173 18717 58207 18751
rect 58207 18717 58216 18751
rect 58164 18708 58216 18717
rect 36084 18640 36136 18692
rect 37188 18683 37240 18692
rect 37188 18649 37197 18683
rect 37197 18649 37231 18683
rect 37231 18649 37240 18683
rect 37188 18640 37240 18649
rect 39764 18640 39816 18692
rect 30472 18572 30524 18624
rect 36820 18615 36872 18624
rect 36820 18581 36829 18615
rect 36829 18581 36863 18615
rect 36863 18581 36872 18615
rect 36820 18572 36872 18581
rect 37004 18572 37056 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 4160 18368 4212 18420
rect 6092 18368 6144 18420
rect 6828 18411 6880 18420
rect 6828 18377 6837 18411
rect 6837 18377 6871 18411
rect 6871 18377 6880 18411
rect 6828 18368 6880 18377
rect 10048 18368 10100 18420
rect 12256 18368 12308 18420
rect 16120 18368 16172 18420
rect 16672 18411 16724 18420
rect 16672 18377 16681 18411
rect 16681 18377 16715 18411
rect 16715 18377 16724 18411
rect 16672 18368 16724 18377
rect 17040 18368 17092 18420
rect 17224 18368 17276 18420
rect 18972 18368 19024 18420
rect 1860 18300 1912 18352
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 2780 18300 2832 18352
rect 4252 18232 4304 18284
rect 6184 18232 6236 18284
rect 8576 18300 8628 18352
rect 11520 18300 11572 18352
rect 15568 18300 15620 18352
rect 7932 18232 7984 18284
rect 8392 18275 8444 18284
rect 8392 18241 8401 18275
rect 8401 18241 8435 18275
rect 8435 18241 8444 18275
rect 8392 18232 8444 18241
rect 9312 18232 9364 18284
rect 18604 18300 18656 18352
rect 5172 18164 5224 18216
rect 5540 18207 5592 18216
rect 5540 18173 5549 18207
rect 5549 18173 5583 18207
rect 5583 18173 5592 18207
rect 5540 18164 5592 18173
rect 7104 18164 7156 18216
rect 3792 18071 3844 18080
rect 3792 18037 3801 18071
rect 3801 18037 3835 18071
rect 3835 18037 3844 18071
rect 3792 18028 3844 18037
rect 4620 18028 4672 18080
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 16856 18275 16908 18284
rect 16856 18241 16865 18275
rect 16865 18241 16899 18275
rect 16899 18241 16908 18275
rect 16856 18232 16908 18241
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 17776 18275 17828 18284
rect 17776 18241 17785 18275
rect 17785 18241 17819 18275
rect 17819 18241 17828 18275
rect 17776 18232 17828 18241
rect 19432 18300 19484 18352
rect 20352 18368 20404 18420
rect 20536 18368 20588 18420
rect 24216 18368 24268 18420
rect 25044 18411 25096 18420
rect 25044 18377 25053 18411
rect 25053 18377 25087 18411
rect 25087 18377 25096 18411
rect 25044 18368 25096 18377
rect 19708 18300 19760 18352
rect 19248 18275 19300 18284
rect 16948 18096 17000 18148
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 19984 18232 20036 18284
rect 20260 18275 20312 18284
rect 20260 18241 20269 18275
rect 20269 18241 20303 18275
rect 20303 18241 20312 18275
rect 20260 18232 20312 18241
rect 32588 18411 32640 18420
rect 32588 18377 32597 18411
rect 32597 18377 32631 18411
rect 32631 18377 32640 18411
rect 32588 18368 32640 18377
rect 33048 18368 33100 18420
rect 35348 18368 35400 18420
rect 20628 18275 20680 18284
rect 20628 18241 20637 18275
rect 20637 18241 20671 18275
rect 20671 18241 20680 18275
rect 20628 18232 20680 18241
rect 20812 18164 20864 18216
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 11704 18071 11756 18080
rect 11704 18037 11713 18071
rect 11713 18037 11747 18071
rect 11747 18037 11756 18071
rect 11704 18028 11756 18037
rect 17408 18028 17460 18080
rect 17684 18071 17736 18080
rect 17684 18037 17693 18071
rect 17693 18037 17727 18071
rect 17727 18037 17736 18071
rect 17684 18028 17736 18037
rect 18420 18028 18472 18080
rect 18604 18028 18656 18080
rect 25780 18300 25832 18352
rect 27344 18300 27396 18352
rect 27896 18300 27948 18352
rect 20996 18232 21048 18284
rect 23756 18275 23808 18284
rect 21732 18164 21784 18216
rect 23756 18241 23765 18275
rect 23765 18241 23799 18275
rect 23799 18241 23808 18275
rect 23756 18232 23808 18241
rect 23940 18275 23992 18284
rect 23940 18241 23949 18275
rect 23949 18241 23983 18275
rect 23983 18241 23992 18275
rect 23940 18232 23992 18241
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 24676 18232 24728 18284
rect 25688 18232 25740 18284
rect 26332 18232 26384 18284
rect 27068 18232 27120 18284
rect 35992 18300 36044 18352
rect 37188 18300 37240 18352
rect 29736 18164 29788 18216
rect 31208 18232 31260 18284
rect 33508 18232 33560 18284
rect 35900 18232 35952 18284
rect 36452 18275 36504 18284
rect 36452 18241 36461 18275
rect 36461 18241 36495 18275
rect 36495 18241 36504 18275
rect 36452 18232 36504 18241
rect 38016 18368 38068 18420
rect 39764 18300 39816 18352
rect 39856 18275 39908 18284
rect 31668 18164 31720 18216
rect 21180 18071 21232 18080
rect 21180 18037 21189 18071
rect 21189 18037 21223 18071
rect 21223 18037 21232 18071
rect 21180 18028 21232 18037
rect 24584 18028 24636 18080
rect 37096 18096 37148 18148
rect 39856 18241 39874 18275
rect 39874 18241 39908 18275
rect 39856 18232 39908 18241
rect 40040 18232 40092 18284
rect 37556 18139 37608 18148
rect 37556 18105 37565 18139
rect 37565 18105 37599 18139
rect 37599 18105 37608 18139
rect 37556 18096 37608 18105
rect 26976 18028 27028 18080
rect 29644 18071 29696 18080
rect 29644 18037 29653 18071
rect 29653 18037 29687 18071
rect 29687 18037 29696 18071
rect 29644 18028 29696 18037
rect 33508 18071 33560 18080
rect 33508 18037 33517 18071
rect 33517 18037 33551 18071
rect 33551 18037 33560 18071
rect 39028 18096 39080 18148
rect 38752 18071 38804 18080
rect 33508 18028 33560 18037
rect 38752 18037 38761 18071
rect 38761 18037 38795 18071
rect 38795 18037 38804 18071
rect 40592 18071 40644 18080
rect 38752 18028 38804 18037
rect 40592 18037 40601 18071
rect 40601 18037 40635 18071
rect 40635 18037 40644 18071
rect 40592 18028 40644 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 1768 17824 1820 17876
rect 4620 17867 4672 17876
rect 4620 17833 4629 17867
rect 4629 17833 4663 17867
rect 4663 17833 4672 17867
rect 4620 17824 4672 17833
rect 9220 17867 9272 17876
rect 9220 17833 9229 17867
rect 9229 17833 9263 17867
rect 9263 17833 9272 17867
rect 9220 17824 9272 17833
rect 11428 17824 11480 17876
rect 20076 17824 20128 17876
rect 21180 17824 21232 17876
rect 25688 17867 25740 17876
rect 25688 17833 25697 17867
rect 25697 17833 25731 17867
rect 25731 17833 25740 17867
rect 25688 17824 25740 17833
rect 27068 17824 27120 17876
rect 30288 17867 30340 17876
rect 30288 17833 30297 17867
rect 30297 17833 30331 17867
rect 30331 17833 30340 17867
rect 30288 17824 30340 17833
rect 30472 17867 30524 17876
rect 30472 17833 30481 17867
rect 30481 17833 30515 17867
rect 30515 17833 30524 17867
rect 30472 17824 30524 17833
rect 2872 17688 2924 17740
rect 2596 17663 2648 17672
rect 2596 17629 2605 17663
rect 2605 17629 2639 17663
rect 2639 17629 2648 17663
rect 2596 17620 2648 17629
rect 3792 17688 3844 17740
rect 9588 17688 9640 17740
rect 10232 17688 10284 17740
rect 13544 17731 13596 17740
rect 3884 17620 3936 17672
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 5908 17620 5960 17672
rect 9312 17663 9364 17672
rect 9312 17629 9321 17663
rect 9321 17629 9355 17663
rect 9355 17629 9364 17663
rect 9312 17620 9364 17629
rect 9404 17663 9456 17672
rect 9404 17629 9413 17663
rect 9413 17629 9447 17663
rect 9447 17629 9456 17663
rect 9404 17620 9456 17629
rect 10508 17620 10560 17672
rect 13544 17697 13553 17731
rect 13553 17697 13587 17731
rect 13587 17697 13596 17731
rect 13544 17688 13596 17697
rect 17500 17620 17552 17672
rect 18052 17688 18104 17740
rect 19984 17688 20036 17740
rect 17960 17620 18012 17672
rect 18236 17663 18288 17672
rect 18236 17629 18245 17663
rect 18245 17629 18279 17663
rect 18279 17629 18288 17663
rect 18236 17620 18288 17629
rect 18512 17620 18564 17672
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 22468 17756 22520 17808
rect 24216 17756 24268 17808
rect 28724 17756 28776 17808
rect 31116 17756 31168 17808
rect 27620 17688 27672 17740
rect 35348 17824 35400 17876
rect 38752 17824 38804 17876
rect 39856 17867 39908 17876
rect 39856 17833 39865 17867
rect 39865 17833 39899 17867
rect 39899 17833 39908 17867
rect 39856 17824 39908 17833
rect 36820 17756 36872 17808
rect 5172 17484 5224 17536
rect 6184 17484 6236 17536
rect 6644 17484 6696 17536
rect 7288 17552 7340 17604
rect 10048 17552 10100 17604
rect 11336 17552 11388 17604
rect 11704 17552 11756 17604
rect 12256 17552 12308 17604
rect 12716 17552 12768 17604
rect 7656 17484 7708 17536
rect 7748 17484 7800 17536
rect 10232 17484 10284 17536
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 17040 17484 17092 17536
rect 17776 17484 17828 17536
rect 18512 17484 18564 17536
rect 21088 17620 21140 17672
rect 23664 17620 23716 17672
rect 24400 17663 24452 17672
rect 24400 17629 24409 17663
rect 24409 17629 24443 17663
rect 24443 17629 24452 17663
rect 24400 17620 24452 17629
rect 24676 17663 24728 17672
rect 24676 17629 24685 17663
rect 24685 17629 24719 17663
rect 24719 17629 24728 17663
rect 24676 17620 24728 17629
rect 25872 17620 25924 17672
rect 22100 17527 22152 17536
rect 22100 17493 22109 17527
rect 22109 17493 22143 17527
rect 22143 17493 22152 17527
rect 22100 17484 22152 17493
rect 25780 17484 25832 17536
rect 26240 17620 26292 17672
rect 26516 17620 26568 17672
rect 26884 17620 26936 17672
rect 27252 17620 27304 17672
rect 27436 17620 27488 17672
rect 30564 17663 30616 17672
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30748 17663 30800 17672
rect 30564 17620 30616 17629
rect 30748 17629 30757 17663
rect 30757 17629 30791 17663
rect 30791 17629 30800 17663
rect 30748 17620 30800 17629
rect 27988 17552 28040 17604
rect 34980 17552 35032 17604
rect 27344 17484 27396 17536
rect 29920 17484 29972 17536
rect 35348 17620 35400 17672
rect 37924 17688 37976 17740
rect 36084 17663 36136 17672
rect 35256 17595 35308 17604
rect 35256 17561 35265 17595
rect 35265 17561 35299 17595
rect 35299 17561 35308 17595
rect 35256 17552 35308 17561
rect 36084 17629 36093 17663
rect 36093 17629 36127 17663
rect 36127 17629 36136 17663
rect 36084 17620 36136 17629
rect 36360 17620 36412 17672
rect 36176 17595 36228 17604
rect 36176 17561 36185 17595
rect 36185 17561 36219 17595
rect 36219 17561 36228 17595
rect 36176 17552 36228 17561
rect 36268 17595 36320 17604
rect 36268 17561 36277 17595
rect 36277 17561 36311 17595
rect 36311 17561 36320 17595
rect 36268 17552 36320 17561
rect 35900 17527 35952 17536
rect 35900 17493 35909 17527
rect 35909 17493 35943 17527
rect 35943 17493 35952 17527
rect 35900 17484 35952 17493
rect 36084 17484 36136 17536
rect 37280 17663 37332 17672
rect 37280 17629 37289 17663
rect 37289 17629 37323 17663
rect 37323 17629 37332 17663
rect 37280 17620 37332 17629
rect 37464 17663 37516 17672
rect 37464 17629 37473 17663
rect 37473 17629 37507 17663
rect 37507 17629 37516 17663
rect 37464 17620 37516 17629
rect 38844 17620 38896 17672
rect 40500 17663 40552 17672
rect 40500 17629 40509 17663
rect 40509 17629 40543 17663
rect 40543 17629 40552 17663
rect 40500 17620 40552 17629
rect 38568 17595 38620 17604
rect 36912 17527 36964 17536
rect 36912 17493 36921 17527
rect 36921 17493 36955 17527
rect 36955 17493 36964 17527
rect 36912 17484 36964 17493
rect 38568 17561 38577 17595
rect 38577 17561 38611 17595
rect 38611 17561 38620 17595
rect 38568 17552 38620 17561
rect 37832 17484 37884 17536
rect 39212 17484 39264 17536
rect 40592 17552 40644 17604
rect 40684 17484 40736 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4896 17280 4948 17332
rect 5264 17280 5316 17332
rect 7288 17280 7340 17332
rect 9312 17323 9364 17332
rect 9312 17289 9321 17323
rect 9321 17289 9355 17323
rect 9355 17289 9364 17323
rect 9312 17280 9364 17289
rect 9404 17280 9456 17332
rect 10692 17212 10744 17264
rect 11888 17212 11940 17264
rect 19984 17280 20036 17332
rect 20168 17280 20220 17332
rect 24216 17280 24268 17332
rect 13268 17255 13320 17264
rect 4620 17144 4672 17196
rect 4896 17144 4948 17196
rect 5264 17144 5316 17196
rect 6644 17144 6696 17196
rect 7748 17187 7800 17196
rect 7748 17153 7757 17187
rect 7757 17153 7791 17187
rect 7791 17153 7800 17187
rect 7748 17144 7800 17153
rect 7932 17187 7984 17196
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 9772 17144 9824 17196
rect 10048 17187 10100 17196
rect 10048 17153 10055 17187
rect 10055 17153 10100 17187
rect 10048 17144 10100 17153
rect 4712 17076 4764 17128
rect 7104 17076 7156 17128
rect 7288 17076 7340 17128
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 4804 17008 4856 17060
rect 9680 17008 9732 17060
rect 11336 17144 11388 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 13268 17221 13277 17255
rect 13277 17221 13311 17255
rect 13311 17221 13320 17255
rect 13268 17212 13320 17221
rect 18420 17212 18472 17264
rect 18788 17212 18840 17264
rect 20812 17212 20864 17264
rect 11704 17144 11756 17153
rect 10416 17076 10468 17128
rect 11796 17076 11848 17128
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 13360 17187 13412 17196
rect 13360 17153 13405 17187
rect 13405 17153 13412 17187
rect 13360 17144 13412 17153
rect 14004 17144 14056 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 20996 17144 21048 17196
rect 21732 17144 21784 17196
rect 21916 17144 21968 17196
rect 22652 17187 22704 17196
rect 22652 17153 22661 17187
rect 22661 17153 22695 17187
rect 22695 17153 22704 17187
rect 22652 17144 22704 17153
rect 26608 17280 26660 17332
rect 27252 17280 27304 17332
rect 35256 17280 35308 17332
rect 36268 17280 36320 17332
rect 37188 17280 37240 17332
rect 39028 17323 39080 17332
rect 39028 17289 39037 17323
rect 39037 17289 39071 17323
rect 39071 17289 39080 17323
rect 39028 17280 39080 17289
rect 25320 17144 25372 17196
rect 35900 17144 35952 17196
rect 36728 17144 36780 17196
rect 38568 17144 38620 17196
rect 10784 17008 10836 17060
rect 19708 17076 19760 17128
rect 19248 17008 19300 17060
rect 6000 16940 6052 16992
rect 6644 16983 6696 16992
rect 6644 16949 6653 16983
rect 6653 16949 6687 16983
rect 6687 16949 6696 16983
rect 6644 16940 6696 16949
rect 9404 16940 9456 16992
rect 13636 16940 13688 16992
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 18236 16940 18288 16992
rect 18788 16940 18840 16992
rect 19524 16983 19576 16992
rect 19524 16949 19533 16983
rect 19533 16949 19567 16983
rect 19567 16949 19576 16983
rect 19524 16940 19576 16949
rect 19984 17051 20036 17060
rect 19984 17017 19993 17051
rect 19993 17017 20027 17051
rect 20027 17017 20036 17051
rect 19984 17008 20036 17017
rect 21916 17008 21968 17060
rect 24400 17076 24452 17128
rect 24124 17008 24176 17060
rect 25228 17076 25280 17128
rect 25872 17076 25924 17128
rect 33784 17119 33836 17128
rect 27160 17008 27212 17060
rect 29552 17008 29604 17060
rect 33784 17085 33793 17119
rect 33793 17085 33827 17119
rect 33827 17085 33836 17119
rect 33784 17076 33836 17085
rect 34612 17076 34664 17128
rect 34980 17076 35032 17128
rect 36084 17076 36136 17128
rect 36820 17076 36872 17128
rect 38200 17076 38252 17128
rect 40500 17076 40552 17128
rect 58164 17051 58216 17060
rect 58164 17017 58173 17051
rect 58173 17017 58207 17051
rect 58207 17017 58216 17051
rect 58164 17008 58216 17017
rect 24768 16940 24820 16992
rect 24952 16983 25004 16992
rect 24952 16949 24961 16983
rect 24961 16949 24995 16983
rect 24995 16949 25004 16983
rect 24952 16940 25004 16949
rect 32864 16940 32916 16992
rect 35532 16940 35584 16992
rect 37740 16940 37792 16992
rect 39764 16940 39816 16992
rect 40040 16940 40092 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 5264 16779 5316 16788
rect 5264 16745 5273 16779
rect 5273 16745 5307 16779
rect 5307 16745 5316 16779
rect 5264 16736 5316 16745
rect 9680 16736 9732 16788
rect 12716 16779 12768 16788
rect 8300 16668 8352 16720
rect 12716 16745 12725 16779
rect 12725 16745 12759 16779
rect 12759 16745 12768 16779
rect 12716 16736 12768 16745
rect 13452 16736 13504 16788
rect 17316 16736 17368 16788
rect 17500 16779 17552 16788
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 18696 16736 18748 16788
rect 19432 16736 19484 16788
rect 19708 16779 19760 16788
rect 19708 16745 19717 16779
rect 19717 16745 19751 16779
rect 19751 16745 19760 16779
rect 19708 16736 19760 16745
rect 20076 16736 20128 16788
rect 21916 16779 21968 16788
rect 21916 16745 21925 16779
rect 21925 16745 21959 16779
rect 21959 16745 21968 16779
rect 21916 16736 21968 16745
rect 24584 16779 24636 16788
rect 14096 16668 14148 16720
rect 24584 16745 24593 16779
rect 24593 16745 24627 16779
rect 24627 16745 24636 16779
rect 24584 16736 24636 16745
rect 25320 16779 25372 16788
rect 25320 16745 25329 16779
rect 25329 16745 25363 16779
rect 25363 16745 25372 16779
rect 25320 16736 25372 16745
rect 26240 16736 26292 16788
rect 27436 16736 27488 16788
rect 27712 16736 27764 16788
rect 34060 16736 34112 16788
rect 35900 16779 35952 16788
rect 35900 16745 35909 16779
rect 35909 16745 35943 16779
rect 35943 16745 35952 16779
rect 35900 16736 35952 16745
rect 36360 16736 36412 16788
rect 27804 16711 27856 16720
rect 5356 16532 5408 16584
rect 9956 16575 10008 16584
rect 9956 16541 9965 16575
rect 9965 16541 9999 16575
rect 9999 16541 10008 16575
rect 9956 16532 10008 16541
rect 10140 16575 10192 16584
rect 10140 16541 10147 16575
rect 10147 16541 10192 16575
rect 10140 16532 10192 16541
rect 10784 16600 10836 16652
rect 15292 16643 15344 16652
rect 10416 16575 10468 16584
rect 10416 16541 10430 16575
rect 10430 16541 10464 16575
rect 10464 16541 10468 16575
rect 11244 16575 11296 16584
rect 10416 16532 10468 16541
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 10324 16507 10376 16516
rect 10324 16473 10333 16507
rect 10333 16473 10367 16507
rect 10367 16473 10376 16507
rect 10324 16464 10376 16473
rect 10968 16464 11020 16516
rect 11796 16532 11848 16584
rect 12164 16532 12216 16584
rect 15292 16609 15301 16643
rect 15301 16609 15335 16643
rect 15335 16609 15344 16643
rect 15292 16600 15344 16609
rect 15936 16600 15988 16652
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 3884 16396 3936 16448
rect 10600 16439 10652 16448
rect 10600 16405 10609 16439
rect 10609 16405 10643 16439
rect 10643 16405 10652 16439
rect 10600 16396 10652 16405
rect 10784 16396 10836 16448
rect 11612 16507 11664 16516
rect 11612 16473 11621 16507
rect 11621 16473 11655 16507
rect 11655 16473 11664 16507
rect 11612 16464 11664 16473
rect 11888 16464 11940 16516
rect 13636 16532 13688 16584
rect 15200 16532 15252 16584
rect 17500 16532 17552 16584
rect 23204 16643 23256 16652
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 14556 16507 14608 16516
rect 14556 16473 14565 16507
rect 14565 16473 14599 16507
rect 14599 16473 14608 16507
rect 14556 16464 14608 16473
rect 12716 16396 12768 16448
rect 13728 16396 13780 16448
rect 19524 16532 19576 16584
rect 20076 16532 20128 16584
rect 20168 16532 20220 16584
rect 23204 16609 23213 16643
rect 23213 16609 23247 16643
rect 23247 16609 23256 16643
rect 23204 16600 23256 16609
rect 22652 16575 22704 16584
rect 19524 16396 19576 16448
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 24492 16600 24544 16652
rect 24768 16600 24820 16652
rect 27804 16677 27813 16711
rect 27813 16677 27847 16711
rect 27847 16677 27856 16711
rect 27804 16668 27856 16677
rect 29552 16643 29604 16652
rect 22652 16532 22704 16541
rect 24676 16575 24728 16584
rect 24676 16541 24685 16575
rect 24685 16541 24719 16575
rect 24719 16541 24728 16575
rect 24676 16532 24728 16541
rect 25044 16532 25096 16584
rect 26608 16532 26660 16584
rect 29552 16609 29561 16643
rect 29561 16609 29595 16643
rect 29595 16609 29604 16643
rect 29552 16600 29604 16609
rect 29920 16600 29972 16652
rect 27712 16532 27764 16584
rect 32588 16600 32640 16652
rect 32864 16643 32916 16652
rect 32864 16609 32873 16643
rect 32873 16609 32907 16643
rect 32907 16609 32916 16643
rect 32864 16600 32916 16609
rect 33784 16668 33836 16720
rect 20628 16464 20680 16516
rect 34704 16600 34756 16652
rect 37924 16711 37976 16720
rect 37924 16677 37933 16711
rect 37933 16677 37967 16711
rect 37967 16677 37976 16711
rect 37924 16668 37976 16677
rect 40040 16600 40092 16652
rect 34980 16575 35032 16584
rect 34980 16541 34989 16575
rect 34989 16541 35023 16575
rect 35023 16541 35032 16575
rect 34980 16532 35032 16541
rect 35532 16532 35584 16584
rect 20812 16396 20864 16448
rect 20996 16396 21048 16448
rect 24308 16396 24360 16448
rect 34704 16396 34756 16448
rect 38660 16464 38712 16516
rect 37096 16396 37148 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 5448 16235 5500 16244
rect 5448 16201 5457 16235
rect 5457 16201 5491 16235
rect 5491 16201 5500 16235
rect 5448 16192 5500 16201
rect 6920 16192 6972 16244
rect 10876 16192 10928 16244
rect 11980 16192 12032 16244
rect 15384 16192 15436 16244
rect 10324 16124 10376 16176
rect 11796 16124 11848 16176
rect 2504 16056 2556 16108
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 9404 16056 9456 16108
rect 10048 16056 10100 16108
rect 10232 16056 10284 16108
rect 11336 16056 11388 16108
rect 3976 15988 4028 16040
rect 11060 15988 11112 16040
rect 12440 16056 12492 16108
rect 4988 15920 5040 15972
rect 2228 15895 2280 15904
rect 2228 15861 2237 15895
rect 2237 15861 2271 15895
rect 2271 15861 2280 15895
rect 2228 15852 2280 15861
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 6644 15852 6696 15904
rect 10048 15852 10100 15904
rect 11704 15852 11756 15904
rect 12164 15988 12216 16040
rect 12716 16056 12768 16108
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 14556 16056 14608 16108
rect 13728 15988 13780 16040
rect 14188 15920 14240 15972
rect 14832 16099 14884 16108
rect 14832 16065 14841 16099
rect 14841 16065 14875 16099
rect 14875 16065 14884 16099
rect 14832 16056 14884 16065
rect 16764 16124 16816 16176
rect 15936 16056 15988 16108
rect 16672 15988 16724 16040
rect 17224 16192 17276 16244
rect 20628 16192 20680 16244
rect 20812 16235 20864 16244
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 21732 16192 21784 16244
rect 22652 16192 22704 16244
rect 24492 16192 24544 16244
rect 34980 16192 35032 16244
rect 36912 16192 36964 16244
rect 37740 16192 37792 16244
rect 17316 16099 17368 16108
rect 17316 16065 17325 16099
rect 17325 16065 17359 16099
rect 17359 16065 17368 16099
rect 17316 16056 17368 16065
rect 17776 16056 17828 16108
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 19432 16099 19484 16108
rect 19432 16065 19441 16099
rect 19441 16065 19475 16099
rect 19475 16065 19484 16099
rect 19432 16056 19484 16065
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 27896 16056 27948 16108
rect 30748 16056 30800 16108
rect 32036 16056 32088 16108
rect 35900 16124 35952 16176
rect 36360 16124 36412 16176
rect 36544 16124 36596 16176
rect 38844 16192 38896 16244
rect 39028 16192 39080 16244
rect 19340 15988 19392 16040
rect 25044 16031 25096 16040
rect 25044 15997 25053 16031
rect 25053 15997 25087 16031
rect 25087 15997 25096 16031
rect 25044 15988 25096 15997
rect 27436 15988 27488 16040
rect 30380 15988 30432 16040
rect 15384 15920 15436 15972
rect 20536 15920 20588 15972
rect 31852 15920 31904 15972
rect 32588 16056 32640 16108
rect 34612 16099 34664 16108
rect 34612 16065 34621 16099
rect 34621 16065 34655 16099
rect 34655 16065 34664 16099
rect 34612 16056 34664 16065
rect 36820 16056 36872 16108
rect 37188 16056 37240 16108
rect 34520 15988 34572 16040
rect 14372 15895 14424 15904
rect 14372 15861 14381 15895
rect 14381 15861 14415 15895
rect 14415 15861 14424 15895
rect 14372 15852 14424 15861
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 18052 15852 18104 15904
rect 20260 15852 20312 15904
rect 20720 15852 20772 15904
rect 24952 15852 25004 15904
rect 25688 15852 25740 15904
rect 33232 15852 33284 15904
rect 36636 15852 36688 15904
rect 36912 15852 36964 15904
rect 38660 16031 38712 16040
rect 38660 15997 38669 16031
rect 38669 15997 38703 16031
rect 38703 15997 38712 16031
rect 38660 15988 38712 15997
rect 37556 15852 37608 15904
rect 39212 16056 39264 16108
rect 58164 15895 58216 15904
rect 58164 15861 58173 15895
rect 58173 15861 58207 15895
rect 58207 15861 58216 15895
rect 58164 15852 58216 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 3976 15648 4028 15700
rect 5264 15648 5316 15700
rect 7196 15691 7248 15700
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 7380 15648 7432 15700
rect 11244 15648 11296 15700
rect 12072 15648 12124 15700
rect 23204 15691 23256 15700
rect 7932 15580 7984 15632
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 23296 15648 23348 15700
rect 24860 15648 24912 15700
rect 25596 15648 25648 15700
rect 25964 15648 26016 15700
rect 27896 15648 27948 15700
rect 29276 15648 29328 15700
rect 34060 15691 34112 15700
rect 2136 15487 2188 15496
rect 2136 15453 2145 15487
rect 2145 15453 2179 15487
rect 2179 15453 2188 15487
rect 2136 15444 2188 15453
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 3424 15444 3476 15496
rect 8208 15512 8260 15564
rect 4160 15444 4212 15496
rect 5908 15444 5960 15496
rect 8300 15444 8352 15496
rect 23020 15580 23072 15632
rect 10876 15512 10928 15564
rect 13544 15512 13596 15564
rect 19248 15512 19300 15564
rect 24768 15580 24820 15632
rect 34060 15657 34069 15691
rect 34069 15657 34103 15691
rect 34103 15657 34112 15691
rect 34060 15648 34112 15657
rect 23572 15555 23624 15564
rect 23572 15521 23581 15555
rect 23581 15521 23615 15555
rect 23615 15521 23624 15555
rect 23572 15512 23624 15521
rect 5356 15376 5408 15428
rect 9404 15444 9456 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 14372 15487 14424 15496
rect 14372 15453 14406 15487
rect 14406 15453 14424 15487
rect 14372 15444 14424 15453
rect 17868 15444 17920 15496
rect 20260 15444 20312 15496
rect 20444 15487 20496 15496
rect 20444 15453 20453 15487
rect 20453 15453 20487 15487
rect 20487 15453 20496 15487
rect 20444 15444 20496 15453
rect 20536 15444 20588 15496
rect 22652 15444 22704 15496
rect 23664 15487 23716 15496
rect 11520 15376 11572 15428
rect 16120 15376 16172 15428
rect 23664 15453 23673 15487
rect 23673 15453 23707 15487
rect 23707 15453 23716 15487
rect 23664 15444 23716 15453
rect 26608 15487 26660 15496
rect 26608 15453 26617 15487
rect 26617 15453 26651 15487
rect 26651 15453 26660 15487
rect 26608 15444 26660 15453
rect 29828 15444 29880 15496
rect 24952 15376 25004 15428
rect 25688 15376 25740 15428
rect 28724 15376 28776 15428
rect 3516 15308 3568 15360
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 5816 15351 5868 15360
rect 5816 15317 5825 15351
rect 5825 15317 5859 15351
rect 5859 15317 5868 15351
rect 5816 15308 5868 15317
rect 7012 15351 7064 15360
rect 7012 15317 7021 15351
rect 7021 15317 7055 15351
rect 7055 15317 7064 15351
rect 7012 15308 7064 15317
rect 9956 15308 10008 15360
rect 11888 15308 11940 15360
rect 15292 15308 15344 15360
rect 18144 15308 18196 15360
rect 20076 15308 20128 15360
rect 20352 15308 20404 15360
rect 27988 15308 28040 15360
rect 30380 15487 30432 15496
rect 30380 15453 30389 15487
rect 30389 15453 30423 15487
rect 30423 15453 30432 15487
rect 30380 15444 30432 15453
rect 30472 15444 30524 15496
rect 31852 15512 31904 15564
rect 32772 15444 32824 15496
rect 34060 15444 34112 15496
rect 34796 15444 34848 15496
rect 36820 15487 36872 15496
rect 34612 15376 34664 15428
rect 36820 15453 36829 15487
rect 36829 15453 36863 15487
rect 36863 15453 36872 15487
rect 36820 15444 36872 15453
rect 37188 15444 37240 15496
rect 37832 15487 37884 15496
rect 37832 15453 37841 15487
rect 37841 15453 37875 15487
rect 37875 15453 37884 15487
rect 37832 15444 37884 15453
rect 37280 15376 37332 15428
rect 37464 15376 37516 15428
rect 31300 15308 31352 15360
rect 37096 15308 37148 15360
rect 37556 15308 37608 15360
rect 38384 15308 38436 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 2964 15147 3016 15156
rect 2964 15113 2973 15147
rect 2973 15113 3007 15147
rect 3007 15113 3016 15147
rect 2964 15104 3016 15113
rect 4160 15104 4212 15156
rect 14188 15147 14240 15156
rect 14188 15113 14197 15147
rect 14197 15113 14231 15147
rect 14231 15113 14240 15147
rect 14188 15104 14240 15113
rect 14832 15104 14884 15156
rect 16672 15147 16724 15156
rect 16672 15113 16681 15147
rect 16681 15113 16715 15147
rect 16715 15113 16724 15147
rect 16672 15104 16724 15113
rect 2780 15036 2832 15088
rect 2228 14968 2280 15020
rect 4620 15036 4672 15088
rect 18144 15104 18196 15156
rect 3516 14968 3568 15020
rect 20812 15036 20864 15088
rect 21088 15104 21140 15156
rect 22008 15104 22060 15156
rect 23204 15104 23256 15156
rect 29828 15147 29880 15156
rect 6920 14968 6972 15020
rect 15292 15011 15344 15020
rect 15292 14977 15301 15011
rect 15301 14977 15335 15011
rect 15335 14977 15344 15011
rect 15292 14968 15344 14977
rect 17776 14968 17828 15020
rect 17868 14968 17920 15020
rect 18052 14968 18104 15020
rect 19340 14875 19392 14884
rect 19340 14841 19349 14875
rect 19349 14841 19383 14875
rect 19383 14841 19392 14875
rect 20536 14968 20588 15020
rect 21456 14900 21508 14952
rect 22100 14900 22152 14952
rect 19340 14832 19392 14841
rect 4804 14807 4856 14816
rect 4804 14773 4813 14807
rect 4813 14773 4847 14807
rect 4847 14773 4856 14807
rect 4804 14764 4856 14773
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 12808 14764 12860 14816
rect 20444 14764 20496 14816
rect 20536 14764 20588 14816
rect 22928 15036 22980 15088
rect 25136 15036 25188 15088
rect 29828 15113 29837 15147
rect 29837 15113 29871 15147
rect 29871 15113 29880 15147
rect 29828 15104 29880 15113
rect 30472 15104 30524 15156
rect 34060 15147 34112 15156
rect 34060 15113 34069 15147
rect 34069 15113 34103 15147
rect 34103 15113 34112 15147
rect 34060 15104 34112 15113
rect 35900 15104 35952 15156
rect 37188 15104 37240 15156
rect 37280 15104 37332 15156
rect 30748 15036 30800 15088
rect 32772 15036 32824 15088
rect 22652 15011 22704 15020
rect 22652 14977 22661 15011
rect 22661 14977 22695 15011
rect 22695 14977 22704 15011
rect 22652 14968 22704 14977
rect 23388 14968 23440 15020
rect 23664 15011 23716 15020
rect 23664 14977 23673 15011
rect 23673 14977 23707 15011
rect 23707 14977 23716 15011
rect 23664 14968 23716 14977
rect 23204 14832 23256 14884
rect 24584 14943 24636 14952
rect 24584 14909 24593 14943
rect 24593 14909 24627 14943
rect 24627 14909 24636 14943
rect 24584 14900 24636 14909
rect 24860 14968 24912 15020
rect 25688 14968 25740 15020
rect 28540 14968 28592 15020
rect 31300 14968 31352 15020
rect 33232 15011 33284 15020
rect 33232 14977 33250 15011
rect 33250 14977 33284 15011
rect 33232 14968 33284 14977
rect 34520 14968 34572 15020
rect 25320 14900 25372 14952
rect 28448 14943 28500 14952
rect 28448 14909 28457 14943
rect 28457 14909 28491 14943
rect 28491 14909 28500 14943
rect 28448 14900 28500 14909
rect 34060 14900 34112 14952
rect 34704 14900 34756 14952
rect 26608 14832 26660 14884
rect 37556 14968 37608 15020
rect 37096 14900 37148 14952
rect 38568 14968 38620 15020
rect 40040 15011 40092 15020
rect 40040 14977 40049 15011
rect 40049 14977 40083 15011
rect 40083 14977 40092 15011
rect 40040 14968 40092 14977
rect 39028 14832 39080 14884
rect 22652 14764 22704 14816
rect 23664 14764 23716 14816
rect 23848 14807 23900 14816
rect 23848 14773 23857 14807
rect 23857 14773 23891 14807
rect 23891 14773 23900 14807
rect 23848 14764 23900 14773
rect 24492 14807 24544 14816
rect 24492 14773 24501 14807
rect 24501 14773 24535 14807
rect 24535 14773 24544 14807
rect 24492 14764 24544 14773
rect 26332 14764 26384 14816
rect 27160 14764 27212 14816
rect 27436 14764 27488 14816
rect 28356 14764 28408 14816
rect 32036 14764 32088 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2320 14560 2372 14612
rect 3056 14560 3108 14612
rect 6920 14603 6972 14612
rect 6920 14569 6929 14603
rect 6929 14569 6963 14603
rect 6963 14569 6972 14603
rect 6920 14560 6972 14569
rect 2136 14492 2188 14544
rect 3884 14492 3936 14544
rect 2964 14467 3016 14476
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 3608 14424 3660 14476
rect 4068 14424 4120 14476
rect 6276 14492 6328 14544
rect 13176 14560 13228 14612
rect 17316 14560 17368 14612
rect 19340 14560 19392 14612
rect 19984 14560 20036 14612
rect 20812 14560 20864 14612
rect 23848 14560 23900 14612
rect 4804 14424 4856 14476
rect 5816 14424 5868 14476
rect 7196 14424 7248 14476
rect 13544 14424 13596 14476
rect 3424 14356 3476 14408
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 5908 14356 5960 14408
rect 6276 14356 6328 14408
rect 5172 14288 5224 14340
rect 6092 14288 6144 14340
rect 7104 14356 7156 14408
rect 7748 14356 7800 14408
rect 8208 14356 8260 14408
rect 10232 14356 10284 14408
rect 10876 14356 10928 14408
rect 21732 14492 21784 14544
rect 7012 14288 7064 14340
rect 10140 14288 10192 14340
rect 11520 14331 11572 14340
rect 11520 14297 11529 14331
rect 11529 14297 11563 14331
rect 11563 14297 11572 14331
rect 11520 14288 11572 14297
rect 7288 14220 7340 14272
rect 9588 14263 9640 14272
rect 9588 14229 9597 14263
rect 9597 14229 9631 14263
rect 9631 14229 9640 14263
rect 9588 14220 9640 14229
rect 20352 14356 20404 14408
rect 20536 14399 20588 14408
rect 20536 14365 20545 14399
rect 20545 14365 20579 14399
rect 20579 14365 20588 14399
rect 20536 14356 20588 14365
rect 21088 14356 21140 14408
rect 15292 14288 15344 14340
rect 21732 14288 21784 14340
rect 22008 14288 22060 14340
rect 23388 14492 23440 14544
rect 24492 14492 24544 14544
rect 27804 14560 27856 14612
rect 28540 14603 28592 14612
rect 28540 14569 28549 14603
rect 28549 14569 28583 14603
rect 28583 14569 28592 14603
rect 28540 14560 28592 14569
rect 34612 14560 34664 14612
rect 23664 14356 23716 14408
rect 23296 14331 23348 14340
rect 23296 14297 23305 14331
rect 23305 14297 23339 14331
rect 23339 14297 23348 14331
rect 23296 14288 23348 14297
rect 24492 14220 24544 14272
rect 25964 14356 26016 14408
rect 28080 14492 28132 14544
rect 32312 14492 32364 14544
rect 27988 14356 28040 14408
rect 25688 14288 25740 14340
rect 26056 14331 26108 14340
rect 26056 14297 26065 14331
rect 26065 14297 26099 14331
rect 26099 14297 26108 14331
rect 26056 14288 26108 14297
rect 27436 14288 27488 14340
rect 28264 14399 28316 14408
rect 28264 14365 28273 14399
rect 28273 14365 28307 14399
rect 28307 14365 28316 14399
rect 28264 14356 28316 14365
rect 29460 14356 29512 14408
rect 30288 14356 30340 14408
rect 34520 14356 34572 14408
rect 36820 14424 36872 14476
rect 40224 14424 40276 14476
rect 36268 14399 36320 14408
rect 36268 14365 36277 14399
rect 36277 14365 36311 14399
rect 36311 14365 36320 14399
rect 36268 14356 36320 14365
rect 37096 14356 37148 14408
rect 38200 14356 38252 14408
rect 28356 14288 28408 14340
rect 28724 14288 28776 14340
rect 38292 14288 38344 14340
rect 40684 14356 40736 14408
rect 58164 14399 58216 14408
rect 58164 14365 58173 14399
rect 58173 14365 58207 14399
rect 58207 14365 58216 14399
rect 58164 14356 58216 14365
rect 25320 14263 25372 14272
rect 25320 14229 25329 14263
rect 25329 14229 25363 14263
rect 25363 14229 25372 14263
rect 25320 14220 25372 14229
rect 25964 14220 26016 14272
rect 28264 14220 28316 14272
rect 29920 14263 29972 14272
rect 29920 14229 29929 14263
rect 29929 14229 29963 14263
rect 29963 14229 29972 14263
rect 29920 14220 29972 14229
rect 35440 14220 35492 14272
rect 37096 14263 37148 14272
rect 37096 14229 37105 14263
rect 37105 14229 37139 14263
rect 37139 14229 37148 14263
rect 37096 14220 37148 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 3976 14016 4028 14068
rect 10140 14059 10192 14068
rect 10140 14025 10149 14059
rect 10149 14025 10183 14059
rect 10183 14025 10192 14059
rect 10140 14016 10192 14025
rect 10232 14016 10284 14068
rect 23204 14016 23256 14068
rect 23296 14016 23348 14068
rect 26056 14016 26108 14068
rect 4804 13948 4856 14000
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 14280 13948 14332 14000
rect 16672 13948 16724 14000
rect 19248 13948 19300 14000
rect 21088 13991 21140 14000
rect 21088 13957 21097 13991
rect 21097 13957 21131 13991
rect 21131 13957 21140 13991
rect 21088 13948 21140 13957
rect 25228 13948 25280 14000
rect 9864 13880 9916 13932
rect 14004 13880 14056 13932
rect 17316 13880 17368 13932
rect 25596 13880 25648 13932
rect 25964 13880 26016 13932
rect 27160 13948 27212 14000
rect 26332 13880 26384 13932
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 34704 14016 34756 14068
rect 27620 13948 27672 14000
rect 29552 13948 29604 14000
rect 32312 13948 32364 14000
rect 26424 13880 26476 13889
rect 29276 13880 29328 13932
rect 30288 13880 30340 13932
rect 6460 13855 6512 13864
rect 6460 13821 6469 13855
rect 6469 13821 6503 13855
rect 6503 13821 6512 13855
rect 6460 13812 6512 13821
rect 7288 13812 7340 13864
rect 9772 13855 9824 13864
rect 9772 13821 9781 13855
rect 9781 13821 9815 13855
rect 9815 13821 9824 13855
rect 9772 13812 9824 13821
rect 14096 13812 14148 13864
rect 17960 13812 18012 13864
rect 5816 13744 5868 13796
rect 11612 13744 11664 13796
rect 12072 13787 12124 13796
rect 12072 13753 12081 13787
rect 12081 13753 12115 13787
rect 12115 13753 12124 13787
rect 12072 13744 12124 13753
rect 14372 13676 14424 13728
rect 20168 13676 20220 13728
rect 25780 13719 25832 13728
rect 25780 13685 25789 13719
rect 25789 13685 25823 13719
rect 25823 13685 25832 13719
rect 25780 13676 25832 13685
rect 35900 14016 35952 14068
rect 37372 14016 37424 14068
rect 37740 14016 37792 14068
rect 37924 14016 37976 14068
rect 36176 13948 36228 14000
rect 33140 13812 33192 13864
rect 35808 13880 35860 13932
rect 40224 13948 40276 14000
rect 38844 13880 38896 13932
rect 40040 13880 40092 13932
rect 35348 13855 35400 13864
rect 35348 13821 35357 13855
rect 35357 13821 35391 13855
rect 35391 13821 35400 13855
rect 35348 13812 35400 13821
rect 35440 13812 35492 13864
rect 38292 13812 38344 13864
rect 26332 13676 26384 13728
rect 28448 13676 28500 13728
rect 28724 13719 28776 13728
rect 28724 13685 28733 13719
rect 28733 13685 28767 13719
rect 28767 13685 28776 13719
rect 28724 13676 28776 13685
rect 31116 13676 31168 13728
rect 36912 13676 36964 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10692 13472 10744 13524
rect 15476 13472 15528 13524
rect 17868 13515 17920 13524
rect 17868 13481 17877 13515
rect 17877 13481 17911 13515
rect 17911 13481 17920 13515
rect 17868 13472 17920 13481
rect 19248 13515 19300 13524
rect 19248 13481 19257 13515
rect 19257 13481 19291 13515
rect 19291 13481 19300 13515
rect 19248 13472 19300 13481
rect 22928 13472 22980 13524
rect 25596 13472 25648 13524
rect 29276 13472 29328 13524
rect 29552 13515 29604 13524
rect 29552 13481 29561 13515
rect 29561 13481 29595 13515
rect 29595 13481 29604 13515
rect 29552 13472 29604 13481
rect 30104 13472 30156 13524
rect 32128 13472 32180 13524
rect 36176 13472 36228 13524
rect 38844 13515 38896 13524
rect 38844 13481 38853 13515
rect 38853 13481 38887 13515
rect 38887 13481 38896 13515
rect 38844 13472 38896 13481
rect 12256 13404 12308 13456
rect 8576 13268 8628 13320
rect 12072 13268 12124 13320
rect 14924 13336 14976 13388
rect 10508 13200 10560 13252
rect 13268 13200 13320 13252
rect 13544 13243 13596 13252
rect 13544 13209 13553 13243
rect 13553 13209 13587 13243
rect 13587 13209 13596 13243
rect 13544 13200 13596 13209
rect 12348 13132 12400 13184
rect 14188 13175 14240 13184
rect 14188 13141 14197 13175
rect 14197 13141 14231 13175
rect 14231 13141 14240 13175
rect 14188 13132 14240 13141
rect 14669 13308 14721 13317
rect 14669 13274 14678 13308
rect 14678 13274 14712 13308
rect 14712 13274 14721 13308
rect 14669 13265 14721 13274
rect 15292 13268 15344 13320
rect 22468 13404 22520 13456
rect 24676 13404 24728 13456
rect 26240 13404 26292 13456
rect 21456 13379 21508 13388
rect 21456 13345 21465 13379
rect 21465 13345 21499 13379
rect 21499 13345 21508 13379
rect 21456 13336 21508 13345
rect 26424 13404 26476 13456
rect 28264 13404 28316 13456
rect 20260 13268 20312 13320
rect 20720 13268 20772 13320
rect 25780 13268 25832 13320
rect 14924 13200 14976 13252
rect 15200 13200 15252 13252
rect 25136 13243 25188 13252
rect 25136 13209 25145 13243
rect 25145 13209 25179 13243
rect 25179 13209 25188 13243
rect 25136 13200 25188 13209
rect 25688 13200 25740 13252
rect 25872 13200 25924 13252
rect 15384 13175 15436 13184
rect 15384 13141 15393 13175
rect 15393 13141 15427 13175
rect 15427 13141 15436 13175
rect 15384 13132 15436 13141
rect 20536 13175 20588 13184
rect 20536 13141 20545 13175
rect 20545 13141 20579 13175
rect 20579 13141 20588 13175
rect 20536 13132 20588 13141
rect 25780 13175 25832 13184
rect 25780 13141 25789 13175
rect 25789 13141 25823 13175
rect 25823 13141 25832 13175
rect 25780 13132 25832 13141
rect 26240 13311 26292 13320
rect 26240 13277 26254 13311
rect 26254 13277 26288 13311
rect 26288 13277 26292 13311
rect 26240 13268 26292 13277
rect 27252 13277 27261 13296
rect 27261 13277 27295 13296
rect 27295 13277 27304 13296
rect 27252 13244 27304 13277
rect 27160 13132 27212 13184
rect 27436 13308 27488 13320
rect 27436 13274 27445 13308
rect 27445 13274 27479 13308
rect 27479 13274 27488 13308
rect 28080 13311 28132 13320
rect 27436 13268 27488 13274
rect 28080 13277 28089 13311
rect 28089 13277 28123 13311
rect 28123 13277 28132 13311
rect 28080 13268 28132 13277
rect 29920 13336 29972 13388
rect 33140 13336 33192 13388
rect 39028 13404 39080 13456
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 28540 13268 28592 13320
rect 32772 13311 32824 13320
rect 32772 13277 32781 13311
rect 32781 13277 32815 13311
rect 32815 13277 32824 13311
rect 32772 13268 32824 13277
rect 34704 13311 34756 13320
rect 34704 13277 34713 13311
rect 34713 13277 34747 13311
rect 34747 13277 34756 13311
rect 34704 13268 34756 13277
rect 36544 13336 36596 13388
rect 37096 13336 37148 13388
rect 30104 13200 30156 13252
rect 33508 13200 33560 13252
rect 34428 13200 34480 13252
rect 34796 13200 34848 13252
rect 37648 13268 37700 13320
rect 37740 13311 37792 13320
rect 37740 13277 37749 13311
rect 37749 13277 37783 13311
rect 37783 13277 37792 13311
rect 38200 13311 38252 13320
rect 37740 13268 37792 13277
rect 38200 13277 38209 13311
rect 38209 13277 38243 13311
rect 38243 13277 38252 13311
rect 38200 13268 38252 13277
rect 38384 13311 38436 13320
rect 38384 13277 38393 13311
rect 38393 13277 38427 13311
rect 38427 13277 38436 13311
rect 38384 13268 38436 13277
rect 37096 13175 37148 13184
rect 37096 13141 37105 13175
rect 37105 13141 37139 13175
rect 37139 13141 37148 13175
rect 37096 13132 37148 13141
rect 38292 13200 38344 13252
rect 38568 13311 38620 13320
rect 38568 13277 38577 13311
rect 38577 13277 38611 13311
rect 38611 13277 38620 13311
rect 38568 13268 38620 13277
rect 40224 13268 40276 13320
rect 58164 13311 58216 13320
rect 58164 13277 58173 13311
rect 58173 13277 58207 13311
rect 58207 13277 58216 13311
rect 58164 13268 58216 13277
rect 39120 13132 39172 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4896 12928 4948 12980
rect 5264 12928 5316 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 13268 12928 13320 12980
rect 14188 12860 14240 12912
rect 15476 12903 15528 12912
rect 15476 12869 15485 12903
rect 15485 12869 15519 12903
rect 15519 12869 15528 12903
rect 15476 12860 15528 12869
rect 16672 12860 16724 12912
rect 17868 12860 17920 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 2320 12656 2372 12708
rect 7380 12792 7432 12844
rect 9128 12792 9180 12844
rect 14372 12792 14424 12844
rect 3424 12767 3476 12776
rect 3424 12733 3433 12767
rect 3433 12733 3467 12767
rect 3467 12733 3476 12767
rect 3424 12724 3476 12733
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 3884 12724 3936 12776
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8576 12767 8628 12776
rect 8116 12724 8168 12733
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 14096 12724 14148 12776
rect 14648 12841 14700 12844
rect 14648 12807 14657 12841
rect 14657 12807 14691 12841
rect 14691 12807 14700 12841
rect 14648 12792 14700 12807
rect 15292 12792 15344 12844
rect 17500 12792 17552 12844
rect 18052 12835 18104 12844
rect 18052 12801 18061 12835
rect 18061 12801 18095 12835
rect 18095 12801 18104 12835
rect 18052 12792 18104 12801
rect 20168 12792 20220 12844
rect 20444 12835 20496 12844
rect 20444 12801 20453 12835
rect 20453 12801 20487 12835
rect 20487 12801 20496 12835
rect 20444 12792 20496 12801
rect 20536 12835 20588 12844
rect 20536 12801 20545 12835
rect 20545 12801 20579 12835
rect 20579 12801 20588 12835
rect 20536 12792 20588 12801
rect 21732 12928 21784 12980
rect 25136 12928 25188 12980
rect 28080 12928 28132 12980
rect 28540 12928 28592 12980
rect 31576 12971 31628 12980
rect 31576 12937 31585 12971
rect 31585 12937 31619 12971
rect 31619 12937 31628 12971
rect 31576 12928 31628 12937
rect 32772 12928 32824 12980
rect 33048 12928 33100 12980
rect 37648 12971 37700 12980
rect 37648 12937 37657 12971
rect 37657 12937 37691 12971
rect 37691 12937 37700 12971
rect 37648 12928 37700 12937
rect 25780 12860 25832 12912
rect 26332 12835 26384 12844
rect 26332 12801 26341 12835
rect 26341 12801 26375 12835
rect 26375 12801 26384 12835
rect 26332 12792 26384 12801
rect 31116 12860 31168 12912
rect 31852 12860 31904 12912
rect 31944 12860 31996 12912
rect 32312 12860 32364 12912
rect 2412 12588 2464 12640
rect 7012 12656 7064 12708
rect 14004 12656 14056 12708
rect 15016 12656 15068 12708
rect 15200 12656 15252 12708
rect 10968 12588 11020 12640
rect 15108 12588 15160 12640
rect 17316 12588 17368 12640
rect 17684 12588 17736 12640
rect 29368 12724 29420 12776
rect 29920 12835 29972 12844
rect 29920 12801 29929 12835
rect 29929 12801 29963 12835
rect 29963 12801 29972 12835
rect 29920 12792 29972 12801
rect 30380 12792 30432 12844
rect 30932 12792 30984 12844
rect 31208 12835 31260 12844
rect 31208 12801 31217 12835
rect 31217 12801 31251 12835
rect 31251 12801 31260 12835
rect 31208 12792 31260 12801
rect 31392 12835 31444 12844
rect 31392 12801 31401 12835
rect 31401 12801 31435 12835
rect 31435 12801 31444 12835
rect 31392 12792 31444 12801
rect 32128 12792 32180 12844
rect 37096 12860 37148 12912
rect 32588 12835 32640 12844
rect 32588 12801 32597 12835
rect 32597 12801 32631 12835
rect 32631 12801 32640 12835
rect 32588 12792 32640 12801
rect 30380 12656 30432 12708
rect 32864 12792 32916 12844
rect 35808 12835 35860 12844
rect 35808 12801 35817 12835
rect 35817 12801 35851 12835
rect 35851 12801 35860 12835
rect 35808 12792 35860 12801
rect 36268 12792 36320 12844
rect 36820 12792 36872 12844
rect 37556 12792 37608 12844
rect 40040 12792 40092 12844
rect 35624 12724 35676 12776
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 27252 12588 27304 12640
rect 29460 12631 29512 12640
rect 29460 12597 29469 12631
rect 29469 12597 29503 12631
rect 29503 12597 29512 12631
rect 29460 12588 29512 12597
rect 32588 12588 32640 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 5816 12384 5868 12436
rect 10508 12427 10560 12436
rect 3424 12248 3476 12300
rect 10508 12393 10517 12427
rect 10517 12393 10551 12427
rect 10551 12393 10560 12427
rect 10508 12384 10560 12393
rect 15476 12427 15528 12436
rect 6920 12316 6972 12368
rect 8116 12316 8168 12368
rect 9772 12316 9824 12368
rect 8484 12248 8536 12300
rect 3148 12180 3200 12232
rect 5816 12223 5868 12232
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 5908 12180 5960 12232
rect 6000 12180 6052 12232
rect 6460 12180 6512 12232
rect 8392 12180 8444 12232
rect 9404 12180 9456 12232
rect 2228 12112 2280 12164
rect 5448 12112 5500 12164
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 17592 12384 17644 12436
rect 20536 12384 20588 12436
rect 20720 12384 20772 12436
rect 29920 12427 29972 12436
rect 29920 12393 29929 12427
rect 29929 12393 29963 12427
rect 29963 12393 29972 12427
rect 29920 12384 29972 12393
rect 34428 12384 34480 12436
rect 35900 12384 35952 12436
rect 36360 12427 36412 12436
rect 36360 12393 36369 12427
rect 36369 12393 36403 12427
rect 36403 12393 36412 12427
rect 36360 12384 36412 12393
rect 37188 12384 37240 12436
rect 18420 12316 18472 12368
rect 23020 12316 23072 12368
rect 24400 12316 24452 12368
rect 32220 12316 32272 12368
rect 17684 12248 17736 12300
rect 11428 12180 11480 12232
rect 11796 12180 11848 12232
rect 5724 12044 5776 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 12256 12112 12308 12164
rect 13268 12180 13320 12232
rect 14096 12223 14148 12232
rect 14096 12189 14105 12223
rect 14105 12189 14139 12223
rect 14139 12189 14148 12223
rect 14096 12180 14148 12189
rect 14740 12180 14792 12232
rect 14648 12112 14700 12164
rect 11060 12044 11112 12096
rect 11428 12044 11480 12096
rect 12348 12044 12400 12096
rect 12992 12044 13044 12096
rect 17592 12180 17644 12232
rect 18052 12248 18104 12300
rect 22836 12248 22888 12300
rect 27344 12248 27396 12300
rect 16672 12155 16724 12164
rect 16672 12121 16681 12155
rect 16681 12121 16715 12155
rect 16715 12121 16724 12155
rect 16672 12112 16724 12121
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 18696 12180 18748 12232
rect 20076 12223 20128 12232
rect 20076 12189 20110 12223
rect 20110 12189 20128 12223
rect 20076 12180 20128 12189
rect 27620 12180 27672 12232
rect 30840 12223 30892 12232
rect 30840 12189 30849 12223
rect 30849 12189 30883 12223
rect 30883 12189 30892 12223
rect 30840 12180 30892 12189
rect 31392 12180 31444 12232
rect 34704 12248 34756 12300
rect 15844 12044 15896 12096
rect 16488 12044 16540 12096
rect 19432 12112 19484 12164
rect 20536 12112 20588 12164
rect 28816 12112 28868 12164
rect 30472 12112 30524 12164
rect 30748 12112 30800 12164
rect 17960 12044 18012 12096
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 20444 12044 20496 12096
rect 25688 12087 25740 12096
rect 25688 12053 25697 12087
rect 25697 12053 25731 12087
rect 25731 12053 25740 12087
rect 25688 12044 25740 12053
rect 32036 12112 32088 12164
rect 31208 12044 31260 12096
rect 31852 12087 31904 12096
rect 31852 12053 31861 12087
rect 31861 12053 31895 12087
rect 31895 12053 31904 12087
rect 31852 12044 31904 12053
rect 32588 12180 32640 12232
rect 35532 12316 35584 12368
rect 35440 12248 35492 12300
rect 35256 12180 35308 12232
rect 35624 12180 35676 12232
rect 34796 12112 34848 12164
rect 34888 12112 34940 12164
rect 38568 12044 38620 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 2228 11883 2280 11892
rect 2228 11849 2237 11883
rect 2237 11849 2271 11883
rect 2271 11849 2280 11883
rect 2228 11840 2280 11849
rect 3148 11840 3200 11892
rect 6920 11840 6972 11892
rect 7380 11840 7432 11892
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9128 11840 9180 11849
rect 12992 11840 13044 11892
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 15016 11840 15068 11892
rect 16488 11840 16540 11892
rect 8484 11772 8536 11824
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 3240 11704 3292 11756
rect 3148 11679 3200 11688
rect 3148 11645 3157 11679
rect 3157 11645 3191 11679
rect 3191 11645 3200 11679
rect 3148 11636 3200 11645
rect 4620 11568 4672 11620
rect 5356 11568 5408 11620
rect 6368 11704 6420 11756
rect 6644 11747 6696 11756
rect 6644 11713 6653 11747
rect 6653 11713 6687 11747
rect 6687 11713 6696 11747
rect 6644 11704 6696 11713
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 6000 11636 6052 11688
rect 7288 11636 7340 11688
rect 7380 11568 7432 11620
rect 10968 11704 11020 11756
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 15200 11772 15252 11824
rect 17684 11840 17736 11892
rect 20168 11840 20220 11892
rect 22836 11840 22888 11892
rect 23112 11840 23164 11892
rect 24492 11840 24544 11892
rect 27620 11840 27672 11892
rect 17224 11772 17276 11824
rect 17868 11772 17920 11824
rect 8668 11679 8720 11688
rect 8668 11645 8677 11679
rect 8677 11645 8711 11679
rect 8711 11645 8720 11679
rect 8668 11636 8720 11645
rect 14740 11636 14792 11688
rect 5632 11500 5684 11552
rect 6000 11500 6052 11552
rect 6368 11500 6420 11552
rect 7932 11500 7984 11552
rect 15292 11747 15344 11756
rect 15292 11713 15301 11747
rect 15301 11713 15335 11747
rect 15335 11713 15344 11747
rect 15292 11704 15344 11713
rect 17500 11704 17552 11756
rect 20444 11772 20496 11824
rect 28632 11840 28684 11892
rect 29460 11772 29512 11824
rect 18880 11704 18932 11756
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 23480 11704 23532 11756
rect 25780 11747 25832 11756
rect 25780 11713 25789 11747
rect 25789 11713 25823 11747
rect 25823 11713 25832 11747
rect 25780 11704 25832 11713
rect 28724 11704 28776 11756
rect 31484 11840 31536 11892
rect 31760 11840 31812 11892
rect 31300 11815 31352 11824
rect 31300 11781 31309 11815
rect 31309 11781 31343 11815
rect 31343 11781 31352 11815
rect 31300 11772 31352 11781
rect 31208 11747 31260 11756
rect 31208 11713 31217 11747
rect 31217 11713 31251 11747
rect 31251 11713 31260 11747
rect 31208 11704 31260 11713
rect 31392 11747 31444 11756
rect 31392 11713 31401 11747
rect 31401 11713 31435 11747
rect 31435 11713 31444 11747
rect 31392 11704 31444 11713
rect 32772 11747 32824 11756
rect 32772 11713 32781 11747
rect 32781 11713 32815 11747
rect 32815 11713 32824 11747
rect 32772 11704 32824 11713
rect 34888 11704 34940 11756
rect 36084 11747 36136 11756
rect 36084 11713 36093 11747
rect 36093 11713 36127 11747
rect 36127 11713 36136 11747
rect 36084 11704 36136 11713
rect 38292 11704 38344 11756
rect 15200 11636 15252 11688
rect 15016 11568 15068 11620
rect 15568 11500 15620 11552
rect 18328 11500 18380 11552
rect 18420 11500 18472 11552
rect 28816 11636 28868 11688
rect 33048 11636 33100 11688
rect 37740 11636 37792 11688
rect 38936 11636 38988 11688
rect 23388 11568 23440 11620
rect 58164 11611 58216 11620
rect 58164 11577 58173 11611
rect 58173 11577 58207 11611
rect 58207 11577 58216 11611
rect 58164 11568 58216 11577
rect 23020 11500 23072 11552
rect 35348 11500 35400 11552
rect 37280 11500 37332 11552
rect 39120 11500 39172 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3240 11339 3292 11348
rect 3240 11305 3249 11339
rect 3249 11305 3283 11339
rect 3283 11305 3292 11339
rect 3240 11296 3292 11305
rect 8668 11296 8720 11348
rect 14096 11296 14148 11348
rect 17224 11296 17276 11348
rect 17500 11339 17552 11348
rect 17500 11305 17509 11339
rect 17509 11305 17543 11339
rect 17543 11305 17552 11339
rect 17500 11296 17552 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 22376 11296 22428 11348
rect 24400 11339 24452 11348
rect 11152 11271 11204 11280
rect 11152 11237 11161 11271
rect 11161 11237 11195 11271
rect 11195 11237 11204 11271
rect 11152 11228 11204 11237
rect 4620 11203 4672 11212
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 5632 11203 5684 11212
rect 5632 11169 5641 11203
rect 5641 11169 5675 11203
rect 5675 11169 5684 11203
rect 5632 11160 5684 11169
rect 5908 11160 5960 11212
rect 6092 11160 6144 11212
rect 6644 11160 6696 11212
rect 15292 11228 15344 11280
rect 16948 11160 17000 11212
rect 17684 11160 17736 11212
rect 22928 11228 22980 11280
rect 24400 11305 24409 11339
rect 24409 11305 24443 11339
rect 24443 11305 24452 11339
rect 24400 11296 24452 11305
rect 26700 11296 26752 11348
rect 29736 11296 29788 11348
rect 32496 11296 32548 11348
rect 35900 11339 35952 11348
rect 35900 11305 35909 11339
rect 35909 11305 35943 11339
rect 35943 11305 35952 11339
rect 35900 11296 35952 11305
rect 28632 11228 28684 11280
rect 3056 11135 3108 11144
rect 3056 11101 3065 11135
rect 3065 11101 3099 11135
rect 3099 11101 3108 11135
rect 3056 11092 3108 11101
rect 6828 11135 6880 11144
rect 6828 11101 6837 11135
rect 6837 11101 6871 11135
rect 6871 11101 6880 11135
rect 6828 11092 6880 11101
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 22652 11160 22704 11212
rect 12624 11092 12676 11101
rect 4620 11024 4672 11076
rect 5540 11067 5592 11076
rect 5540 11033 5549 11067
rect 5549 11033 5583 11067
rect 5583 11033 5592 11067
rect 5540 11024 5592 11033
rect 5724 11024 5776 11076
rect 4252 10956 4304 11008
rect 7380 11024 7432 11076
rect 11520 11024 11572 11076
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 18696 11092 18748 11144
rect 22836 11135 22888 11144
rect 22836 11101 22845 11135
rect 22845 11101 22879 11135
rect 22879 11101 22888 11135
rect 22836 11092 22888 11101
rect 23020 11135 23072 11144
rect 23020 11101 23034 11135
rect 23034 11101 23068 11135
rect 23068 11101 23072 11135
rect 23020 11092 23072 11101
rect 23388 11092 23440 11144
rect 25780 11092 25832 11144
rect 34704 11228 34756 11280
rect 36360 11228 36412 11280
rect 38568 11228 38620 11280
rect 32772 11203 32824 11212
rect 29460 11092 29512 11144
rect 29736 11135 29788 11144
rect 29736 11101 29745 11135
rect 29745 11101 29779 11135
rect 29779 11101 29788 11135
rect 29736 11092 29788 11101
rect 32772 11169 32781 11203
rect 32781 11169 32815 11203
rect 32815 11169 32824 11203
rect 32772 11160 32824 11169
rect 32864 11160 32916 11212
rect 31852 11135 31904 11144
rect 31852 11101 31861 11135
rect 31861 11101 31895 11135
rect 31895 11101 31904 11135
rect 31852 11092 31904 11101
rect 18512 11024 18564 11076
rect 28724 11024 28776 11076
rect 30380 11024 30432 11076
rect 30472 11024 30524 11076
rect 31576 11024 31628 11076
rect 35256 11067 35308 11076
rect 35256 11033 35265 11067
rect 35265 11033 35299 11067
rect 35299 11033 35308 11067
rect 35256 11024 35308 11033
rect 35900 11092 35952 11144
rect 37188 11092 37240 11144
rect 37648 11024 37700 11076
rect 38936 11135 38988 11144
rect 38936 11101 38945 11135
rect 38945 11101 38979 11135
rect 38979 11101 38988 11135
rect 38936 11092 38988 11101
rect 39120 11092 39172 11144
rect 7196 10956 7248 11008
rect 11612 10956 11664 11008
rect 22284 10956 22336 11008
rect 35440 10956 35492 11008
rect 35900 10956 35952 11008
rect 39304 10999 39356 11008
rect 39304 10965 39313 10999
rect 39313 10965 39347 10999
rect 39347 10965 39356 10999
rect 39304 10956 39356 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 3056 10752 3108 10804
rect 12440 10752 12492 10804
rect 22468 10752 22520 10804
rect 23480 10752 23532 10804
rect 24768 10752 24820 10804
rect 27620 10752 27672 10804
rect 29184 10752 29236 10804
rect 30104 10795 30156 10804
rect 30104 10761 30113 10795
rect 30113 10761 30147 10795
rect 30147 10761 30156 10795
rect 30104 10752 30156 10761
rect 31024 10752 31076 10804
rect 32312 10752 32364 10804
rect 37648 10795 37700 10804
rect 5908 10684 5960 10736
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 5816 10616 5868 10668
rect 4620 10548 4672 10600
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 13176 10684 13228 10736
rect 21088 10684 21140 10736
rect 22560 10684 22612 10736
rect 28632 10727 28684 10736
rect 28632 10693 28641 10727
rect 28641 10693 28675 10727
rect 28675 10693 28684 10727
rect 28632 10684 28684 10693
rect 30380 10684 30432 10736
rect 31208 10727 31260 10736
rect 31208 10693 31217 10727
rect 31217 10693 31251 10727
rect 31251 10693 31260 10727
rect 31208 10684 31260 10693
rect 37648 10761 37657 10795
rect 37657 10761 37691 10795
rect 37691 10761 37700 10795
rect 37648 10752 37700 10761
rect 34704 10684 34756 10736
rect 38568 10684 38620 10736
rect 7840 10659 7892 10668
rect 7840 10625 7849 10659
rect 7849 10625 7883 10659
rect 7883 10625 7892 10659
rect 7840 10616 7892 10625
rect 11612 10659 11664 10668
rect 11612 10625 11621 10659
rect 11621 10625 11655 10659
rect 11655 10625 11664 10659
rect 11612 10616 11664 10625
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 17132 10616 17184 10668
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 20076 10616 20128 10668
rect 22008 10659 22060 10668
rect 9588 10548 9640 10600
rect 12532 10548 12584 10600
rect 18604 10548 18656 10600
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 23296 10616 23348 10668
rect 24032 10616 24084 10668
rect 24400 10659 24452 10668
rect 24400 10625 24409 10659
rect 24409 10625 24443 10659
rect 24443 10625 24452 10659
rect 24400 10616 24452 10625
rect 27620 10659 27672 10668
rect 27620 10625 27629 10659
rect 27629 10625 27663 10659
rect 27663 10625 27672 10659
rect 27620 10616 27672 10625
rect 21916 10548 21968 10600
rect 25228 10548 25280 10600
rect 27896 10548 27948 10600
rect 9312 10412 9364 10464
rect 12440 10412 12492 10464
rect 18512 10412 18564 10464
rect 23296 10480 23348 10532
rect 29552 10616 29604 10668
rect 29736 10616 29788 10668
rect 31116 10659 31168 10668
rect 31116 10625 31125 10659
rect 31125 10625 31159 10659
rect 31159 10625 31168 10659
rect 31116 10616 31168 10625
rect 31300 10548 31352 10600
rect 30564 10480 30616 10532
rect 31208 10480 31260 10532
rect 32220 10616 32272 10668
rect 32496 10659 32548 10668
rect 32496 10625 32505 10659
rect 32505 10625 32539 10659
rect 32539 10625 32548 10659
rect 32496 10616 32548 10625
rect 32956 10616 33008 10668
rect 34796 10659 34848 10668
rect 34796 10625 34830 10659
rect 34830 10625 34848 10659
rect 37280 10659 37332 10668
rect 34796 10616 34848 10625
rect 37280 10625 37289 10659
rect 37289 10625 37323 10659
rect 37323 10625 37332 10659
rect 37280 10616 37332 10625
rect 32864 10548 32916 10600
rect 37004 10548 37056 10600
rect 39304 10616 39356 10668
rect 24676 10412 24728 10464
rect 24952 10412 25004 10464
rect 34428 10480 34480 10532
rect 33232 10412 33284 10464
rect 35900 10455 35952 10464
rect 35900 10421 35909 10455
rect 35909 10421 35943 10455
rect 35943 10421 35952 10455
rect 35900 10412 35952 10421
rect 58164 10455 58216 10464
rect 58164 10421 58173 10455
rect 58173 10421 58207 10455
rect 58207 10421 58216 10455
rect 58164 10412 58216 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 11060 10208 11112 10260
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 6276 10004 6328 10056
rect 7196 10047 7248 10056
rect 7196 10013 7205 10047
rect 7205 10013 7239 10047
rect 7239 10013 7248 10047
rect 7196 10004 7248 10013
rect 19156 10140 19208 10192
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 12624 10072 12676 10124
rect 16580 10072 16632 10124
rect 21916 10208 21968 10260
rect 22560 10208 22612 10260
rect 24676 10208 24728 10260
rect 32220 10208 32272 10260
rect 32496 10251 32548 10260
rect 32496 10217 32505 10251
rect 32505 10217 32539 10251
rect 32539 10217 32548 10251
rect 32496 10208 32548 10217
rect 34796 10208 34848 10260
rect 22928 10072 22980 10124
rect 13268 10047 13320 10056
rect 4620 9936 4672 9988
rect 13268 10013 13277 10047
rect 13277 10013 13311 10047
rect 13311 10013 13320 10047
rect 13268 10004 13320 10013
rect 20812 10047 20864 10056
rect 20812 10013 20821 10047
rect 20821 10013 20855 10047
rect 20855 10013 20864 10047
rect 20812 10004 20864 10013
rect 22284 10004 22336 10056
rect 27712 10072 27764 10124
rect 29368 10140 29420 10192
rect 32312 10140 32364 10192
rect 34520 10140 34572 10192
rect 34980 10208 35032 10260
rect 12164 9979 12216 9988
rect 12164 9945 12173 9979
rect 12173 9945 12207 9979
rect 12207 9945 12216 9979
rect 12164 9936 12216 9945
rect 16580 9936 16632 9988
rect 19432 9936 19484 9988
rect 22100 9936 22152 9988
rect 2412 9911 2464 9920
rect 2412 9877 2421 9911
rect 2421 9877 2455 9911
rect 2455 9877 2464 9911
rect 2412 9868 2464 9877
rect 7288 9911 7340 9920
rect 7288 9877 7297 9911
rect 7297 9877 7331 9911
rect 7331 9877 7340 9911
rect 7288 9868 7340 9877
rect 9128 9868 9180 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 9680 9868 9732 9920
rect 13360 9868 13412 9920
rect 18880 9868 18932 9920
rect 19248 9868 19300 9920
rect 19340 9868 19392 9920
rect 21088 9868 21140 9920
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 22744 9936 22796 9988
rect 23388 9936 23440 9988
rect 24032 10004 24084 10056
rect 24676 10004 24728 10056
rect 26700 10004 26752 10056
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 29736 10072 29788 10124
rect 34980 10047 35032 10056
rect 27344 9979 27396 9988
rect 27344 9945 27353 9979
rect 27353 9945 27387 9979
rect 27387 9945 27396 9979
rect 27344 9936 27396 9945
rect 31116 9936 31168 9988
rect 31576 9979 31628 9988
rect 31576 9945 31585 9979
rect 31585 9945 31619 9979
rect 31619 9945 31628 9979
rect 31576 9936 31628 9945
rect 32128 9936 32180 9988
rect 23204 9911 23256 9920
rect 23204 9877 23213 9911
rect 23213 9877 23247 9911
rect 23247 9877 23256 9911
rect 23204 9868 23256 9877
rect 28540 9868 28592 9920
rect 34980 10013 34989 10047
rect 34989 10013 35023 10047
rect 35023 10013 35032 10047
rect 34980 10004 35032 10013
rect 37740 10140 37792 10192
rect 35440 10072 35492 10124
rect 35348 10047 35400 10056
rect 35348 10013 35357 10047
rect 35357 10013 35391 10047
rect 35391 10013 35400 10047
rect 38016 10072 38068 10124
rect 35348 10004 35400 10013
rect 36820 10047 36872 10056
rect 36820 10013 36829 10047
rect 36829 10013 36863 10047
rect 36863 10013 36872 10047
rect 36820 10004 36872 10013
rect 37280 10004 37332 10056
rect 35256 9868 35308 9920
rect 35348 9868 35400 9920
rect 36268 9868 36320 9920
rect 36544 9868 36596 9920
rect 37280 9911 37332 9920
rect 37280 9877 37289 9911
rect 37289 9877 37323 9911
rect 37323 9877 37332 9911
rect 37280 9868 37332 9877
rect 37464 9868 37516 9920
rect 38384 9936 38436 9988
rect 39948 9868 40000 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 9680 9707 9732 9716
rect 9680 9673 9689 9707
rect 9689 9673 9723 9707
rect 9723 9673 9732 9707
rect 9680 9664 9732 9673
rect 2412 9639 2464 9648
rect 2412 9605 2446 9639
rect 2446 9605 2464 9639
rect 2412 9596 2464 9605
rect 5264 9528 5316 9580
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 7840 9596 7892 9648
rect 7932 9596 7984 9648
rect 6368 9528 6420 9580
rect 7012 9528 7064 9580
rect 8208 9528 8260 9580
rect 8944 9528 8996 9580
rect 4620 9460 4672 9469
rect 5632 9460 5684 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 5540 9392 5592 9444
rect 10048 9596 10100 9648
rect 12164 9664 12216 9716
rect 22376 9664 22428 9716
rect 23664 9664 23716 9716
rect 28080 9664 28132 9716
rect 13452 9596 13504 9648
rect 12440 9571 12492 9580
rect 12440 9537 12474 9571
rect 12474 9537 12492 9571
rect 12440 9528 12492 9537
rect 10324 9503 10376 9512
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 10784 9503 10836 9512
rect 10784 9469 10793 9503
rect 10793 9469 10827 9503
rect 10827 9469 10836 9503
rect 10784 9460 10836 9469
rect 18144 9596 18196 9648
rect 14556 9528 14608 9580
rect 17960 9460 18012 9512
rect 20168 9596 20220 9648
rect 19340 9528 19392 9580
rect 19984 9571 20036 9580
rect 19984 9537 19993 9571
rect 19993 9537 20027 9571
rect 20027 9537 20036 9571
rect 19984 9528 20036 9537
rect 25596 9596 25648 9648
rect 23204 9528 23256 9580
rect 20444 9503 20496 9512
rect 20444 9469 20453 9503
rect 20453 9469 20487 9503
rect 20487 9469 20496 9503
rect 20444 9460 20496 9469
rect 3976 9367 4028 9376
rect 3976 9333 3985 9367
rect 3985 9333 4019 9367
rect 4019 9333 4028 9367
rect 3976 9324 4028 9333
rect 5264 9367 5316 9376
rect 5264 9333 5273 9367
rect 5273 9333 5307 9367
rect 5307 9333 5316 9367
rect 5264 9324 5316 9333
rect 13176 9324 13228 9376
rect 14556 9367 14608 9376
rect 14556 9333 14565 9367
rect 14565 9333 14599 9367
rect 14599 9333 14608 9367
rect 14556 9324 14608 9333
rect 15384 9324 15436 9376
rect 16856 9324 16908 9376
rect 19432 9392 19484 9444
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 24768 9528 24820 9580
rect 25320 9571 25372 9580
rect 25320 9537 25329 9571
rect 25329 9537 25363 9571
rect 25363 9537 25372 9571
rect 25320 9528 25372 9537
rect 25504 9571 25556 9580
rect 25504 9537 25513 9571
rect 25513 9537 25547 9571
rect 25547 9537 25556 9571
rect 25504 9528 25556 9537
rect 31576 9596 31628 9648
rect 33232 9639 33284 9648
rect 33232 9605 33250 9639
rect 33250 9605 33284 9639
rect 33232 9596 33284 9605
rect 30380 9528 30432 9580
rect 27988 9460 28040 9512
rect 28908 9460 28960 9512
rect 25320 9392 25372 9444
rect 27804 9392 27856 9444
rect 23296 9324 23348 9376
rect 24032 9367 24084 9376
rect 24032 9333 24041 9367
rect 24041 9333 24075 9367
rect 24075 9333 24084 9367
rect 24032 9324 24084 9333
rect 25412 9324 25464 9376
rect 26148 9324 26200 9376
rect 27344 9324 27396 9376
rect 32128 9367 32180 9376
rect 32128 9333 32137 9367
rect 32137 9333 32171 9367
rect 32171 9333 32180 9367
rect 32128 9324 32180 9333
rect 32772 9324 32824 9376
rect 34704 9664 34756 9716
rect 35900 9596 35952 9648
rect 35992 9596 36044 9648
rect 36636 9664 36688 9716
rect 37280 9664 37332 9716
rect 39948 9707 40000 9716
rect 34704 9571 34756 9580
rect 34704 9537 34713 9571
rect 34713 9537 34747 9571
rect 34747 9537 34756 9571
rect 34704 9528 34756 9537
rect 34796 9528 34848 9580
rect 36268 9571 36320 9580
rect 35440 9460 35492 9512
rect 35624 9460 35676 9512
rect 36268 9537 36277 9571
rect 36277 9537 36311 9571
rect 36311 9537 36320 9571
rect 36268 9528 36320 9537
rect 37188 9528 37240 9580
rect 37280 9460 37332 9512
rect 37464 9392 37516 9444
rect 37727 9577 37779 9583
rect 37727 9543 37736 9577
rect 37736 9543 37770 9577
rect 37770 9543 37779 9577
rect 37727 9531 37779 9543
rect 39948 9673 39957 9707
rect 39957 9673 39991 9707
rect 39991 9673 40000 9707
rect 39948 9664 40000 9673
rect 38568 9571 38620 9580
rect 38568 9537 38577 9571
rect 38577 9537 38611 9571
rect 38611 9537 38620 9571
rect 38568 9528 38620 9537
rect 36636 9324 36688 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2596 9120 2648 9172
rect 8944 9163 8996 9172
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 3884 9052 3936 9104
rect 3976 8984 4028 9036
rect 4712 8984 4764 9036
rect 6828 8984 6880 9036
rect 4620 8916 4672 8968
rect 6276 8916 6328 8968
rect 5724 8848 5776 8900
rect 7196 8916 7248 8968
rect 7380 8916 7432 8968
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 10324 8984 10376 9036
rect 10784 9027 10836 9036
rect 10784 8993 10793 9027
rect 10793 8993 10827 9027
rect 10827 8993 10836 9027
rect 10784 8984 10836 8993
rect 12532 9052 12584 9104
rect 6736 8848 6788 8900
rect 13268 9120 13320 9172
rect 15568 9120 15620 9172
rect 18604 9163 18656 9172
rect 18604 9129 18613 9163
rect 18613 9129 18647 9163
rect 18647 9129 18656 9163
rect 18604 9120 18656 9129
rect 23204 9120 23256 9172
rect 24124 9120 24176 9172
rect 25320 9120 25372 9172
rect 28264 9120 28316 9172
rect 28632 9120 28684 9172
rect 31116 9120 31168 9172
rect 38016 9120 38068 9172
rect 12808 8984 12860 9036
rect 17224 9027 17276 9036
rect 17224 8993 17233 9027
rect 17233 8993 17267 9027
rect 17267 8993 17276 9027
rect 17224 8984 17276 8993
rect 13176 8916 13228 8968
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 13452 8916 13504 8968
rect 14924 8916 14976 8968
rect 19984 8984 20036 9036
rect 20444 8984 20496 9036
rect 23940 9052 23992 9104
rect 25044 9052 25096 9104
rect 25504 9052 25556 9104
rect 19248 8959 19300 8968
rect 11980 8848 12032 8900
rect 12072 8848 12124 8900
rect 4988 8780 5040 8832
rect 6920 8780 6972 8832
rect 11152 8780 11204 8832
rect 11244 8780 11296 8832
rect 12532 8780 12584 8832
rect 13544 8823 13596 8832
rect 13544 8789 13553 8823
rect 13553 8789 13587 8823
rect 13587 8789 13596 8823
rect 13544 8780 13596 8789
rect 15476 8848 15528 8900
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 19432 8959 19484 8968
rect 19432 8925 19441 8959
rect 19441 8925 19475 8959
rect 19475 8925 19484 8959
rect 19432 8916 19484 8925
rect 21272 8916 21324 8968
rect 24032 8984 24084 9036
rect 25596 9027 25648 9036
rect 25596 8993 25605 9027
rect 25605 8993 25639 9027
rect 25639 8993 25648 9027
rect 25596 8984 25648 8993
rect 27712 8984 27764 9036
rect 36360 9027 36412 9036
rect 36360 8993 36369 9027
rect 36369 8993 36403 9027
rect 36403 8993 36412 9027
rect 36360 8984 36412 8993
rect 23296 8959 23348 8968
rect 23296 8925 23305 8959
rect 23305 8925 23339 8959
rect 23339 8925 23348 8959
rect 23296 8916 23348 8925
rect 18052 8848 18104 8900
rect 18512 8848 18564 8900
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 16856 8780 16908 8832
rect 19156 8780 19208 8832
rect 19340 8823 19392 8832
rect 19340 8789 19349 8823
rect 19349 8789 19383 8823
rect 19383 8789 19392 8823
rect 19340 8780 19392 8789
rect 21180 8848 21232 8900
rect 22008 8848 22060 8900
rect 27804 8916 27856 8968
rect 27988 8916 28040 8968
rect 29828 8959 29880 8968
rect 29828 8925 29837 8959
rect 29837 8925 29871 8959
rect 29871 8925 29880 8959
rect 29828 8916 29880 8925
rect 36636 8959 36688 8968
rect 36636 8925 36670 8959
rect 36670 8925 36688 8959
rect 36636 8916 36688 8925
rect 58164 8959 58216 8968
rect 58164 8925 58173 8959
rect 58173 8925 58207 8959
rect 58207 8925 58216 8959
rect 58164 8916 58216 8925
rect 25872 8891 25924 8900
rect 25872 8857 25906 8891
rect 25906 8857 25924 8891
rect 25872 8848 25924 8857
rect 29000 8848 29052 8900
rect 25320 8780 25372 8832
rect 25504 8780 25556 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 3792 8508 3844 8560
rect 6184 8576 6236 8628
rect 7840 8576 7892 8628
rect 12808 8576 12860 8628
rect 5540 8483 5592 8492
rect 3240 8415 3292 8424
rect 3240 8381 3249 8415
rect 3249 8381 3283 8415
rect 3283 8381 3292 8415
rect 3240 8372 3292 8381
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 1768 8304 1820 8356
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 5632 8483 5684 8492
rect 5632 8449 5641 8483
rect 5641 8449 5675 8483
rect 5675 8449 5684 8483
rect 7196 8508 7248 8560
rect 7472 8508 7524 8560
rect 15016 8576 15068 8628
rect 15568 8619 15620 8628
rect 5632 8440 5684 8449
rect 6736 8440 6788 8492
rect 4620 8372 4672 8424
rect 5356 8372 5408 8424
rect 3976 8347 4028 8356
rect 3976 8313 3985 8347
rect 3985 8313 4019 8347
rect 4019 8313 4028 8347
rect 3976 8304 4028 8313
rect 6276 8372 6328 8424
rect 11796 8440 11848 8492
rect 7564 8372 7616 8424
rect 12532 8415 12584 8424
rect 12532 8381 12541 8415
rect 12541 8381 12575 8415
rect 12575 8381 12584 8415
rect 12532 8372 12584 8381
rect 13544 8440 13596 8492
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 18052 8619 18104 8628
rect 18052 8585 18061 8619
rect 18061 8585 18095 8619
rect 18095 8585 18104 8619
rect 18052 8576 18104 8585
rect 18144 8576 18196 8628
rect 18696 8576 18748 8628
rect 23112 8576 23164 8628
rect 24676 8576 24728 8628
rect 25872 8619 25924 8628
rect 16764 8508 16816 8560
rect 18328 8483 18380 8492
rect 13912 8372 13964 8424
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 15108 8372 15160 8424
rect 16580 8372 16632 8424
rect 18328 8449 18337 8483
rect 18337 8449 18371 8483
rect 18371 8449 18380 8483
rect 18328 8440 18380 8449
rect 18512 8483 18564 8492
rect 18512 8449 18521 8483
rect 18521 8449 18555 8483
rect 18555 8449 18564 8483
rect 18512 8440 18564 8449
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 21180 8440 21232 8492
rect 25044 8508 25096 8560
rect 25872 8585 25881 8619
rect 25881 8585 25915 8619
rect 25915 8585 25924 8619
rect 25872 8576 25924 8585
rect 22560 8440 22612 8492
rect 23480 8440 23532 8492
rect 23940 8440 23992 8492
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25412 8483 25464 8492
rect 25412 8449 25421 8483
rect 25421 8449 25455 8483
rect 25455 8449 25464 8483
rect 25412 8440 25464 8449
rect 25688 8508 25740 8560
rect 27896 8576 27948 8628
rect 28632 8576 28684 8628
rect 29000 8619 29052 8628
rect 27160 8508 27212 8560
rect 19340 8372 19392 8424
rect 19524 8372 19576 8424
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 23204 8372 23256 8424
rect 24768 8372 24820 8424
rect 27436 8440 27488 8492
rect 27804 8440 27856 8492
rect 28540 8483 28592 8492
rect 28540 8449 28549 8483
rect 28549 8449 28583 8483
rect 28583 8449 28592 8483
rect 28540 8440 28592 8449
rect 29000 8585 29009 8619
rect 29009 8585 29043 8619
rect 29043 8585 29052 8619
rect 29000 8576 29052 8585
rect 30012 8619 30064 8628
rect 30012 8585 30021 8619
rect 30021 8585 30055 8619
rect 30055 8585 30064 8619
rect 30012 8576 30064 8585
rect 28908 8508 28960 8560
rect 32128 8508 32180 8560
rect 27988 8372 28040 8424
rect 28816 8440 28868 8492
rect 29552 8440 29604 8492
rect 34520 8483 34572 8492
rect 8392 8347 8444 8356
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 2780 8236 2832 8245
rect 4068 8236 4120 8288
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 8392 8313 8401 8347
rect 8401 8313 8435 8347
rect 8435 8313 8444 8347
rect 8392 8304 8444 8313
rect 6920 8236 6972 8288
rect 9220 8236 9272 8288
rect 10416 8304 10468 8356
rect 18788 8304 18840 8356
rect 19156 8304 19208 8356
rect 24676 8347 24728 8356
rect 24676 8313 24685 8347
rect 24685 8313 24719 8347
rect 24719 8313 24728 8347
rect 24676 8304 24728 8313
rect 25228 8304 25280 8356
rect 27160 8304 27212 8356
rect 27712 8304 27764 8356
rect 27896 8304 27948 8356
rect 34520 8449 34529 8483
rect 34529 8449 34563 8483
rect 34563 8449 34572 8483
rect 34520 8440 34572 8449
rect 35992 8508 36044 8560
rect 34704 8483 34756 8492
rect 34704 8449 34713 8483
rect 34713 8449 34747 8483
rect 34747 8449 34756 8483
rect 34704 8440 34756 8449
rect 35624 8440 35676 8492
rect 11980 8236 12032 8288
rect 12440 8236 12492 8288
rect 15568 8236 15620 8288
rect 22008 8236 22060 8288
rect 22100 8236 22152 8288
rect 27436 8236 27488 8288
rect 28080 8236 28132 8288
rect 34244 8279 34296 8288
rect 34244 8245 34253 8279
rect 34253 8245 34287 8279
rect 34287 8245 34296 8279
rect 34244 8236 34296 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1584 7896 1636 7948
rect 4068 8032 4120 8084
rect 5540 8032 5592 8084
rect 9956 8032 10008 8084
rect 13268 8075 13320 8084
rect 2780 7828 2832 7880
rect 2872 7760 2924 7812
rect 6460 7964 6512 8016
rect 3332 7896 3384 7948
rect 5816 7939 5868 7948
rect 5816 7905 5825 7939
rect 5825 7905 5859 7939
rect 5859 7905 5868 7939
rect 5816 7896 5868 7905
rect 6736 7896 6788 7948
rect 4712 7828 4764 7880
rect 5724 7871 5776 7880
rect 5724 7837 5733 7871
rect 5733 7837 5767 7871
rect 5767 7837 5776 7871
rect 5724 7828 5776 7837
rect 5908 7871 5960 7880
rect 5908 7837 5917 7871
rect 5917 7837 5951 7871
rect 5951 7837 5960 7871
rect 5908 7828 5960 7837
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 3240 7760 3292 7812
rect 3976 7760 4028 7812
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 9496 7828 9548 7880
rect 11612 7964 11664 8016
rect 11152 7939 11204 7948
rect 11152 7905 11161 7939
rect 11161 7905 11195 7939
rect 11195 7905 11204 7939
rect 11152 7896 11204 7905
rect 12440 7939 12492 7948
rect 12440 7905 12449 7939
rect 12449 7905 12483 7939
rect 12483 7905 12492 7939
rect 12440 7896 12492 7905
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 5816 7692 5868 7744
rect 6184 7692 6236 7744
rect 8392 7760 8444 7812
rect 7196 7735 7248 7744
rect 7196 7701 7205 7735
rect 7205 7701 7239 7735
rect 7239 7701 7248 7735
rect 7196 7692 7248 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 8484 7692 8536 7744
rect 11244 7760 11296 7812
rect 11980 7828 12032 7880
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 13268 8041 13277 8075
rect 13277 8041 13311 8075
rect 13311 8041 13320 8075
rect 13268 8032 13320 8041
rect 15016 8032 15068 8084
rect 18144 8032 18196 8084
rect 18512 8032 18564 8084
rect 23572 8032 23624 8084
rect 28724 8032 28776 8084
rect 34704 8075 34756 8084
rect 34704 8041 34713 8075
rect 34713 8041 34747 8075
rect 34747 8041 34756 8075
rect 34704 8032 34756 8041
rect 19248 7964 19300 8016
rect 34796 7964 34848 8016
rect 37372 7964 37424 8016
rect 17132 7896 17184 7948
rect 32772 7939 32824 7948
rect 13912 7828 13964 7880
rect 15108 7828 15160 7880
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 18604 7828 18656 7880
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 32772 7905 32781 7939
rect 32781 7905 32815 7939
rect 32815 7905 32824 7939
rect 32772 7896 32824 7905
rect 22560 7871 22612 7880
rect 12624 7760 12676 7812
rect 18328 7760 18380 7812
rect 11152 7692 11204 7744
rect 11520 7735 11572 7744
rect 11520 7701 11529 7735
rect 11529 7701 11563 7735
rect 11563 7701 11572 7735
rect 11520 7692 11572 7701
rect 12808 7692 12860 7744
rect 14372 7692 14424 7744
rect 15568 7692 15620 7744
rect 17224 7735 17276 7744
rect 17224 7701 17233 7735
rect 17233 7701 17267 7735
rect 17267 7701 17276 7735
rect 17224 7692 17276 7701
rect 18788 7760 18840 7812
rect 22560 7837 22569 7871
rect 22569 7837 22603 7871
rect 22603 7837 22612 7871
rect 22560 7828 22612 7837
rect 23480 7828 23532 7880
rect 27068 7828 27120 7880
rect 29828 7828 29880 7880
rect 34244 7828 34296 7880
rect 34796 7828 34848 7880
rect 35348 7828 35400 7880
rect 35532 7828 35584 7880
rect 37188 7871 37240 7880
rect 37188 7837 37197 7871
rect 37197 7837 37231 7871
rect 37231 7837 37240 7871
rect 37188 7828 37240 7837
rect 37740 7896 37792 7948
rect 58164 7871 58216 7880
rect 24952 7760 25004 7812
rect 25688 7760 25740 7812
rect 27712 7803 27764 7812
rect 27712 7769 27746 7803
rect 27746 7769 27764 7803
rect 27712 7760 27764 7769
rect 19248 7735 19300 7744
rect 19248 7701 19257 7735
rect 19257 7701 19291 7735
rect 19291 7701 19300 7735
rect 19248 7692 19300 7701
rect 23296 7692 23348 7744
rect 25964 7692 26016 7744
rect 33784 7692 33836 7744
rect 58164 7837 58173 7871
rect 58173 7837 58207 7871
rect 58207 7837 58216 7871
rect 58164 7828 58216 7837
rect 37832 7735 37884 7744
rect 37832 7701 37841 7735
rect 37841 7701 37875 7735
rect 37875 7701 37884 7735
rect 37832 7692 37884 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 3976 7488 4028 7540
rect 7932 7488 7984 7540
rect 11060 7488 11112 7540
rect 12164 7531 12216 7540
rect 12164 7497 12173 7531
rect 12173 7497 12207 7531
rect 12207 7497 12216 7531
rect 12164 7488 12216 7497
rect 5908 7420 5960 7472
rect 11612 7463 11664 7472
rect 2136 7352 2188 7404
rect 2688 7395 2740 7404
rect 2688 7361 2722 7395
rect 2722 7361 2740 7395
rect 2688 7352 2740 7361
rect 7840 7352 7892 7404
rect 11612 7429 11621 7463
rect 11621 7429 11655 7463
rect 11655 7429 11664 7463
rect 11612 7420 11664 7429
rect 11244 7284 11296 7336
rect 12164 7216 12216 7268
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 14924 7352 14976 7404
rect 16764 7352 16816 7404
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 19432 7488 19484 7540
rect 21272 7531 21324 7540
rect 20812 7420 20864 7472
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 22560 7488 22612 7540
rect 24584 7488 24636 7540
rect 24768 7488 24820 7540
rect 27804 7488 27856 7540
rect 34428 7531 34480 7540
rect 34428 7497 34437 7531
rect 34437 7497 34471 7531
rect 34471 7497 34480 7531
rect 34428 7488 34480 7497
rect 34796 7488 34848 7540
rect 35808 7488 35860 7540
rect 37372 7488 37424 7540
rect 23296 7420 23348 7472
rect 19984 7352 20036 7404
rect 20720 7352 20772 7404
rect 17408 7284 17460 7336
rect 19432 7327 19484 7336
rect 19432 7293 19441 7327
rect 19441 7293 19475 7327
rect 19475 7293 19484 7327
rect 19432 7284 19484 7293
rect 18052 7216 18104 7268
rect 23388 7352 23440 7404
rect 24860 7420 24912 7472
rect 25688 7463 25740 7472
rect 25688 7429 25697 7463
rect 25697 7429 25731 7463
rect 25731 7429 25740 7463
rect 25688 7420 25740 7429
rect 26792 7420 26844 7472
rect 31024 7463 31076 7472
rect 31024 7429 31033 7463
rect 31033 7429 31067 7463
rect 31067 7429 31076 7463
rect 31024 7420 31076 7429
rect 34060 7420 34112 7472
rect 23204 7284 23256 7336
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 24400 7352 24452 7404
rect 24492 7352 24544 7404
rect 24768 7395 24820 7404
rect 24768 7361 24782 7395
rect 24782 7361 24816 7395
rect 24816 7361 24820 7395
rect 24768 7352 24820 7361
rect 23480 7216 23532 7268
rect 23664 7216 23716 7268
rect 24860 7216 24912 7268
rect 1952 7191 2004 7200
rect 1952 7157 1961 7191
rect 1961 7157 1995 7191
rect 1995 7157 2004 7191
rect 1952 7148 2004 7157
rect 4804 7191 4856 7200
rect 4804 7157 4813 7191
rect 4813 7157 4847 7191
rect 4847 7157 4856 7191
rect 4804 7148 4856 7157
rect 7656 7148 7708 7200
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 9588 7148 9640 7200
rect 14648 7148 14700 7200
rect 15292 7148 15344 7200
rect 15844 7148 15896 7200
rect 23572 7148 23624 7200
rect 24216 7148 24268 7200
rect 24400 7148 24452 7200
rect 25228 7352 25280 7404
rect 25872 7395 25924 7404
rect 25872 7361 25881 7395
rect 25881 7361 25915 7395
rect 25915 7361 25924 7395
rect 25872 7352 25924 7361
rect 26148 7352 26200 7404
rect 28724 7352 28776 7404
rect 35440 7420 35492 7472
rect 37188 7420 37240 7472
rect 34796 7395 34848 7404
rect 34796 7361 34805 7395
rect 34805 7361 34839 7395
rect 34839 7361 34848 7395
rect 34796 7352 34848 7361
rect 35348 7352 35400 7404
rect 35808 7395 35860 7404
rect 35808 7361 35817 7395
rect 35817 7361 35851 7395
rect 35851 7361 35860 7395
rect 35808 7352 35860 7361
rect 35992 7395 36044 7404
rect 35992 7361 36001 7395
rect 36001 7361 36035 7395
rect 36035 7361 36044 7395
rect 35992 7352 36044 7361
rect 36084 7352 36136 7404
rect 36728 7395 36780 7404
rect 36728 7361 36737 7395
rect 36737 7361 36771 7395
rect 36771 7361 36780 7395
rect 36728 7352 36780 7361
rect 37096 7352 37148 7404
rect 37464 7395 37516 7404
rect 37464 7361 37468 7395
rect 37468 7361 37502 7395
rect 37502 7361 37516 7395
rect 37464 7352 37516 7361
rect 37924 7352 37976 7404
rect 38384 7395 38436 7404
rect 38384 7361 38393 7395
rect 38393 7361 38427 7395
rect 38427 7361 38436 7395
rect 38384 7352 38436 7361
rect 25136 7216 25188 7268
rect 29828 7148 29880 7200
rect 30196 7148 30248 7200
rect 37740 7216 37792 7268
rect 39120 7284 39172 7336
rect 38016 7148 38068 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 2688 6944 2740 6996
rect 20812 6944 20864 6996
rect 22008 6944 22060 6996
rect 24492 6987 24544 6996
rect 24492 6953 24501 6987
rect 24501 6953 24535 6987
rect 24535 6953 24544 6987
rect 24492 6944 24544 6953
rect 27252 6944 27304 6996
rect 36084 6944 36136 6996
rect 2412 6808 2464 6860
rect 6092 6808 6144 6860
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 9496 6876 9548 6928
rect 7196 6808 7248 6860
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7840 6851 7892 6860
rect 7472 6808 7524 6817
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8024 6808 8076 6860
rect 14924 6876 14976 6928
rect 7656 6783 7708 6792
rect 7196 6672 7248 6724
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8208 6740 8260 6792
rect 3056 6604 3108 6656
rect 3976 6647 4028 6656
rect 3976 6613 3985 6647
rect 3985 6613 4019 6647
rect 4019 6613 4028 6647
rect 3976 6604 4028 6613
rect 4620 6604 4672 6656
rect 5448 6604 5500 6656
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6000 6604 6052 6613
rect 6552 6647 6604 6656
rect 6552 6613 6561 6647
rect 6561 6613 6595 6647
rect 6595 6613 6604 6647
rect 6552 6604 6604 6613
rect 8668 6672 8720 6724
rect 8852 6604 8904 6656
rect 15476 6808 15528 6860
rect 9496 6740 9548 6792
rect 11244 6783 11296 6792
rect 11244 6749 11253 6783
rect 11253 6749 11287 6783
rect 11287 6749 11296 6783
rect 11244 6740 11296 6749
rect 13084 6740 13136 6792
rect 34060 6851 34112 6860
rect 34060 6817 34069 6851
rect 34069 6817 34103 6851
rect 34103 6817 34112 6851
rect 34060 6808 34112 6817
rect 11520 6715 11572 6724
rect 11520 6681 11554 6715
rect 11554 6681 11572 6715
rect 11520 6672 11572 6681
rect 14556 6672 14608 6724
rect 15844 6783 15896 6792
rect 15844 6749 15853 6783
rect 15853 6749 15887 6783
rect 15887 6749 15896 6783
rect 15844 6740 15896 6749
rect 15292 6672 15344 6724
rect 17132 6740 17184 6792
rect 19248 6740 19300 6792
rect 22192 6740 22244 6792
rect 26792 6783 26844 6792
rect 16672 6715 16724 6724
rect 16672 6681 16681 6715
rect 16681 6681 16715 6715
rect 16715 6681 16724 6715
rect 16672 6672 16724 6681
rect 18052 6715 18104 6724
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 15108 6604 15160 6656
rect 18052 6681 18061 6715
rect 18061 6681 18095 6715
rect 18095 6681 18104 6715
rect 18052 6672 18104 6681
rect 26792 6749 26801 6783
rect 26801 6749 26835 6783
rect 26835 6749 26844 6783
rect 26792 6740 26844 6749
rect 28816 6740 28868 6792
rect 30196 6783 30248 6792
rect 30196 6749 30205 6783
rect 30205 6749 30239 6783
rect 30239 6749 30248 6783
rect 30196 6740 30248 6749
rect 32772 6740 32824 6792
rect 29276 6672 29328 6724
rect 30748 6672 30800 6724
rect 38016 6740 38068 6792
rect 37280 6672 37332 6724
rect 17040 6604 17092 6656
rect 17868 6604 17920 6656
rect 18696 6604 18748 6656
rect 20444 6604 20496 6656
rect 25596 6604 25648 6656
rect 27436 6604 27488 6656
rect 29184 6604 29236 6656
rect 30564 6604 30616 6656
rect 31484 6604 31536 6656
rect 37188 6604 37240 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4896 6400 4948 6452
rect 8024 6400 8076 6452
rect 4068 6332 4120 6384
rect 2412 6307 2464 6316
rect 2412 6273 2421 6307
rect 2421 6273 2455 6307
rect 2455 6273 2464 6307
rect 2412 6264 2464 6273
rect 5172 6264 5224 6316
rect 7288 6332 7340 6384
rect 7840 6332 7892 6384
rect 5724 6264 5776 6316
rect 6000 6264 6052 6316
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 3884 6196 3936 6248
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 6460 6264 6512 6316
rect 8024 6264 8076 6316
rect 15200 6400 15252 6452
rect 15568 6400 15620 6452
rect 19984 6400 20036 6452
rect 24952 6400 25004 6452
rect 28816 6400 28868 6452
rect 30748 6443 30800 6452
rect 30748 6409 30757 6443
rect 30757 6409 30791 6443
rect 30791 6409 30800 6443
rect 30748 6400 30800 6409
rect 33784 6443 33836 6452
rect 33784 6409 33793 6443
rect 33793 6409 33827 6443
rect 33827 6409 33836 6443
rect 33784 6400 33836 6409
rect 35900 6400 35952 6452
rect 39120 6443 39172 6452
rect 39120 6409 39129 6443
rect 39129 6409 39163 6443
rect 39163 6409 39172 6443
rect 39120 6400 39172 6409
rect 12808 6375 12860 6384
rect 12808 6341 12826 6375
rect 12826 6341 12860 6375
rect 12808 6332 12860 6341
rect 8300 6264 8352 6316
rect 8760 6307 8812 6316
rect 8760 6273 8769 6307
rect 8769 6273 8803 6307
rect 8803 6273 8812 6307
rect 8760 6264 8812 6273
rect 8852 6264 8904 6316
rect 7564 6196 7616 6248
rect 13084 6307 13136 6316
rect 13084 6273 13093 6307
rect 13093 6273 13127 6307
rect 13127 6273 13136 6307
rect 13084 6264 13136 6273
rect 14464 6264 14516 6316
rect 15200 6307 15252 6316
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 17868 6332 17920 6384
rect 3516 6128 3568 6180
rect 2872 6060 2924 6112
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 5632 6128 5684 6180
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 8392 6128 8444 6180
rect 14924 6196 14976 6248
rect 15660 6264 15712 6316
rect 20720 6332 20772 6384
rect 21272 6332 21324 6384
rect 22192 6375 22244 6384
rect 22192 6341 22201 6375
rect 22201 6341 22235 6375
rect 22235 6341 22244 6375
rect 22192 6332 22244 6341
rect 20076 6307 20128 6316
rect 20076 6273 20085 6307
rect 20085 6273 20119 6307
rect 20119 6273 20128 6307
rect 20076 6264 20128 6273
rect 20444 6307 20496 6316
rect 17040 6196 17092 6248
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 19340 6239 19392 6248
rect 19340 6205 19349 6239
rect 19349 6205 19383 6239
rect 19383 6205 19392 6239
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 24860 6332 24912 6384
rect 25596 6332 25648 6384
rect 29276 6375 29328 6384
rect 29276 6341 29285 6375
rect 29285 6341 29319 6375
rect 29319 6341 29328 6375
rect 29276 6332 29328 6341
rect 31484 6332 31536 6384
rect 23572 6307 23624 6316
rect 23572 6273 23606 6307
rect 23606 6273 23624 6307
rect 23572 6264 23624 6273
rect 27068 6307 27120 6316
rect 27068 6273 27077 6307
rect 27077 6273 27111 6307
rect 27111 6273 27120 6307
rect 27068 6264 27120 6273
rect 27160 6264 27212 6316
rect 30012 6264 30064 6316
rect 19340 6196 19392 6205
rect 9312 6060 9364 6112
rect 10324 6060 10376 6112
rect 10508 6060 10560 6112
rect 11612 6060 11664 6112
rect 11980 6060 12032 6112
rect 18972 6128 19024 6180
rect 26976 6196 27028 6248
rect 30564 6264 30616 6316
rect 34796 6307 34848 6316
rect 34796 6273 34805 6307
rect 34805 6273 34839 6307
rect 34839 6273 34848 6307
rect 34796 6264 34848 6273
rect 35624 6264 35676 6316
rect 35900 6307 35952 6316
rect 35900 6273 35909 6307
rect 35909 6273 35943 6307
rect 35943 6273 35952 6307
rect 35900 6264 35952 6273
rect 37832 6332 37884 6384
rect 36084 6307 36136 6316
rect 36084 6273 36093 6307
rect 36093 6273 36127 6307
rect 36127 6273 36136 6307
rect 36084 6264 36136 6273
rect 37280 6264 37332 6316
rect 14648 6103 14700 6112
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 14648 6060 14700 6069
rect 15660 6060 15712 6112
rect 15752 6060 15804 6112
rect 20076 6060 20128 6112
rect 30472 6128 30524 6180
rect 58164 6171 58216 6180
rect 58164 6137 58173 6171
rect 58173 6137 58207 6171
rect 58207 6137 58216 6171
rect 58164 6128 58216 6137
rect 34336 6103 34388 6112
rect 34336 6069 34345 6103
rect 34345 6069 34379 6103
rect 34379 6069 34388 6103
rect 34336 6060 34388 6069
rect 37004 6060 37056 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 2136 5856 2188 5908
rect 5724 5899 5776 5908
rect 5724 5865 5733 5899
rect 5733 5865 5767 5899
rect 5767 5865 5776 5899
rect 5724 5856 5776 5865
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 7564 5856 7616 5908
rect 8024 5788 8076 5840
rect 9772 5856 9824 5908
rect 11888 5856 11940 5908
rect 10416 5788 10468 5840
rect 11796 5788 11848 5840
rect 17040 5899 17092 5908
rect 3608 5720 3660 5772
rect 6460 5720 6512 5772
rect 10600 5720 10652 5772
rect 14924 5788 14976 5840
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 19432 5856 19484 5908
rect 20444 5856 20496 5908
rect 24768 5856 24820 5908
rect 27160 5856 27212 5908
rect 18512 5788 18564 5840
rect 20904 5788 20956 5840
rect 4528 5652 4580 5704
rect 4896 5652 4948 5704
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 6828 5652 6880 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7104 5652 7156 5704
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9128 5652 9180 5704
rect 9680 5652 9732 5704
rect 10048 5695 10100 5704
rect 10048 5661 10054 5695
rect 10054 5661 10100 5695
rect 10048 5652 10100 5661
rect 11336 5652 11388 5704
rect 13360 5695 13412 5704
rect 2964 5584 3016 5636
rect 5448 5584 5500 5636
rect 7380 5584 7432 5636
rect 9864 5627 9916 5636
rect 9864 5593 9873 5627
rect 9873 5593 9907 5627
rect 9907 5593 9916 5627
rect 9864 5584 9916 5593
rect 10232 5584 10284 5636
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 14832 5695 14884 5704
rect 14832 5661 14841 5695
rect 14841 5661 14875 5695
rect 14875 5661 14884 5695
rect 14832 5652 14884 5661
rect 15108 5652 15160 5704
rect 15292 5652 15344 5704
rect 15752 5652 15804 5704
rect 19340 5720 19392 5772
rect 26976 5720 27028 5772
rect 20628 5652 20680 5704
rect 23480 5652 23532 5704
rect 25872 5652 25924 5704
rect 26240 5652 26292 5704
rect 27252 5695 27304 5704
rect 27252 5661 27261 5695
rect 27261 5661 27295 5695
rect 27295 5661 27304 5695
rect 27252 5652 27304 5661
rect 27436 5695 27488 5704
rect 27436 5661 27445 5695
rect 27445 5661 27479 5695
rect 27479 5661 27488 5695
rect 27436 5652 27488 5661
rect 17868 5584 17920 5636
rect 18512 5627 18564 5636
rect 4896 5516 4948 5568
rect 6276 5516 6328 5568
rect 6460 5516 6512 5568
rect 6828 5516 6880 5568
rect 7012 5516 7064 5568
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 18512 5593 18521 5627
rect 18521 5593 18555 5627
rect 18555 5593 18564 5627
rect 18512 5584 18564 5593
rect 21272 5584 21324 5636
rect 27160 5584 27212 5636
rect 29276 5652 29328 5704
rect 30840 5856 30892 5908
rect 34796 5856 34848 5908
rect 35900 5856 35952 5908
rect 37464 5856 37516 5908
rect 32772 5720 32824 5772
rect 35348 5652 35400 5704
rect 35992 5652 36044 5704
rect 37188 5695 37240 5704
rect 37188 5661 37197 5695
rect 37197 5661 37231 5695
rect 37231 5661 37240 5695
rect 37188 5652 37240 5661
rect 30840 5584 30892 5636
rect 35532 5584 35584 5636
rect 38384 5584 38436 5636
rect 19432 5516 19484 5568
rect 30380 5516 30432 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 6368 5312 6420 5364
rect 8576 5312 8628 5364
rect 1584 5244 1636 5296
rect 2136 5244 2188 5296
rect 4620 5244 4672 5296
rect 6460 5244 6512 5296
rect 11704 5244 11756 5296
rect 14832 5312 14884 5364
rect 16672 5312 16724 5364
rect 19340 5312 19392 5364
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 5172 5176 5224 5228
rect 6276 5176 6328 5228
rect 6920 5176 6972 5228
rect 7564 5176 7616 5228
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 8668 5176 8720 5228
rect 10784 5176 10836 5228
rect 6644 5151 6696 5160
rect 6644 5117 6653 5151
rect 6653 5117 6687 5151
rect 6687 5117 6696 5151
rect 6644 5108 6696 5117
rect 10416 5108 10468 5160
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 10876 5108 10928 5160
rect 11060 5108 11112 5160
rect 7104 5083 7156 5092
rect 7104 5049 7113 5083
rect 7113 5049 7147 5083
rect 7147 5049 7156 5083
rect 7104 5040 7156 5049
rect 10048 5083 10100 5092
rect 10048 5049 10057 5083
rect 10057 5049 10091 5083
rect 10091 5049 10100 5083
rect 10048 5040 10100 5049
rect 1676 4972 1728 5024
rect 5632 4972 5684 5024
rect 6184 4972 6236 5024
rect 9864 4972 9916 5024
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 10600 4972 10652 5024
rect 11796 4972 11848 5024
rect 11888 4972 11940 5024
rect 12072 4972 12124 5024
rect 14556 5244 14608 5296
rect 14464 5176 14516 5228
rect 15292 5176 15344 5228
rect 16948 5108 17000 5160
rect 17868 5108 17920 5160
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 19248 5244 19300 5296
rect 19432 5244 19484 5296
rect 23480 5312 23532 5364
rect 30380 5312 30432 5364
rect 30840 5355 30892 5364
rect 30840 5321 30849 5355
rect 30849 5321 30883 5355
rect 30883 5321 30892 5355
rect 30840 5312 30892 5321
rect 36084 5312 36136 5364
rect 18880 5176 18932 5185
rect 19064 5108 19116 5160
rect 19984 5219 20036 5228
rect 19984 5185 19993 5219
rect 19993 5185 20027 5219
rect 20027 5185 20036 5219
rect 19984 5176 20036 5185
rect 20168 5176 20220 5228
rect 24216 5219 24268 5228
rect 24216 5185 24234 5219
rect 24234 5185 24268 5219
rect 24216 5176 24268 5185
rect 24860 5176 24912 5228
rect 30012 5176 30064 5228
rect 24952 5151 25004 5160
rect 24952 5117 24961 5151
rect 24961 5117 24995 5151
rect 24995 5117 25004 5151
rect 24952 5108 25004 5117
rect 27160 5108 27212 5160
rect 30288 5108 30340 5160
rect 19248 5040 19300 5092
rect 27436 5040 27488 5092
rect 29736 5040 29788 5092
rect 53748 5108 53800 5160
rect 54116 5040 54168 5092
rect 17960 4972 18012 5024
rect 18328 4972 18380 5024
rect 18880 4972 18932 5024
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 20260 5015 20312 5024
rect 20260 4981 20269 5015
rect 20269 4981 20303 5015
rect 20303 4981 20312 5015
rect 20260 4972 20312 4981
rect 25780 4972 25832 5024
rect 30564 4972 30616 5024
rect 53656 4972 53708 5024
rect 58164 5015 58216 5024
rect 58164 4981 58173 5015
rect 58173 4981 58207 5015
rect 58207 4981 58216 5015
rect 58164 4972 58216 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 3884 4768 3936 4820
rect 5356 4811 5408 4820
rect 5356 4777 5365 4811
rect 5365 4777 5399 4811
rect 5399 4777 5408 4811
rect 5356 4768 5408 4777
rect 6460 4811 6512 4820
rect 6460 4777 6469 4811
rect 6469 4777 6503 4811
rect 6503 4777 6512 4811
rect 6460 4768 6512 4777
rect 8300 4768 8352 4820
rect 10140 4768 10192 4820
rect 5264 4700 5316 4752
rect 7104 4700 7156 4752
rect 1952 4632 2004 4684
rect 10048 4700 10100 4752
rect 11520 4768 11572 4820
rect 11796 4768 11848 4820
rect 12716 4768 12768 4820
rect 10600 4743 10652 4752
rect 10600 4709 10609 4743
rect 10609 4709 10643 4743
rect 10643 4709 10652 4743
rect 10600 4700 10652 4709
rect 25780 4768 25832 4820
rect 16948 4743 17000 4752
rect 2596 4607 2648 4616
rect 2596 4573 2605 4607
rect 2605 4573 2639 4607
rect 2639 4573 2648 4607
rect 2596 4564 2648 4573
rect 3056 4607 3108 4616
rect 3056 4573 3057 4607
rect 3057 4573 3091 4607
rect 3091 4573 3108 4607
rect 3056 4564 3108 4573
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4804 4564 4856 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 6276 4564 6328 4616
rect 8944 4632 8996 4684
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 6736 4564 6788 4616
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 8024 4564 8076 4616
rect 8392 4564 8444 4616
rect 5264 4496 5316 4548
rect 8852 4496 8904 4548
rect 9220 4496 9272 4548
rect 10876 4632 10928 4684
rect 10416 4564 10468 4616
rect 11520 4564 11572 4616
rect 16948 4709 16957 4743
rect 16957 4709 16991 4743
rect 16991 4709 17000 4743
rect 16948 4700 17000 4709
rect 18328 4743 18380 4752
rect 18328 4709 18337 4743
rect 18337 4709 18371 4743
rect 18371 4709 18380 4743
rect 18328 4700 18380 4709
rect 21272 4743 21324 4752
rect 21272 4709 21281 4743
rect 21281 4709 21315 4743
rect 21315 4709 21324 4743
rect 21272 4700 21324 4709
rect 12256 4632 12308 4684
rect 12716 4564 12768 4616
rect 14096 4564 14148 4616
rect 19340 4564 19392 4616
rect 20628 4564 20680 4616
rect 2320 4428 2372 4480
rect 4620 4471 4672 4480
rect 4620 4437 4629 4471
rect 4629 4437 4663 4471
rect 4663 4437 4672 4471
rect 4620 4428 4672 4437
rect 5540 4428 5592 4480
rect 19156 4496 19208 4548
rect 13360 4428 13412 4480
rect 13452 4471 13504 4480
rect 13452 4437 13461 4471
rect 13461 4437 13495 4471
rect 13495 4437 13504 4471
rect 13452 4428 13504 4437
rect 17868 4428 17920 4480
rect 24952 4564 25004 4616
rect 21272 4496 21324 4548
rect 31208 4768 31260 4820
rect 35992 4768 36044 4820
rect 27160 4700 27212 4752
rect 27620 4632 27672 4684
rect 26056 4607 26108 4616
rect 26056 4573 26065 4607
rect 26065 4573 26099 4607
rect 26099 4573 26108 4607
rect 26056 4564 26108 4573
rect 26516 4564 26568 4616
rect 26884 4607 26936 4616
rect 26884 4573 26893 4607
rect 26893 4573 26927 4607
rect 26927 4573 26936 4607
rect 26884 4564 26936 4573
rect 27160 4607 27212 4616
rect 26332 4428 26384 4480
rect 27160 4573 27169 4607
rect 27169 4573 27203 4607
rect 27203 4573 27212 4607
rect 27160 4564 27212 4573
rect 29276 4632 29328 4684
rect 30564 4700 30616 4752
rect 52184 4700 52236 4752
rect 53932 4700 53984 4752
rect 30012 4607 30064 4616
rect 30012 4573 30021 4607
rect 30021 4573 30055 4607
rect 30055 4573 30064 4607
rect 30012 4564 30064 4573
rect 37280 4675 37332 4684
rect 37280 4641 37289 4675
rect 37289 4641 37323 4675
rect 37323 4641 37332 4675
rect 37280 4632 37332 4641
rect 53196 4632 53248 4684
rect 54300 4632 54352 4684
rect 30380 4607 30432 4616
rect 30380 4573 30389 4607
rect 30389 4573 30423 4607
rect 30423 4573 30432 4607
rect 30380 4564 30432 4573
rect 30656 4564 30708 4616
rect 30932 4564 30984 4616
rect 31576 4564 31628 4616
rect 37004 4607 37056 4616
rect 37004 4573 37022 4607
rect 37022 4573 37056 4607
rect 37004 4564 37056 4573
rect 52092 4564 52144 4616
rect 52644 4564 52696 4616
rect 30472 4496 30524 4548
rect 29000 4471 29052 4480
rect 29000 4437 29009 4471
rect 29009 4437 29043 4471
rect 29043 4437 29052 4471
rect 29000 4428 29052 4437
rect 29276 4428 29328 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 2596 4156 2648 4208
rect 3792 4224 3844 4276
rect 3976 4224 4028 4276
rect 5356 4156 5408 4208
rect 6828 4224 6880 4276
rect 7564 4267 7616 4276
rect 7564 4233 7573 4267
rect 7573 4233 7607 4267
rect 7607 4233 7616 4267
rect 7564 4224 7616 4233
rect 29000 4224 29052 4276
rect 30380 4224 30432 4276
rect 31576 4267 31628 4276
rect 31576 4233 31585 4267
rect 31585 4233 31619 4267
rect 31619 4233 31628 4267
rect 31576 4224 31628 4233
rect 6920 4156 6972 4208
rect 20260 4156 20312 4208
rect 30564 4156 30616 4208
rect 1676 4131 1728 4140
rect 1676 4097 1685 4131
rect 1685 4097 1719 4131
rect 1719 4097 1728 4131
rect 1676 4088 1728 4097
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 2412 4131 2464 4140
rect 2412 4097 2421 4131
rect 2421 4097 2455 4131
rect 2455 4097 2464 4131
rect 2412 4088 2464 4097
rect 2872 4088 2924 4140
rect 4068 4088 4120 4140
rect 6552 4088 6604 4140
rect 7288 4088 7340 4140
rect 7472 4088 7524 4140
rect 3516 4020 3568 4072
rect 4896 4020 4948 4072
rect 6368 4020 6420 4072
rect 2964 3995 3016 4004
rect 2964 3961 2973 3995
rect 2973 3961 3007 3995
rect 3007 3961 3016 3995
rect 2964 3952 3016 3961
rect 4528 3952 4580 4004
rect 4620 3952 4672 4004
rect 1952 3884 2004 3936
rect 5356 3884 5408 3936
rect 5724 3884 5776 3936
rect 6276 3884 6328 3936
rect 6644 3952 6696 4004
rect 8300 4088 8352 4140
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 11612 4088 11664 4140
rect 14740 4088 14792 4140
rect 19340 4131 19392 4140
rect 19340 4097 19349 4131
rect 19349 4097 19383 4131
rect 19383 4097 19392 4131
rect 19340 4088 19392 4097
rect 30196 4131 30248 4140
rect 30196 4097 30205 4131
rect 30205 4097 30239 4131
rect 30239 4097 30248 4131
rect 30196 4088 30248 4097
rect 32772 4088 32824 4140
rect 34336 4088 34388 4140
rect 53012 4088 53064 4140
rect 8392 4020 8444 4072
rect 10048 4020 10100 4072
rect 51816 4020 51868 4072
rect 54024 4020 54076 4072
rect 9312 3952 9364 4004
rect 35348 3952 35400 4004
rect 52828 3952 52880 4004
rect 8392 3884 8444 3936
rect 8576 3884 8628 3936
rect 8852 3884 8904 3936
rect 9220 3884 9272 3936
rect 11612 3884 11664 3936
rect 12164 3884 12216 3936
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 12440 3884 12492 3893
rect 13268 3884 13320 3936
rect 13820 3884 13872 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 14832 3927 14884 3936
rect 14832 3893 14841 3927
rect 14841 3893 14875 3927
rect 14875 3893 14884 3927
rect 14832 3884 14884 3893
rect 20904 3884 20956 3936
rect 29460 3884 29512 3936
rect 51080 3884 51132 3936
rect 51356 3884 51408 3936
rect 52460 3884 52512 3936
rect 55312 3927 55364 3936
rect 55312 3893 55321 3927
rect 55321 3893 55355 3927
rect 55355 3893 55364 3927
rect 55312 3884 55364 3893
rect 58440 3884 58492 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2136 3680 2188 3732
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 5632 3680 5684 3732
rect 7564 3680 7616 3732
rect 7656 3680 7708 3732
rect 8668 3680 8720 3732
rect 9128 3680 9180 3732
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 10968 3680 11020 3732
rect 26056 3680 26108 3732
rect 27620 3680 27672 3732
rect 52736 3680 52788 3732
rect 5448 3612 5500 3664
rect 6552 3612 6604 3664
rect 8300 3612 8352 3664
rect 6736 3544 6788 3596
rect 8668 3544 8720 3596
rect 11244 3612 11296 3664
rect 12256 3612 12308 3664
rect 14004 3612 14056 3664
rect 9496 3587 9548 3596
rect 9496 3553 9505 3587
rect 9505 3553 9539 3587
rect 9539 3553 9548 3587
rect 9496 3544 9548 3553
rect 13544 3544 13596 3596
rect 13912 3544 13964 3596
rect 46296 3612 46348 3664
rect 51448 3612 51500 3664
rect 24860 3544 24912 3596
rect 50804 3544 50856 3596
rect 51632 3544 51684 3596
rect 53840 3544 53892 3596
rect 1952 3476 2004 3528
rect 5080 3476 5132 3528
rect 5264 3476 5316 3528
rect 6460 3476 6512 3528
rect 8484 3476 8536 3528
rect 9036 3476 9088 3528
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 11152 3476 11204 3528
rect 12992 3476 13044 3528
rect 14188 3476 14240 3528
rect 15200 3476 15252 3528
rect 15936 3476 15988 3528
rect 16764 3476 16816 3528
rect 17592 3476 17644 3528
rect 18420 3476 18472 3528
rect 19432 3476 19484 3528
rect 20352 3476 20404 3528
rect 21180 3476 21232 3528
rect 22284 3476 22336 3528
rect 22560 3476 22612 3528
rect 23388 3476 23440 3528
rect 24492 3476 24544 3528
rect 25596 3519 25648 3528
rect 25596 3485 25605 3519
rect 25605 3485 25639 3519
rect 25639 3485 25648 3519
rect 25596 3476 25648 3485
rect 26332 3519 26384 3528
rect 26332 3485 26366 3519
rect 26366 3485 26384 3519
rect 26332 3476 26384 3485
rect 27528 3476 27580 3528
rect 28632 3476 28684 3528
rect 34704 3476 34756 3528
rect 35348 3476 35400 3528
rect 35808 3476 35860 3528
rect 36636 3476 36688 3528
rect 37464 3476 37516 3528
rect 38568 3476 38620 3528
rect 39948 3476 40000 3528
rect 40500 3476 40552 3528
rect 41052 3476 41104 3528
rect 42432 3476 42484 3528
rect 42708 3476 42760 3528
rect 44364 3476 44416 3528
rect 45192 3476 45244 3528
rect 46020 3476 46072 3528
rect 47676 3476 47728 3528
rect 48228 3476 48280 3528
rect 50160 3476 50212 3528
rect 50620 3476 50672 3528
rect 51172 3476 51224 3528
rect 52276 3476 52328 3528
rect 5724 3451 5776 3460
rect 5724 3417 5733 3451
rect 5733 3417 5767 3451
rect 5767 3417 5776 3451
rect 5724 3408 5776 3417
rect 6644 3408 6696 3460
rect 8392 3408 8444 3460
rect 2596 3340 2648 3392
rect 4068 3340 4120 3392
rect 5632 3340 5684 3392
rect 8024 3340 8076 3392
rect 11152 3340 11204 3392
rect 14832 3451 14884 3460
rect 14832 3417 14841 3451
rect 14841 3417 14875 3451
rect 14875 3417 14884 3451
rect 14832 3408 14884 3417
rect 53288 3408 53340 3460
rect 57520 3519 57572 3528
rect 57520 3485 57529 3519
rect 57529 3485 57563 3519
rect 57563 3485 57572 3519
rect 57520 3476 57572 3485
rect 58164 3519 58216 3528
rect 58164 3485 58173 3519
rect 58173 3485 58207 3519
rect 58207 3485 58216 3519
rect 58164 3476 58216 3485
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 5724 3136 5776 3188
rect 5908 3136 5960 3188
rect 7564 3136 7616 3188
rect 7840 3136 7892 3188
rect 3332 3111 3384 3120
rect 3332 3077 3366 3111
rect 3366 3077 3384 3111
rect 3332 3068 3384 3077
rect 5080 3068 5132 3120
rect 7104 3068 7156 3120
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 4988 3000 5040 3052
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 5908 3000 5960 3052
rect 6276 3000 6328 3052
rect 6828 3000 6880 3052
rect 7748 3000 7800 3052
rect 2136 2932 2188 2984
rect 4804 2932 4856 2984
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 5724 2864 5776 2916
rect 5816 2864 5868 2916
rect 8760 3068 8812 3120
rect 9404 3068 9456 3120
rect 10416 3111 10468 3120
rect 10416 3077 10425 3111
rect 10425 3077 10459 3111
rect 10459 3077 10468 3111
rect 10416 3068 10468 3077
rect 12072 3136 12124 3188
rect 10968 3068 11020 3120
rect 14280 3136 14332 3188
rect 26240 3068 26292 3120
rect 51908 3068 51960 3120
rect 8576 3000 8628 3052
rect 8852 3000 8904 3052
rect 9496 3000 9548 3052
rect 12624 3000 12676 3052
rect 13452 3000 13504 3052
rect 14464 3000 14516 3052
rect 51724 3000 51776 3052
rect 54760 3000 54812 3052
rect 4712 2796 4764 2848
rect 4988 2796 5040 2848
rect 5080 2839 5132 2848
rect 5080 2805 5089 2839
rect 5089 2805 5123 2839
rect 5123 2805 5132 2839
rect 5080 2796 5132 2805
rect 8024 2796 8076 2848
rect 9128 2932 9180 2984
rect 9312 2932 9364 2984
rect 11704 2932 11756 2984
rect 18696 2932 18748 2984
rect 19984 2932 20036 2984
rect 26424 2932 26476 2984
rect 32772 2932 32824 2984
rect 38292 2932 38344 2984
rect 42156 2932 42208 2984
rect 53104 2932 53156 2984
rect 56600 2975 56652 2984
rect 56600 2941 56609 2975
rect 56609 2941 56643 2975
rect 56643 2941 56652 2975
rect 56600 2932 56652 2941
rect 8852 2864 8904 2916
rect 14924 2864 14976 2916
rect 33876 2864 33928 2916
rect 37188 2864 37240 2916
rect 39120 2864 39172 2916
rect 40224 2864 40276 2916
rect 42984 2864 43036 2916
rect 44088 2864 44140 2916
rect 8668 2796 8720 2848
rect 14648 2796 14700 2848
rect 15384 2796 15436 2848
rect 15660 2796 15712 2848
rect 16488 2796 16540 2848
rect 17868 2796 17920 2848
rect 19248 2796 19300 2848
rect 20536 2796 20588 2848
rect 20904 2796 20956 2848
rect 21732 2796 21784 2848
rect 23112 2796 23164 2848
rect 23664 2796 23716 2848
rect 24216 2796 24268 2848
rect 25044 2796 25096 2848
rect 25872 2796 25924 2848
rect 26976 2796 27028 2848
rect 27804 2796 27856 2848
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 29184 2796 29236 2848
rect 29736 2796 29788 2848
rect 30012 2839 30064 2848
rect 30012 2805 30021 2839
rect 30021 2805 30055 2839
rect 30055 2805 30064 2839
rect 30012 2796 30064 2805
rect 30564 2796 30616 2848
rect 31668 2796 31720 2848
rect 32220 2796 32272 2848
rect 33324 2796 33376 2848
rect 34428 2796 34480 2848
rect 35440 2796 35492 2848
rect 36360 2796 36412 2848
rect 37740 2796 37792 2848
rect 39672 2796 39724 2848
rect 41604 2796 41656 2848
rect 43536 2796 43588 2848
rect 44916 2796 44968 2848
rect 47400 2864 47452 2916
rect 48780 2864 48832 2916
rect 49884 2864 49936 2916
rect 50988 2864 51040 2916
rect 54208 2864 54260 2916
rect 45468 2796 45520 2848
rect 46848 2796 46900 2848
rect 47952 2796 48004 2848
rect 49332 2796 49384 2848
rect 50712 2796 50764 2848
rect 51540 2796 51592 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 2780 2592 2832 2644
rect 5908 2592 5960 2644
rect 6644 2635 6696 2644
rect 6644 2601 6653 2635
rect 6653 2601 6687 2635
rect 6687 2601 6696 2635
rect 6644 2592 6696 2601
rect 8576 2592 8628 2644
rect 13912 2592 13964 2644
rect 5264 2524 5316 2576
rect 3792 2456 3844 2508
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 2228 2388 2280 2440
rect 2872 2388 2924 2440
rect 4068 2388 4120 2440
rect 4988 2456 5040 2508
rect 9404 2524 9456 2576
rect 9680 2524 9732 2576
rect 11520 2524 11572 2576
rect 5632 2388 5684 2440
rect 6092 2388 6144 2440
rect 7196 2388 7248 2440
rect 7472 2456 7524 2508
rect 9496 2456 9548 2508
rect 16212 2524 16264 2576
rect 21456 2592 21508 2644
rect 52000 2592 52052 2644
rect 27436 2524 27488 2576
rect 28356 2524 28408 2576
rect 34152 2524 34204 2576
rect 38016 2524 38068 2576
rect 41880 2524 41932 2576
rect 45744 2524 45796 2576
rect 49608 2524 49660 2576
rect 9404 2388 9456 2440
rect 5908 2252 5960 2304
rect 7932 2320 7984 2372
rect 8208 2320 8260 2372
rect 9496 2320 9548 2372
rect 9588 2320 9640 2372
rect 11704 2388 11756 2440
rect 12256 2431 12308 2440
rect 12256 2397 12265 2431
rect 12265 2397 12299 2431
rect 12299 2397 12308 2431
rect 12256 2388 12308 2397
rect 17040 2456 17092 2508
rect 18144 2456 18196 2508
rect 20076 2456 20128 2508
rect 22008 2456 22060 2508
rect 25320 2456 25372 2508
rect 26700 2456 26752 2508
rect 31944 2456 31996 2508
rect 33048 2456 33100 2508
rect 35532 2456 35584 2508
rect 38844 2456 38896 2508
rect 40776 2456 40828 2508
rect 43260 2456 43312 2508
rect 46572 2456 46624 2508
rect 48504 2456 48556 2508
rect 17316 2388 17368 2440
rect 15016 2320 15068 2372
rect 7380 2252 7432 2304
rect 9404 2252 9456 2304
rect 9864 2295 9916 2304
rect 9864 2261 9873 2295
rect 9873 2261 9907 2295
rect 9907 2261 9916 2295
rect 9864 2252 9916 2261
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 18972 2320 19024 2372
rect 22836 2320 22888 2372
rect 24768 2388 24820 2440
rect 26148 2388 26200 2440
rect 27252 2388 27304 2440
rect 28908 2388 28960 2440
rect 29460 2388 29512 2440
rect 30288 2388 30340 2440
rect 30840 2388 30892 2440
rect 31116 2388 31168 2440
rect 31392 2388 31444 2440
rect 32496 2388 32548 2440
rect 33600 2388 33652 2440
rect 36084 2388 36136 2440
rect 23940 2320 23992 2372
rect 36912 2320 36964 2372
rect 39396 2388 39448 2440
rect 41328 2388 41380 2440
rect 43812 2388 43864 2440
rect 44640 2320 44692 2372
rect 47124 2388 47176 2440
rect 49056 2388 49108 2440
rect 50896 2388 50948 2440
rect 57888 2499 57940 2508
rect 52552 2388 52604 2440
rect 51264 2252 51316 2304
rect 57888 2465 57897 2499
rect 57897 2465 57931 2499
rect 57931 2465 57940 2499
rect 57888 2456 57940 2465
rect 55956 2431 56008 2440
rect 55956 2397 55965 2431
rect 55965 2397 55999 2431
rect 55999 2397 56008 2431
rect 55956 2388 56008 2397
rect 56600 2431 56652 2440
rect 56600 2397 56609 2431
rect 56609 2397 56643 2431
rect 56643 2397 56652 2431
rect 56600 2388 56652 2397
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 5264 2048 5316 2100
rect 6644 2048 6696 2100
rect 52368 2048 52420 2100
rect 55956 2048 56008 2100
rect 11520 1980 11572 2032
rect 17224 1980 17276 2032
rect 53564 1980 53616 2032
rect 57888 1980 57940 2032
rect 12348 1912 12400 1964
rect 20168 1912 20220 1964
rect 1584 1844 1636 1896
rect 7472 1844 7524 1896
rect 7932 1708 7984 1760
rect 8208 1708 8260 1760
rect 5908 1504 5960 1556
rect 7748 1504 7800 1556
rect 3056 1368 3108 1420
rect 5908 1368 5960 1420
rect 7472 1368 7524 1420
rect 52736 1368 52788 1420
rect 53012 1368 53064 1420
rect 5356 1300 5408 1352
rect 6000 1300 6052 1352
rect 7840 1300 7892 1352
rect 52552 1096 52604 1148
rect 50988 892 51040 944
rect 52552 892 52604 944
rect 52920 892 52972 944
rect 56600 1368 56652 1420
rect 54760 824 54812 876
<< metal2 >>
rect 1766 59200 1822 60000
rect 3330 59200 3386 60000
rect 4894 59200 4950 60000
rect 6458 59200 6514 60000
rect 8022 59200 8078 60000
rect 9586 59200 9642 60000
rect 11150 59200 11206 60000
rect 12714 59200 12770 60000
rect 14278 59200 14334 60000
rect 15842 59200 15898 60000
rect 17406 59200 17462 60000
rect 18970 59200 19026 60000
rect 20534 59200 20590 60000
rect 22098 59200 22154 60000
rect 23662 59200 23718 60000
rect 25226 59200 25282 60000
rect 26790 59200 26846 60000
rect 28354 59200 28410 60000
rect 29918 59200 29974 60000
rect 31482 59200 31538 60000
rect 33046 59200 33102 60000
rect 34610 59200 34666 60000
rect 36174 59200 36230 60000
rect 37738 59200 37794 60000
rect 39302 59200 39358 60000
rect 40866 59200 40922 60000
rect 42430 59200 42486 60000
rect 43994 59200 44050 60000
rect 45558 59200 45614 60000
rect 47122 59200 47178 60000
rect 48686 59200 48742 60000
rect 50250 59200 50306 60000
rect 51814 59200 51870 60000
rect 53378 59200 53434 60000
rect 54942 59200 54998 60000
rect 56506 59200 56562 60000
rect 58070 59200 58126 60000
rect 58438 59256 58494 59265
rect 1780 57458 1808 59200
rect 3344 57458 3372 59200
rect 4908 57458 4936 59200
rect 6472 57458 6500 59200
rect 8036 57458 8064 59200
rect 1768 57452 1820 57458
rect 1768 57394 1820 57400
rect 3332 57452 3384 57458
rect 3332 57394 3384 57400
rect 4896 57452 4948 57458
rect 4896 57394 4948 57400
rect 6460 57452 6512 57458
rect 6460 57394 6512 57400
rect 8024 57452 8076 57458
rect 9600 57440 9628 59200
rect 11164 57458 11192 59200
rect 12728 57458 12756 59200
rect 14292 57458 14320 59200
rect 15856 57458 15884 59200
rect 17420 57458 17448 59200
rect 18984 57458 19012 59200
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 20548 57458 20576 59200
rect 22112 57458 22140 59200
rect 23676 57458 23704 59200
rect 25240 57458 25268 59200
rect 26804 57458 26832 59200
rect 28368 57458 28396 59200
rect 29932 57458 29960 59200
rect 31496 57458 31524 59200
rect 9680 57452 9732 57458
rect 9600 57412 9680 57440
rect 8024 57394 8076 57400
rect 9680 57394 9732 57400
rect 11152 57452 11204 57458
rect 11152 57394 11204 57400
rect 12716 57452 12768 57458
rect 12716 57394 12768 57400
rect 14280 57452 14332 57458
rect 14280 57394 14332 57400
rect 15844 57452 15896 57458
rect 15844 57394 15896 57400
rect 17408 57452 17460 57458
rect 17408 57394 17460 57400
rect 18972 57452 19024 57458
rect 18972 57394 19024 57400
rect 20536 57452 20588 57458
rect 20536 57394 20588 57400
rect 22100 57452 22152 57458
rect 22100 57394 22152 57400
rect 23664 57452 23716 57458
rect 23664 57394 23716 57400
rect 25228 57452 25280 57458
rect 25228 57394 25280 57400
rect 26792 57452 26844 57458
rect 26792 57394 26844 57400
rect 28356 57452 28408 57458
rect 28356 57394 28408 57400
rect 29920 57452 29972 57458
rect 29920 57394 29972 57400
rect 31484 57452 31536 57458
rect 33060 57440 33088 59200
rect 34624 57458 34652 59200
rect 36188 57458 36216 59200
rect 37752 57458 37780 59200
rect 39316 57458 39344 59200
rect 40880 57458 40908 59200
rect 42444 57458 42472 59200
rect 44008 57458 44036 59200
rect 45572 57458 45600 59200
rect 47136 57458 47164 59200
rect 48700 57458 48728 59200
rect 50264 57882 50292 59200
rect 50172 57854 50292 57882
rect 50172 57458 50200 57854
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 51828 57458 51856 59200
rect 53392 57458 53420 59200
rect 33140 57452 33192 57458
rect 33060 57412 33140 57440
rect 31484 57394 31536 57400
rect 33140 57394 33192 57400
rect 34612 57452 34664 57458
rect 34612 57394 34664 57400
rect 36176 57452 36228 57458
rect 36176 57394 36228 57400
rect 37740 57452 37792 57458
rect 37740 57394 37792 57400
rect 39304 57452 39356 57458
rect 39304 57394 39356 57400
rect 40868 57452 40920 57458
rect 40868 57394 40920 57400
rect 42432 57452 42484 57458
rect 42432 57394 42484 57400
rect 43996 57452 44048 57458
rect 43996 57394 44048 57400
rect 45560 57452 45612 57458
rect 45560 57394 45612 57400
rect 47124 57452 47176 57458
rect 47124 57394 47176 57400
rect 48688 57452 48740 57458
rect 48688 57394 48740 57400
rect 50160 57452 50212 57458
rect 50160 57394 50212 57400
rect 51816 57452 51868 57458
rect 51816 57394 51868 57400
rect 53380 57452 53432 57458
rect 53380 57394 53432 57400
rect 54956 57390 54984 59200
rect 56520 57882 56548 59200
rect 57518 57896 57574 57905
rect 56520 57854 56640 57882
rect 56612 57458 56640 57854
rect 57518 57831 57574 57840
rect 56600 57452 56652 57458
rect 56600 57394 56652 57400
rect 54944 57384 54996 57390
rect 54944 57326 54996 57332
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 57532 57050 57560 57831
rect 58084 57458 58112 59200
rect 58438 59191 58494 59200
rect 58072 57452 58124 57458
rect 58072 57394 58124 57400
rect 57520 57044 57572 57050
rect 57520 56986 57572 56992
rect 57888 56840 57940 56846
rect 57888 56782 57940 56788
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 57900 56545 57928 56782
rect 57886 56536 57942 56545
rect 57886 56471 57942 56480
rect 58452 56370 58480 59191
rect 58440 56364 58492 56370
rect 58440 56306 58492 56312
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 58162 55176 58218 55185
rect 58162 55111 58164 55120
rect 58216 55111 58218 55120
rect 58164 55082 58216 55088
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 57888 53984 57940 53990
rect 57888 53926 57940 53932
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 57900 53825 57928 53926
rect 57886 53816 57942 53825
rect 57886 53751 57942 53760
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 57888 52488 57940 52494
rect 57886 52456 57888 52465
rect 57940 52456 57942 52465
rect 57886 52391 57942 52400
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 58164 51400 58216 51406
rect 58164 51342 58216 51348
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 58176 51105 58204 51342
rect 58162 51096 58218 51105
rect 58162 51031 58218 51040
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 58164 49768 58216 49774
rect 58162 49736 58164 49745
rect 58216 49736 58218 49745
rect 58162 49671 58218 49680
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 58164 48544 58216 48550
rect 58164 48486 58216 48492
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 58176 48385 58204 48486
rect 58162 48376 58218 48385
rect 58162 48311 58218 48320
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 58164 47048 58216 47054
rect 58162 47016 58164 47025
rect 58216 47016 58218 47025
rect 58162 46951 58218 46960
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 58164 45960 58216 45966
rect 58164 45902 58216 45908
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 58176 45665 58204 45902
rect 58162 45656 58218 45665
rect 58162 45591 58218 45600
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 58162 44296 58218 44305
rect 58162 44231 58164 44240
rect 58216 44231 58218 44240
rect 58164 44202 58216 44208
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 58164 43104 58216 43110
rect 58164 43046 58216 43052
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 58176 42945 58204 43046
rect 58162 42936 58218 42945
rect 58162 42871 58218 42880
rect 12716 42696 12768 42702
rect 12716 42638 12768 42644
rect 20444 42696 20496 42702
rect 20444 42638 20496 42644
rect 12164 42356 12216 42362
rect 12164 42298 12216 42304
rect 12072 42016 12124 42022
rect 12072 41958 12124 41964
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 12084 41614 12112 41958
rect 12072 41608 12124 41614
rect 12072 41550 12124 41556
rect 11244 41540 11296 41546
rect 11244 41482 11296 41488
rect 11428 41540 11480 41546
rect 11428 41482 11480 41488
rect 5172 41472 5224 41478
rect 5172 41414 5224 41420
rect 4620 40928 4672 40934
rect 4620 40870 4672 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4632 40526 4660 40870
rect 5184 40526 5212 41414
rect 11256 41206 11284 41482
rect 11440 41414 11468 41482
rect 11440 41386 11560 41414
rect 6368 41200 6420 41206
rect 6368 41142 6420 41148
rect 11244 41200 11296 41206
rect 11244 41142 11296 41148
rect 6000 41132 6052 41138
rect 6000 41074 6052 41080
rect 4436 40520 4488 40526
rect 4436 40462 4488 40468
rect 4620 40520 4672 40526
rect 4620 40462 4672 40468
rect 4712 40520 4764 40526
rect 4712 40462 4764 40468
rect 5172 40520 5224 40526
rect 5172 40462 5224 40468
rect 2412 40044 2464 40050
rect 2412 39986 2464 39992
rect 2424 39642 2452 39986
rect 4448 39982 4476 40462
rect 4068 39976 4120 39982
rect 4068 39918 4120 39924
rect 4436 39976 4488 39982
rect 4436 39918 4488 39924
rect 3240 39908 3292 39914
rect 3240 39850 3292 39856
rect 2780 39840 2832 39846
rect 2780 39782 2832 39788
rect 2412 39636 2464 39642
rect 2412 39578 2464 39584
rect 2596 39364 2648 39370
rect 2596 39306 2648 39312
rect 2608 38010 2636 39306
rect 2596 38004 2648 38010
rect 2596 37946 2648 37952
rect 2320 37664 2372 37670
rect 2320 37606 2372 37612
rect 2332 37194 2360 37606
rect 2608 37466 2636 37946
rect 2792 37738 2820 39782
rect 3252 39438 3280 39850
rect 3976 39840 4028 39846
rect 3976 39782 4028 39788
rect 2872 39432 2924 39438
rect 2872 39374 2924 39380
rect 3240 39432 3292 39438
rect 3240 39374 3292 39380
rect 3792 39432 3844 39438
rect 3792 39374 3844 39380
rect 2884 38758 2912 39374
rect 2872 38752 2924 38758
rect 2872 38694 2924 38700
rect 3148 38208 3200 38214
rect 3148 38150 3200 38156
rect 2872 37868 2924 37874
rect 2872 37810 2924 37816
rect 2780 37732 2832 37738
rect 2780 37674 2832 37680
rect 2596 37460 2648 37466
rect 2596 37402 2648 37408
rect 2792 37194 2820 37674
rect 2320 37188 2372 37194
rect 2320 37130 2372 37136
rect 2780 37188 2832 37194
rect 2780 37130 2832 37136
rect 2792 35630 2820 37130
rect 2884 36922 2912 37810
rect 3160 37806 3188 38150
rect 3252 37874 3280 39374
rect 3804 38350 3832 39374
rect 3988 39370 4016 39782
rect 3976 39364 4028 39370
rect 3976 39306 4028 39312
rect 3792 38344 3844 38350
rect 3792 38286 3844 38292
rect 3240 37868 3292 37874
rect 3240 37810 3292 37816
rect 3804 37806 3832 38286
rect 3884 38276 3936 38282
rect 3884 38218 3936 38224
rect 3148 37800 3200 37806
rect 3148 37742 3200 37748
rect 3792 37800 3844 37806
rect 3792 37742 3844 37748
rect 3056 37120 3108 37126
rect 3056 37062 3108 37068
rect 2872 36916 2924 36922
rect 2872 36858 2924 36864
rect 3068 36786 3096 37062
rect 3056 36780 3108 36786
rect 3056 36722 3108 36728
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2792 34746 2820 35566
rect 2780 34740 2832 34746
rect 2780 34682 2832 34688
rect 2136 32360 2188 32366
rect 2136 32302 2188 32308
rect 1952 31816 2004 31822
rect 2148 31770 2176 32302
rect 2004 31764 2176 31770
rect 1952 31758 2176 31764
rect 1964 31742 2176 31758
rect 3068 31754 3096 36722
rect 3160 33998 3188 37742
rect 3804 37126 3832 37742
rect 3896 37466 3924 38218
rect 3884 37460 3936 37466
rect 3884 37402 3936 37408
rect 3792 37120 3844 37126
rect 3792 37062 3844 37068
rect 3792 34604 3844 34610
rect 3792 34546 3844 34552
rect 3804 34202 3832 34546
rect 3792 34196 3844 34202
rect 3792 34138 3844 34144
rect 3424 34060 3476 34066
rect 3424 34002 3476 34008
rect 3148 33992 3200 33998
rect 3148 33934 3200 33940
rect 3332 33856 3384 33862
rect 3332 33798 3384 33804
rect 2148 31346 2176 31742
rect 2596 31748 2648 31754
rect 3068 31726 3188 31754
rect 2596 31690 2648 31696
rect 2136 31340 2188 31346
rect 2136 31282 2188 31288
rect 2608 30938 2636 31690
rect 2964 31476 3016 31482
rect 2964 31418 3016 31424
rect 2688 31340 2740 31346
rect 2688 31282 2740 31288
rect 2596 30932 2648 30938
rect 2596 30874 2648 30880
rect 2700 30394 2728 31282
rect 2976 30598 3004 31418
rect 2964 30592 3016 30598
rect 2964 30534 3016 30540
rect 2976 30394 3004 30534
rect 2688 30388 2740 30394
rect 2688 30330 2740 30336
rect 2964 30388 3016 30394
rect 2964 30330 3016 30336
rect 2780 29640 2832 29646
rect 2780 29582 2832 29588
rect 2792 28558 2820 29582
rect 2780 28552 2832 28558
rect 2780 28494 2832 28500
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2320 28008 2372 28014
rect 2320 27950 2372 27956
rect 2332 25906 2360 27950
rect 2608 27674 2636 28018
rect 2596 27668 2648 27674
rect 2596 27610 2648 27616
rect 2976 27334 3004 30330
rect 3160 29714 3188 31726
rect 3344 30734 3372 33798
rect 3436 31482 3464 34002
rect 3792 32768 3844 32774
rect 3792 32710 3844 32716
rect 3804 32434 3832 32710
rect 3792 32428 3844 32434
rect 3792 32370 3844 32376
rect 3884 31680 3936 31686
rect 3884 31622 3936 31628
rect 3424 31476 3476 31482
rect 3424 31418 3476 31424
rect 3792 31476 3844 31482
rect 3792 31418 3844 31424
rect 3516 31136 3568 31142
rect 3516 31078 3568 31084
rect 3332 30728 3384 30734
rect 3332 30670 3384 30676
rect 3240 30388 3292 30394
rect 3240 30330 3292 30336
rect 3252 29850 3280 30330
rect 3344 30258 3372 30670
rect 3332 30252 3384 30258
rect 3332 30194 3384 30200
rect 3240 29844 3292 29850
rect 3240 29786 3292 29792
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 3148 28416 3200 28422
rect 3148 28358 3200 28364
rect 3160 27402 3188 28358
rect 3344 27470 3372 30194
rect 3424 30116 3476 30122
rect 3424 30058 3476 30064
rect 3332 27464 3384 27470
rect 3332 27406 3384 27412
rect 3148 27396 3200 27402
rect 3148 27338 3200 27344
rect 2964 27328 3016 27334
rect 2964 27270 3016 27276
rect 3436 26994 3464 30058
rect 3528 29646 3556 31078
rect 3516 29640 3568 29646
rect 3516 29582 3568 29588
rect 3700 28552 3752 28558
rect 3700 28494 3752 28500
rect 3712 28218 3740 28494
rect 3700 28212 3752 28218
rect 3700 28154 3752 28160
rect 3608 27328 3660 27334
rect 3608 27270 3660 27276
rect 3516 27124 3568 27130
rect 3516 27066 3568 27072
rect 2688 26988 2740 26994
rect 2688 26930 2740 26936
rect 3424 26988 3476 26994
rect 3424 26930 3476 26936
rect 2700 26790 2728 26930
rect 2688 26784 2740 26790
rect 2688 26726 2740 26732
rect 3148 26784 3200 26790
rect 3148 26726 3200 26732
rect 2596 26376 2648 26382
rect 2596 26318 2648 26324
rect 2320 25900 2372 25906
rect 2320 25842 2372 25848
rect 2332 24886 2360 25842
rect 2608 24954 2636 26318
rect 2596 24948 2648 24954
rect 2596 24890 2648 24896
rect 2320 24880 2372 24886
rect 2320 24822 2372 24828
rect 1860 23724 1912 23730
rect 1860 23666 1912 23672
rect 1872 21894 1900 23666
rect 2700 23254 2728 26726
rect 3160 25974 3188 26726
rect 3528 26246 3556 27066
rect 3620 26994 3648 27270
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 3700 26920 3752 26926
rect 3700 26862 3752 26868
rect 3712 26450 3740 26862
rect 3700 26444 3752 26450
rect 3700 26386 3752 26392
rect 3700 26308 3752 26314
rect 3700 26250 3752 26256
rect 3516 26240 3568 26246
rect 3516 26182 3568 26188
rect 3148 25968 3200 25974
rect 3148 25910 3200 25916
rect 3712 24818 3740 26250
rect 3804 25430 3832 31418
rect 3896 30734 3924 31622
rect 3884 30728 3936 30734
rect 3884 30670 3936 30676
rect 3896 30258 3924 30670
rect 3988 30326 4016 39306
rect 4080 39098 4108 39918
rect 4724 39914 4752 40462
rect 5080 40384 5132 40390
rect 5080 40326 5132 40332
rect 4712 39908 4764 39914
rect 4712 39850 4764 39856
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4724 39506 4752 39850
rect 4712 39500 4764 39506
rect 4712 39442 4764 39448
rect 5092 39438 5120 40326
rect 5080 39432 5132 39438
rect 5080 39374 5132 39380
rect 4068 39092 4120 39098
rect 4068 39034 4120 39040
rect 4712 38752 4764 38758
rect 4712 38694 4764 38700
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4620 37868 4672 37874
rect 4620 37810 4672 37816
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37448 4660 37810
rect 4448 37420 4660 37448
rect 4448 37262 4476 37420
rect 4724 37346 4752 38694
rect 4632 37318 4752 37346
rect 4436 37256 4488 37262
rect 4436 37198 4488 37204
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 35692 4120 35698
rect 4068 35634 4120 35640
rect 4080 34746 4108 35634
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 34740 4120 34746
rect 4068 34682 4120 34688
rect 4632 34610 4660 37318
rect 4988 37188 5040 37194
rect 4988 37130 5040 37136
rect 5000 36038 5028 37130
rect 4988 36032 5040 36038
rect 4988 35974 5040 35980
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4724 35018 4752 35430
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4804 34944 4856 34950
rect 4804 34886 4856 34892
rect 5080 34944 5132 34950
rect 5080 34886 5132 34892
rect 4816 34610 4844 34886
rect 5092 34610 5120 34886
rect 4620 34604 4672 34610
rect 4620 34546 4672 34552
rect 4804 34604 4856 34610
rect 4804 34546 4856 34552
rect 5080 34604 5132 34610
rect 5080 34546 5132 34552
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 33992 4120 33998
rect 4068 33934 4120 33940
rect 4252 33992 4304 33998
rect 4252 33934 4304 33940
rect 4080 31482 4108 33934
rect 4264 33658 4292 33934
rect 4252 33652 4304 33658
rect 4252 33594 4304 33600
rect 4632 33425 4660 34546
rect 4896 34536 4948 34542
rect 4896 34478 4948 34484
rect 4908 33930 4936 34478
rect 5092 34406 5120 34546
rect 4988 34400 5040 34406
rect 4988 34342 5040 34348
rect 5080 34400 5132 34406
rect 5080 34342 5132 34348
rect 4896 33924 4948 33930
rect 4896 33866 4948 33872
rect 4908 33658 4936 33866
rect 4896 33652 4948 33658
rect 4896 33594 4948 33600
rect 4712 33584 4764 33590
rect 4908 33538 4936 33594
rect 5000 33590 5028 34342
rect 5092 33998 5120 34342
rect 5080 33992 5132 33998
rect 5080 33934 5132 33940
rect 4712 33526 4764 33532
rect 4618 33416 4674 33425
rect 4618 33351 4674 33360
rect 4620 33312 4672 33318
rect 4620 33254 4672 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4632 32978 4660 33254
rect 4620 32972 4672 32978
rect 4620 32914 4672 32920
rect 4724 32298 4752 33526
rect 4816 33510 4936 33538
rect 4988 33584 5040 33590
rect 4988 33526 5040 33532
rect 4816 33046 4844 33510
rect 5000 33454 5028 33526
rect 4988 33448 5040 33454
rect 4988 33390 5040 33396
rect 4896 33312 4948 33318
rect 4896 33254 4948 33260
rect 4986 33280 5042 33289
rect 4804 33040 4856 33046
rect 4804 32982 4856 32988
rect 4712 32292 4764 32298
rect 4712 32234 4764 32240
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4068 31476 4120 31482
rect 4068 31418 4120 31424
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30870 4108 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4068 30864 4120 30870
rect 4068 30806 4120 30812
rect 3976 30320 4028 30326
rect 3976 30262 4028 30268
rect 3884 30252 3936 30258
rect 3884 30194 3936 30200
rect 3884 27464 3936 27470
rect 3884 27406 3936 27412
rect 3896 26586 3924 27406
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3884 26580 3936 26586
rect 3884 26522 3936 26528
rect 3896 26382 3924 26522
rect 3884 26376 3936 26382
rect 3884 26318 3936 26324
rect 3988 26042 4016 27338
rect 4080 26382 4108 30806
rect 4620 30728 4672 30734
rect 4620 30670 4672 30676
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29782 4660 30670
rect 4804 30048 4856 30054
rect 4804 29990 4856 29996
rect 4620 29776 4672 29782
rect 4620 29718 4672 29724
rect 4712 29504 4764 29510
rect 4712 29446 4764 29452
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4620 27872 4672 27878
rect 4620 27814 4672 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27538 4660 27814
rect 4620 27532 4672 27538
rect 4620 27474 4672 27480
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4068 26376 4120 26382
rect 4068 26318 4120 26324
rect 4080 26042 4108 26318
rect 4632 26314 4660 27474
rect 4724 27470 4752 29446
rect 4712 27464 4764 27470
rect 4712 27406 4764 27412
rect 4816 26994 4844 29990
rect 4908 27606 4936 33254
rect 4986 33215 5042 33224
rect 5000 30376 5028 33215
rect 5092 32978 5120 33934
rect 5080 32972 5132 32978
rect 5080 32914 5132 32920
rect 5184 32842 5212 40462
rect 5540 40384 5592 40390
rect 5540 40326 5592 40332
rect 5552 40118 5580 40326
rect 6012 40186 6040 41074
rect 6000 40180 6052 40186
rect 6000 40122 6052 40128
rect 5540 40112 5592 40118
rect 5540 40054 5592 40060
rect 6012 39370 6040 40122
rect 6380 39642 6408 41142
rect 9312 41132 9364 41138
rect 9312 41074 9364 41080
rect 10140 41132 10192 41138
rect 10140 41074 10192 41080
rect 6920 40928 6972 40934
rect 6920 40870 6972 40876
rect 8116 40928 8168 40934
rect 8116 40870 8168 40876
rect 6932 40526 6960 40870
rect 6920 40520 6972 40526
rect 6920 40462 6972 40468
rect 8128 40458 8156 40870
rect 9324 40730 9352 41074
rect 9956 41064 10008 41070
rect 9956 41006 10008 41012
rect 9312 40724 9364 40730
rect 9312 40666 9364 40672
rect 8484 40520 8536 40526
rect 8484 40462 8536 40468
rect 7012 40452 7064 40458
rect 7012 40394 7064 40400
rect 8116 40452 8168 40458
rect 8116 40394 8168 40400
rect 7024 39982 7052 40394
rect 8496 40050 8524 40462
rect 9036 40452 9088 40458
rect 9036 40394 9088 40400
rect 9048 40118 9076 40394
rect 9864 40384 9916 40390
rect 9864 40326 9916 40332
rect 9772 40180 9824 40186
rect 9772 40122 9824 40128
rect 8576 40112 8628 40118
rect 8576 40054 8628 40060
rect 9036 40112 9088 40118
rect 9036 40054 9088 40060
rect 7104 40044 7156 40050
rect 7104 39986 7156 39992
rect 8484 40044 8536 40050
rect 8484 39986 8536 39992
rect 7012 39976 7064 39982
rect 7012 39918 7064 39924
rect 6644 39908 6696 39914
rect 6644 39850 6696 39856
rect 6368 39636 6420 39642
rect 6368 39578 6420 39584
rect 6000 39364 6052 39370
rect 6000 39306 6052 39312
rect 5724 38956 5776 38962
rect 5724 38898 5776 38904
rect 5264 38208 5316 38214
rect 5264 38150 5316 38156
rect 5540 38208 5592 38214
rect 5540 38150 5592 38156
rect 5276 36768 5304 38150
rect 5356 37256 5408 37262
rect 5552 37244 5580 38150
rect 5736 37874 5764 38898
rect 6012 38282 6040 39306
rect 6000 38276 6052 38282
rect 6000 38218 6052 38224
rect 5724 37868 5776 37874
rect 5724 37810 5776 37816
rect 5736 37670 5764 37810
rect 5724 37664 5776 37670
rect 5724 37606 5776 37612
rect 5408 37216 5580 37244
rect 5356 37198 5408 37204
rect 5632 37120 5684 37126
rect 5632 37062 5684 37068
rect 5276 36740 5396 36768
rect 5264 35012 5316 35018
rect 5264 34954 5316 34960
rect 5172 32836 5224 32842
rect 5172 32778 5224 32784
rect 5184 32570 5212 32778
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5000 30348 5212 30376
rect 5080 30252 5132 30258
rect 5080 30194 5132 30200
rect 4988 30184 5040 30190
rect 4988 30126 5040 30132
rect 5000 29578 5028 30126
rect 5092 29646 5120 30194
rect 5080 29640 5132 29646
rect 5080 29582 5132 29588
rect 4988 29572 5040 29578
rect 4988 29514 5040 29520
rect 5000 28626 5028 29514
rect 4988 28620 5040 28626
rect 4988 28562 5040 28568
rect 5092 28558 5120 29582
rect 5080 28552 5132 28558
rect 5080 28494 5132 28500
rect 4896 27600 4948 27606
rect 4896 27542 4948 27548
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 4896 27328 4948 27334
rect 4896 27270 4948 27276
rect 4908 27130 4936 27270
rect 5000 27130 5028 27406
rect 5080 27328 5132 27334
rect 5080 27270 5132 27276
rect 4896 27124 4948 27130
rect 4896 27066 4948 27072
rect 4988 27124 5040 27130
rect 4988 27066 5040 27072
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4908 26382 4936 27066
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 3792 25424 3844 25430
rect 3792 25366 3844 25372
rect 3700 24812 3752 24818
rect 3700 24754 3752 24760
rect 3792 23792 3844 23798
rect 3792 23734 3844 23740
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3332 23588 3384 23594
rect 3332 23530 3384 23536
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2688 23248 2740 23254
rect 2688 23190 2740 23196
rect 3160 23050 3188 23462
rect 3148 23044 3200 23050
rect 3148 22986 3200 22992
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 1860 21888 1912 21894
rect 1860 21830 1912 21836
rect 1872 21078 1900 21830
rect 2700 21554 2728 22918
rect 3344 22642 3372 23530
rect 3332 22636 3384 22642
rect 3332 22578 3384 22584
rect 2964 22432 3016 22438
rect 2964 22374 3016 22380
rect 2976 22030 3004 22374
rect 2964 22024 3016 22030
rect 2964 21966 3016 21972
rect 3436 21894 3464 23666
rect 3608 23180 3660 23186
rect 3608 23122 3660 23128
rect 3516 23112 3568 23118
rect 3516 23054 3568 23060
rect 3528 22642 3556 23054
rect 3620 22710 3648 23122
rect 3608 22704 3660 22710
rect 3608 22646 3660 22652
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3424 21888 3476 21894
rect 3424 21830 3476 21836
rect 3712 21570 3740 22510
rect 3804 21962 3832 23734
rect 4080 22658 4108 25978
rect 4908 25974 4936 26318
rect 4988 26308 5040 26314
rect 4988 26250 5040 26256
rect 4896 25968 4948 25974
rect 4896 25910 4948 25916
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4712 23248 4764 23254
rect 4764 23208 4844 23236
rect 4712 23190 4764 23196
rect 3896 22630 4108 22658
rect 4712 22636 4764 22642
rect 3896 22574 3924 22630
rect 4712 22578 4764 22584
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 4068 22500 4120 22506
rect 4068 22442 4120 22448
rect 4080 22234 4108 22442
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22228 4120 22234
rect 4068 22170 4120 22176
rect 4252 22024 4304 22030
rect 4252 21966 4304 21972
rect 3792 21956 3844 21962
rect 3792 21898 3844 21904
rect 3976 21956 4028 21962
rect 3976 21898 4028 21904
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3896 21690 3924 21830
rect 3988 21690 4016 21898
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 3976 21684 4028 21690
rect 3976 21626 4028 21632
rect 2688 21548 2740 21554
rect 3712 21542 4016 21570
rect 4264 21554 4292 21966
rect 4632 21622 4660 22374
rect 4724 21894 4752 22578
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 2688 21490 2740 21496
rect 1860 21072 1912 21078
rect 1860 21014 1912 21020
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2148 18766 2176 19654
rect 2424 19514 2452 19790
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3896 19514 3924 19722
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3792 19372 3844 19378
rect 3792 19314 3844 19320
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 1860 18760 1912 18766
rect 1860 18702 1912 18708
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1872 18358 1900 18702
rect 1860 18352 1912 18358
rect 1860 18294 1912 18300
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17882 1808 18226
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 2608 17678 2636 19110
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2228 15904 2280 15910
rect 2228 15846 2280 15852
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 2148 14550 2176 15438
rect 2240 15026 2268 15846
rect 2516 15706 2544 16050
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2332 14618 2360 15438
rect 2792 15094 2820 18294
rect 2884 17746 2912 19246
rect 3804 18970 3832 19314
rect 3884 19236 3936 19242
rect 3884 19178 3936 19184
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3896 18850 3924 19178
rect 3804 18822 3924 18850
rect 3804 18086 3832 18822
rect 3792 18080 3844 18086
rect 3792 18022 3844 18028
rect 3804 17746 3832 18022
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 3792 17740 3844 17746
rect 3792 17682 3844 17688
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3896 16454 3924 17614
rect 3884 16448 3936 16454
rect 3884 16390 3936 16396
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 3424 15496 3476 15502
rect 3424 15438 3476 15444
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2148 12850 2176 14486
rect 2976 14482 3004 15098
rect 3068 14618 3096 15438
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 3436 14414 3464 15438
rect 3516 15360 3568 15366
rect 3516 15302 3568 15308
rect 3528 15026 3556 15302
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3896 14550 3924 16390
rect 3988 16046 4016 21542
rect 4252 21548 4304 21554
rect 4252 21490 4304 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4724 19854 4752 21830
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 4080 18970 4108 19246
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3988 15706 4016 15982
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 3884 14544 3936 14550
rect 3884 14486 3936 14492
rect 4080 14482 4108 18906
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4172 18426 4200 18566
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4264 18290 4292 18770
rect 4724 18698 4752 19110
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 18022
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4632 17202 4660 17818
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4724 17134 4752 18634
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 15162 4200 15438
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4632 15094 4660 15846
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3436 14074 3464 14350
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3436 13954 3464 14010
rect 3436 13926 3556 13954
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2240 11898 2268 12106
rect 2228 11892 2280 11898
rect 2228 11834 2280 11840
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1504 3754 1532 8298
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1596 7002 1624 7890
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1596 5302 1624 6938
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4146 1716 4966
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1504 3726 1624 3754
rect 1596 2446 1624 3726
rect 1780 3346 1808 8298
rect 2148 7410 2176 9454
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 4690 1992 7142
rect 2148 5914 2176 7346
rect 2332 6914 2360 12650
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 11762 2452 12582
rect 3436 12306 3464 12718
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3160 11898 3188 12174
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 3160 11694 3188 11834
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3252 11354 3280 11698
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10810 3096 11086
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2412 9920 2464 9926
rect 2412 9862 2464 9868
rect 2424 9654 2452 9862
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2608 9178 2636 9998
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7886 2820 8230
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 3252 7818 3280 8366
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 2872 7812 2924 7818
rect 2872 7754 2924 7760
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2700 7002 2728 7346
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2240 6886 2360 6914
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2148 5302 2176 5850
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1964 3534 1992 3878
rect 2148 3738 2176 5238
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1688 3318 1808 3346
rect 1688 3058 1716 3318
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1688 2961 1716 2994
rect 2148 2990 2176 3674
rect 2136 2984 2188 2990
rect 1674 2952 1730 2961
rect 2136 2926 2188 2932
rect 1674 2887 1730 2896
rect 2240 2446 2268 6886
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2424 6322 2452 6802
rect 2792 6798 2820 7686
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2884 6202 2912 7754
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2792 6174 2912 6202
rect 2410 5808 2466 5817
rect 2410 5743 2466 5752
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4146 2360 4422
rect 2424 4146 2452 5743
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2608 4214 2636 4558
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2792 3482 2820 6174
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 4146 2912 6054
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2976 4010 3004 5578
rect 3068 4622 3096 6598
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2792 3454 2912 3482
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2608 3058 2636 3334
rect 2778 3224 2834 3233
rect 2778 3159 2834 3168
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2792 2650 2820 3159
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 2884 2446 2912 3454
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 1596 1902 1624 2382
rect 1584 1896 1636 1902
rect 1584 1838 1636 1844
rect 3068 1426 3096 4558
rect 3344 3126 3372 7890
rect 3528 6186 3556 13926
rect 3620 12782 3648 14418
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 14074 4016 14350
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3896 9110 3924 12718
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12434 4752 17070
rect 4816 17066 4844 23208
rect 5000 22642 5028 26250
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 5092 22094 5120 27270
rect 5000 22066 5120 22094
rect 5184 22094 5212 30348
rect 5276 26858 5304 34954
rect 5368 28490 5396 36740
rect 5540 36032 5592 36038
rect 5540 35974 5592 35980
rect 5448 35012 5500 35018
rect 5448 34954 5500 34960
rect 5460 32366 5488 34954
rect 5552 32434 5580 35974
rect 5644 34202 5672 37062
rect 5632 34196 5684 34202
rect 5632 34138 5684 34144
rect 5540 32428 5592 32434
rect 5540 32370 5592 32376
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5460 30734 5488 32302
rect 5736 31822 5764 37606
rect 6012 36854 6040 38218
rect 6380 37942 6408 39578
rect 6656 38418 6684 39850
rect 6644 38412 6696 38418
rect 6644 38354 6696 38360
rect 6368 37936 6420 37942
rect 6368 37878 6420 37884
rect 6828 37868 6880 37874
rect 6828 37810 6880 37816
rect 6840 37126 6868 37810
rect 6184 37120 6236 37126
rect 6184 37062 6236 37068
rect 6828 37120 6880 37126
rect 6828 37062 6880 37068
rect 6000 36848 6052 36854
rect 6000 36790 6052 36796
rect 6092 36168 6144 36174
rect 6092 36110 6144 36116
rect 6000 34944 6052 34950
rect 6000 34886 6052 34892
rect 6012 34490 6040 34886
rect 6104 34610 6132 36110
rect 6196 35086 6224 37062
rect 6920 36100 6972 36106
rect 6920 36042 6972 36048
rect 6932 35834 6960 36042
rect 6920 35828 6972 35834
rect 6920 35770 6972 35776
rect 6276 35488 6328 35494
rect 6276 35430 6328 35436
rect 6184 35080 6236 35086
rect 6184 35022 6236 35028
rect 6092 34604 6144 34610
rect 6092 34546 6144 34552
rect 6012 34462 6132 34490
rect 6104 33998 6132 34462
rect 5908 33992 5960 33998
rect 5908 33934 5960 33940
rect 6092 33992 6144 33998
rect 6092 33934 6144 33940
rect 5724 31816 5776 31822
rect 5724 31758 5776 31764
rect 5448 30728 5500 30734
rect 5448 30670 5500 30676
rect 5632 30252 5684 30258
rect 5632 30194 5684 30200
rect 5356 28484 5408 28490
rect 5356 28426 5408 28432
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5460 26926 5488 27406
rect 5448 26920 5500 26926
rect 5448 26862 5500 26868
rect 5264 26852 5316 26858
rect 5264 26794 5316 26800
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5460 26353 5488 26726
rect 5446 26344 5502 26353
rect 5446 26279 5502 26288
rect 5540 25220 5592 25226
rect 5540 25162 5592 25168
rect 5552 24818 5580 25162
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5552 24274 5580 24754
rect 5540 24268 5592 24274
rect 5540 24210 5592 24216
rect 5552 23186 5580 24210
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 5460 23066 5488 23122
rect 5644 23066 5672 30194
rect 5920 27470 5948 33934
rect 6184 33856 6236 33862
rect 6184 33798 6236 33804
rect 6196 33386 6224 33798
rect 6184 33380 6236 33386
rect 6184 33322 6236 33328
rect 6092 32564 6144 32570
rect 6092 32506 6144 32512
rect 6000 28484 6052 28490
rect 6000 28426 6052 28432
rect 5908 27464 5960 27470
rect 5908 27406 5960 27412
rect 6012 26382 6040 28426
rect 6000 26376 6052 26382
rect 6000 26318 6052 26324
rect 6104 24818 6132 32506
rect 6184 32496 6236 32502
rect 6184 32438 6236 32444
rect 6196 31278 6224 32438
rect 6288 31754 6316 35430
rect 6736 35012 6788 35018
rect 6736 34954 6788 34960
rect 6644 33652 6696 33658
rect 6644 33594 6696 33600
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 6472 32366 6500 32506
rect 6460 32360 6512 32366
rect 6460 32302 6512 32308
rect 6552 32292 6604 32298
rect 6552 32234 6604 32240
rect 6460 32224 6512 32230
rect 6460 32166 6512 32172
rect 6288 31726 6408 31754
rect 6184 31272 6236 31278
rect 6184 31214 6236 31220
rect 6196 30734 6224 31214
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 6380 30258 6408 31726
rect 6472 31414 6500 32166
rect 6460 31408 6512 31414
rect 6460 31350 6512 31356
rect 6460 30660 6512 30666
rect 6460 30602 6512 30608
rect 6472 30394 6500 30602
rect 6460 30388 6512 30394
rect 6460 30330 6512 30336
rect 6368 30252 6420 30258
rect 6368 30194 6420 30200
rect 6564 28150 6592 32234
rect 6656 32230 6684 33594
rect 6748 33590 6776 34954
rect 6828 34604 6880 34610
rect 6828 34546 6880 34552
rect 6736 33584 6788 33590
rect 6736 33526 6788 33532
rect 6748 33114 6776 33526
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 6748 32910 6776 33050
rect 6736 32904 6788 32910
rect 6736 32846 6788 32852
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6840 32026 6868 34546
rect 7116 34406 7144 39986
rect 8588 37874 8616 40054
rect 9220 40044 9272 40050
rect 9220 39986 9272 39992
rect 9232 39642 9260 39986
rect 9220 39636 9272 39642
rect 9220 39578 9272 39584
rect 9680 39432 9732 39438
rect 9680 39374 9732 39380
rect 9692 38554 9720 39374
rect 9680 38548 9732 38554
rect 9680 38490 9732 38496
rect 9784 38418 9812 40122
rect 9772 38412 9824 38418
rect 9772 38354 9824 38360
rect 9876 38214 9904 40326
rect 9968 39914 9996 41006
rect 9956 39908 10008 39914
rect 9956 39850 10008 39856
rect 9968 39370 9996 39850
rect 10152 39794 10180 41074
rect 10968 40996 11020 41002
rect 10968 40938 11020 40944
rect 10508 40520 10560 40526
rect 10508 40462 10560 40468
rect 10232 40452 10284 40458
rect 10232 40394 10284 40400
rect 10244 39982 10272 40394
rect 10324 40112 10376 40118
rect 10324 40054 10376 40060
rect 10232 39976 10284 39982
rect 10232 39918 10284 39924
rect 10232 39840 10284 39846
rect 10152 39788 10232 39794
rect 10152 39782 10284 39788
rect 10152 39766 10272 39782
rect 10244 39370 10272 39766
rect 10336 39438 10364 40054
rect 10324 39432 10376 39438
rect 10324 39374 10376 39380
rect 9956 39364 10008 39370
rect 9956 39306 10008 39312
rect 10232 39364 10284 39370
rect 10232 39306 10284 39312
rect 9864 38208 9916 38214
rect 9864 38150 9916 38156
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 8576 37868 8628 37874
rect 8576 37810 8628 37816
rect 8312 36242 8340 37810
rect 8668 37664 8720 37670
rect 8668 37606 8720 37612
rect 8944 37664 8996 37670
rect 8944 37606 8996 37612
rect 8300 36236 8352 36242
rect 8300 36178 8352 36184
rect 7380 36100 7432 36106
rect 7380 36042 7432 36048
rect 8300 36100 8352 36106
rect 8300 36042 8352 36048
rect 7392 35698 7420 36042
rect 7380 35692 7432 35698
rect 7380 35634 7432 35640
rect 7656 35624 7708 35630
rect 7656 35566 7708 35572
rect 7564 35556 7616 35562
rect 7564 35498 7616 35504
rect 7472 34604 7524 34610
rect 7472 34546 7524 34552
rect 7104 34400 7156 34406
rect 7104 34342 7156 34348
rect 7116 34202 7144 34342
rect 7484 34202 7512 34546
rect 7104 34196 7156 34202
rect 7104 34138 7156 34144
rect 7472 34196 7524 34202
rect 7472 34138 7524 34144
rect 7116 33998 7144 34138
rect 7104 33992 7156 33998
rect 7156 33940 7236 33946
rect 7104 33934 7236 33940
rect 7116 33918 7236 33934
rect 7012 32972 7064 32978
rect 7012 32914 7064 32920
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6932 32434 6960 32710
rect 7024 32434 7052 32914
rect 7104 32836 7156 32842
rect 7104 32778 7156 32784
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 7012 32428 7064 32434
rect 7012 32370 7064 32376
rect 6828 32020 6880 32026
rect 6828 31962 6880 31968
rect 6840 30734 6868 31962
rect 7116 31142 7144 32778
rect 7104 31136 7156 31142
rect 7104 31078 7156 31084
rect 7104 30932 7156 30938
rect 7104 30874 7156 30880
rect 6828 30728 6880 30734
rect 6828 30670 6880 30676
rect 6736 28416 6788 28422
rect 6736 28358 6788 28364
rect 6552 28144 6604 28150
rect 6552 28086 6604 28092
rect 6748 26994 6776 28358
rect 6840 28082 6868 30670
rect 6920 30252 6972 30258
rect 6920 30194 6972 30200
rect 6932 29850 6960 30194
rect 6920 29844 6972 29850
rect 6920 29786 6972 29792
rect 7116 29646 7144 30874
rect 7104 29640 7156 29646
rect 7104 29582 7156 29588
rect 7012 29572 7064 29578
rect 7012 29514 7064 29520
rect 7024 28490 7052 29514
rect 7012 28484 7064 28490
rect 7012 28426 7064 28432
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 6932 27674 6960 28018
rect 6920 27668 6972 27674
rect 6920 27610 6972 27616
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6368 26376 6420 26382
rect 6368 26318 6420 26324
rect 6380 26042 6408 26318
rect 6564 26314 6592 26386
rect 6840 26382 6868 26930
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6552 26308 6604 26314
rect 6552 26250 6604 26256
rect 6736 26308 6788 26314
rect 6736 26250 6788 26256
rect 6368 26036 6420 26042
rect 6368 25978 6420 25984
rect 6748 25974 6776 26250
rect 6736 25968 6788 25974
rect 6736 25910 6788 25916
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6092 24812 6144 24818
rect 6092 24754 6144 24760
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 5828 23730 5856 24346
rect 6104 24138 6132 24754
rect 6840 24750 6868 25638
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 6460 24608 6512 24614
rect 6460 24550 6512 24556
rect 6472 24206 6500 24550
rect 6840 24274 6868 24686
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6460 24200 6512 24206
rect 6460 24142 6512 24148
rect 6092 24132 6144 24138
rect 6092 24074 6144 24080
rect 6828 24132 6880 24138
rect 6828 24074 6880 24080
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6288 23798 6316 24006
rect 6276 23792 6328 23798
rect 6276 23734 6328 23740
rect 5816 23724 5868 23730
rect 5816 23666 5868 23672
rect 5460 23038 5672 23066
rect 6288 23050 6316 23734
rect 6368 23656 6420 23662
rect 6368 23598 6420 23604
rect 6276 23044 6328 23050
rect 5552 22234 5580 23038
rect 6276 22986 6328 22992
rect 6288 22778 6316 22986
rect 6380 22982 6408 23598
rect 6368 22976 6420 22982
rect 6368 22918 6420 22924
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6380 22642 6408 22918
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6840 22386 6868 24074
rect 6920 23656 6972 23662
rect 6920 23598 6972 23604
rect 6932 23322 6960 23598
rect 6920 23316 6972 23322
rect 6920 23258 6972 23264
rect 6932 22574 6960 23258
rect 7116 22642 7144 27406
rect 7208 26466 7236 33918
rect 7472 33108 7524 33114
rect 7472 33050 7524 33056
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 7300 32366 7328 32506
rect 7288 32360 7340 32366
rect 7288 32302 7340 32308
rect 7392 32026 7420 32846
rect 7484 32502 7512 33050
rect 7472 32496 7524 32502
rect 7472 32438 7524 32444
rect 7380 32020 7432 32026
rect 7380 31962 7432 31968
rect 7576 30258 7604 35498
rect 7668 34066 7696 35566
rect 8312 35086 8340 36042
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8576 35012 8628 35018
rect 8576 34954 8628 34960
rect 7932 34944 7984 34950
rect 7932 34886 7984 34892
rect 7656 34060 7708 34066
rect 7656 34002 7708 34008
rect 7668 33046 7696 34002
rect 7944 33998 7972 34886
rect 8588 34746 8616 34954
rect 8576 34740 8628 34746
rect 8576 34682 8628 34688
rect 8208 34060 8260 34066
rect 8208 34002 8260 34008
rect 7932 33992 7984 33998
rect 7932 33934 7984 33940
rect 8024 33924 8076 33930
rect 8024 33866 8076 33872
rect 8036 33590 8064 33866
rect 8024 33584 8076 33590
rect 8024 33526 8076 33532
rect 7656 33040 7708 33046
rect 7656 32982 7708 32988
rect 7748 31136 7800 31142
rect 7748 31078 7800 31084
rect 7564 30252 7616 30258
rect 7564 30194 7616 30200
rect 7472 30184 7524 30190
rect 7472 30126 7524 30132
rect 7484 29102 7512 30126
rect 7576 30054 7604 30194
rect 7564 30048 7616 30054
rect 7564 29990 7616 29996
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 7380 28416 7432 28422
rect 7380 28358 7432 28364
rect 7392 27470 7420 28358
rect 7484 27538 7512 29038
rect 7472 27532 7524 27538
rect 7472 27474 7524 27480
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7208 26438 7328 26466
rect 7194 26344 7250 26353
rect 7194 26279 7250 26288
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 7116 22438 7144 22578
rect 6656 22358 6868 22386
rect 7012 22432 7064 22438
rect 7012 22374 7064 22380
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 5540 22228 5592 22234
rect 5540 22170 5592 22176
rect 5552 22094 5580 22170
rect 5184 22066 5304 22094
rect 5552 22066 5764 22094
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4908 17338 4936 19790
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4804 14816 4856 14822
rect 4804 14758 4856 14764
rect 4816 14482 4844 14758
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4816 14006 4844 14418
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4908 12986 4936 17138
rect 5000 15978 5028 22066
rect 5276 22001 5304 22066
rect 5262 21992 5318 22001
rect 5262 21927 5318 21936
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5184 17542 5212 18158
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 4988 15972 5040 15978
rect 4988 15914 5040 15920
rect 5184 15366 5212 17478
rect 5276 17338 5304 21927
rect 5736 19990 5764 22066
rect 6656 20534 6684 22358
rect 6736 22228 6788 22234
rect 6736 22170 6788 22176
rect 6748 21622 6776 22170
rect 7024 21962 7052 22374
rect 7012 21956 7064 21962
rect 7012 21898 7064 21904
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 6932 20602 6960 20810
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 6184 19780 6236 19786
rect 6184 19722 6236 19728
rect 5736 19174 5764 19722
rect 6196 19174 6224 19722
rect 5724 19168 5776 19174
rect 5722 19136 5724 19145
rect 6184 19168 6236 19174
rect 5776 19136 5778 19145
rect 6184 19110 6236 19116
rect 5722 19071 5778 19080
rect 6196 18714 6224 19110
rect 6104 18686 6224 18714
rect 6828 18692 6880 18698
rect 6104 18426 6132 18686
rect 6828 18634 6880 18640
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6196 18290 6224 18566
rect 6840 18426 6868 18634
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 5540 18216 5592 18222
rect 5540 18158 5592 18164
rect 5552 17678 5580 18158
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5276 16794 5304 17138
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5276 15706 5304 16730
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5368 15434 5396 16526
rect 5448 16244 5500 16250
rect 5448 16186 5500 16192
rect 5356 15428 5408 15434
rect 5356 15370 5408 15376
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 14346 5212 15302
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 4724 12406 4936 12434
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11218 4660 11562
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10674 4292 10950
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4632 10606 4660 11018
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 9994 4660 10542
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4632 9738 4660 9930
rect 4632 9710 4752 9738
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3528 4078 3556 6122
rect 3620 5778 3648 6190
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3804 4706 3832 8502
rect 3896 6254 3924 9046
rect 3988 9042 4016 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4632 8974 4660 9454
rect 4724 9042 4752 9710
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4632 8430 4660 8910
rect 4620 8424 4672 8430
rect 3974 8392 4030 8401
rect 4620 8366 4672 8372
rect 3974 8327 3976 8336
rect 4028 8327 4030 8336
rect 3976 8298 4028 8304
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 8090 4108 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3988 7546 4016 7754
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 3882 5536 3938 5545
rect 3882 5471 3938 5480
rect 3896 4826 3924 5471
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3804 4678 3924 4706
rect 3792 4616 3844 4622
rect 3790 4584 3792 4593
rect 3844 4584 3846 4593
rect 3790 4519 3846 4528
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 3804 2514 3832 4218
rect 3896 2774 3924 4678
rect 3988 4282 4016 6598
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 4080 4146 4108 6326
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4540 5114 4568 5646
rect 4632 5302 4660 6598
rect 4620 5296 4672 5302
rect 4620 5238 4672 5244
rect 4540 5086 4660 5114
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4570 4660 5086
rect 4540 4542 4660 4570
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4080 3398 4108 4082
rect 4540 4010 4568 4542
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4010 4660 4422
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4724 2854 4752 7822
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 4622 4844 7142
rect 4908 6458 4936 12406
rect 5276 9738 5304 12922
rect 5368 11626 5396 15370
rect 5460 12170 5488 16186
rect 5920 15502 5948 17614
rect 6196 17542 6224 18226
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5828 14482 5856 15302
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5920 14414 5948 15438
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5828 12442 5856 13738
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5920 12322 5948 14350
rect 5828 12294 5948 12322
rect 5828 12238 5856 12294
rect 6012 12238 6040 16934
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5356 11620 5408 11626
rect 5356 11562 5408 11568
rect 5276 9710 5396 9738
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5276 9382 5304 9522
rect 5264 9376 5316 9382
rect 5262 9344 5264 9353
rect 5316 9344 5318 9353
rect 5262 9279 5318 9288
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4908 5710 4936 6394
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 5234 4936 5510
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4816 2990 4844 4558
rect 4908 4078 4936 5170
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 5000 3097 5028 8774
rect 5368 8430 5396 9710
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5092 3534 5120 6054
rect 5184 5234 5212 6258
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5184 3738 5212 5170
rect 5368 4826 5396 8366
rect 5460 6662 5488 12106
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11218 5672 11494
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5538 11112 5594 11121
rect 5736 11082 5764 12038
rect 5538 11047 5540 11056
rect 5592 11047 5594 11056
rect 5724 11076 5776 11082
rect 5540 11018 5592 11024
rect 5724 11018 5776 11024
rect 5828 10674 5856 12174
rect 5920 11218 5948 12174
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11694 6040 12038
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6000 11552 6052 11558
rect 6000 11494 6052 11500
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5920 10742 5948 11154
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5540 9444 5592 9450
rect 5540 9386 5592 9392
rect 5552 8498 5580 9386
rect 5644 8498 5672 9454
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5552 6254 5580 8026
rect 5736 7886 5764 8842
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5828 7954 5856 8230
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5632 6180 5684 6186
rect 5632 6122 5684 6128
rect 5644 5794 5672 6122
rect 5736 5914 5764 6258
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5644 5766 5764 5794
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5264 4752 5316 4758
rect 5316 4700 5396 4706
rect 5264 4694 5396 4700
rect 5276 4678 5396 4694
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3534 5304 4490
rect 5368 4214 5396 4678
rect 5460 4622 5488 5578
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5356 3936 5408 3942
rect 5354 3904 5356 3913
rect 5408 3904 5410 3913
rect 5354 3839 5410 3848
rect 5460 3670 5488 4558
rect 5552 4486 5580 5646
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5538 4040 5594 4049
rect 5538 3975 5594 3984
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5080 3120 5132 3126
rect 4986 3088 5042 3097
rect 5080 3062 5132 3068
rect 4986 3023 4988 3032
rect 5040 3023 5042 3032
rect 4988 2994 5040 3000
rect 4804 2984 4856 2990
rect 5000 2963 5028 2994
rect 4804 2926 4856 2932
rect 5092 2854 5120 3062
rect 5354 2952 5410 2961
rect 5354 2887 5410 2896
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 3896 2746 4108 2774
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 4080 2446 4108 2746
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5000 2514 5028 2790
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 5276 2106 5304 2518
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 3056 1420 3108 1426
rect 3056 1362 3108 1368
rect 5368 1358 5396 2887
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5552 800 5580 3975
rect 5644 3738 5672 4966
rect 5736 3942 5764 5766
rect 5828 4570 5856 7686
rect 5920 7478 5948 7822
rect 5908 7472 5960 7478
rect 5908 7414 5960 7420
rect 6012 6662 6040 11494
rect 6104 11218 6132 14282
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6104 10130 6132 11154
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6196 8634 6224 17478
rect 6656 17202 6684 17478
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6656 16998 6684 17138
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6932 16250 6960 20538
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 19718 7144 20402
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7116 17134 7144 18158
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6288 14414 6316 14486
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6288 12434 6316 14350
rect 6460 13864 6512 13870
rect 6458 13832 6460 13841
rect 6512 13832 6514 13841
rect 6458 13767 6514 13776
rect 6288 12406 6408 12434
rect 6380 11762 6408 12406
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11558 6408 11698
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 8974 6316 9998
rect 6380 9586 6408 10542
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6288 8430 6316 8910
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6104 6866 6132 7822
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6012 6322 6040 6598
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6196 5250 6224 7686
rect 6288 5574 6316 8366
rect 6472 8022 6500 12174
rect 6656 11762 6684 15846
rect 7208 15706 7236 26279
rect 7300 23254 7328 26438
rect 7288 23248 7340 23254
rect 7288 23190 7340 23196
rect 7300 22234 7328 23190
rect 7288 22228 7340 22234
rect 7288 22170 7340 22176
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7300 17338 7328 17546
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7300 15586 7328 17070
rect 7392 15706 7420 26726
rect 7484 26518 7512 27474
rect 7576 27470 7604 29990
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7760 27062 7788 31078
rect 8220 30938 8248 34002
rect 8588 33930 8616 34682
rect 8576 33924 8628 33930
rect 8576 33866 8628 33872
rect 8300 33856 8352 33862
rect 8300 33798 8352 33804
rect 8312 33658 8340 33798
rect 8300 33652 8352 33658
rect 8300 33594 8352 33600
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 8208 28484 8260 28490
rect 8208 28426 8260 28432
rect 8220 28218 8248 28426
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8680 28082 8708 37606
rect 8956 33998 8984 37606
rect 9968 36106 9996 39306
rect 10140 36780 10192 36786
rect 10140 36722 10192 36728
rect 10152 36378 10180 36722
rect 10140 36372 10192 36378
rect 10140 36314 10192 36320
rect 9956 36100 10008 36106
rect 9956 36042 10008 36048
rect 10244 35698 10272 39306
rect 10336 38350 10364 39374
rect 10520 38758 10548 40462
rect 10600 40384 10652 40390
rect 10600 40326 10652 40332
rect 10612 39370 10640 40326
rect 10692 40044 10744 40050
rect 10692 39986 10744 39992
rect 10704 39642 10732 39986
rect 10692 39636 10744 39642
rect 10692 39578 10744 39584
rect 10600 39364 10652 39370
rect 10600 39306 10652 39312
rect 10508 38752 10560 38758
rect 10508 38694 10560 38700
rect 10324 38344 10376 38350
rect 10324 38286 10376 38292
rect 10336 37262 10364 38286
rect 10324 37256 10376 37262
rect 10324 37198 10376 37204
rect 10336 35766 10364 37198
rect 10416 37188 10468 37194
rect 10416 37130 10468 37136
rect 10428 36922 10456 37130
rect 10416 36916 10468 36922
rect 10416 36858 10468 36864
rect 10520 36854 10548 38694
rect 10612 37738 10640 39306
rect 10600 37732 10652 37738
rect 10600 37674 10652 37680
rect 10600 37120 10652 37126
rect 10600 37062 10652 37068
rect 10508 36848 10560 36854
rect 10508 36790 10560 36796
rect 10520 36038 10548 36790
rect 10612 36174 10640 37062
rect 10600 36168 10652 36174
rect 10600 36110 10652 36116
rect 10876 36168 10928 36174
rect 10876 36110 10928 36116
rect 10416 36032 10468 36038
rect 10416 35974 10468 35980
rect 10508 36032 10560 36038
rect 10508 35974 10560 35980
rect 10324 35760 10376 35766
rect 10324 35702 10376 35708
rect 10232 35692 10284 35698
rect 10232 35634 10284 35640
rect 10244 34610 10272 35634
rect 10232 34604 10284 34610
rect 10232 34546 10284 34552
rect 9864 34060 9916 34066
rect 9864 34002 9916 34008
rect 8944 33992 8996 33998
rect 8944 33934 8996 33940
rect 9588 33856 9640 33862
rect 9588 33798 9640 33804
rect 9128 33516 9180 33522
rect 9128 33458 9180 33464
rect 9036 33108 9088 33114
rect 9036 33050 9088 33056
rect 8944 31884 8996 31890
rect 8944 31826 8996 31832
rect 8956 29714 8984 31826
rect 8944 29708 8996 29714
rect 8944 29650 8996 29656
rect 8668 28076 8720 28082
rect 8668 28018 8720 28024
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 8956 27538 8984 28018
rect 8944 27532 8996 27538
rect 8944 27474 8996 27480
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 7748 27056 7800 27062
rect 7748 26998 7800 27004
rect 8128 26586 8156 27270
rect 8956 27130 8984 27474
rect 8944 27124 8996 27130
rect 8944 27066 8996 27072
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 7472 26512 7524 26518
rect 7472 26454 7524 26460
rect 7484 26246 7512 26454
rect 7576 26314 7604 26522
rect 7564 26308 7616 26314
rect 7564 26250 7616 26256
rect 7472 26240 7524 26246
rect 7472 26182 7524 26188
rect 9048 25498 9076 33050
rect 9140 32434 9168 33458
rect 9128 32428 9180 32434
rect 9128 32370 9180 32376
rect 9404 32428 9456 32434
rect 9404 32370 9456 32376
rect 9416 30598 9444 32370
rect 9404 30592 9456 30598
rect 9404 30534 9456 30540
rect 9416 28558 9444 30534
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9508 29646 9536 29990
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 9312 28552 9364 28558
rect 9312 28494 9364 28500
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9324 28422 9352 28494
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 9140 26994 9168 28018
rect 9220 27872 9272 27878
rect 9220 27814 9272 27820
rect 9128 26988 9180 26994
rect 9128 26930 9180 26936
rect 9036 25492 9088 25498
rect 9036 25434 9088 25440
rect 9048 25294 9076 25434
rect 9036 25288 9088 25294
rect 9036 25230 9088 25236
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 8036 24342 8064 24550
rect 8024 24336 8076 24342
rect 8024 24278 8076 24284
rect 7472 23588 7524 23594
rect 7472 23530 7524 23536
rect 7484 22574 7512 23530
rect 7472 22568 7524 22574
rect 7472 22510 7524 22516
rect 7484 22234 7512 22510
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7576 19922 7604 22374
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7760 21486 7788 21966
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 7760 20874 7788 21422
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 7760 20398 7788 20810
rect 7944 20806 7972 21558
rect 7932 20800 7984 20806
rect 7932 20742 7984 20748
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7564 19916 7616 19922
rect 7564 19858 7616 19864
rect 7760 18834 7788 20334
rect 7944 19378 7972 20742
rect 7932 19372 7984 19378
rect 7932 19314 7984 19320
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 18290 8432 18566
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7668 17134 7696 17478
rect 7760 17202 7788 17478
rect 7944 17202 7972 18226
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7654 16144 7710 16153
rect 7654 16079 7656 16088
rect 7708 16079 7710 16088
rect 7656 16050 7708 16056
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7944 15638 7972 17138
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 7208 15558 7328 15586
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 8208 15564 8260 15570
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 6932 14618 6960 14962
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7024 14346 7052 15302
rect 7208 14482 7236 15558
rect 8208 15506 8260 15512
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 7012 12708 7064 12714
rect 7012 12650 7064 12656
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6932 11898 6960 12310
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 7024 11762 7052 12650
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 6656 11121 6684 11154
rect 6828 11144 6880 11150
rect 6642 11112 6698 11121
rect 6828 11086 6880 11092
rect 6642 11047 6698 11056
rect 6840 9518 6868 11086
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6840 9042 6868 9454
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 8498 6776 8842
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6748 7954 6776 8434
rect 6932 8294 6960 8774
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 7024 7886 7052 9522
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7024 7562 7052 7822
rect 6840 7534 7052 7562
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6104 5222 6224 5250
rect 6288 5234 6316 5510
rect 6380 5370 6408 6054
rect 6472 5778 6500 6258
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6472 5574 6500 5714
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6276 5228 6328 5234
rect 5906 4584 5962 4593
rect 5828 4542 5906 4570
rect 5906 4519 5962 4528
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5814 3904 5870 3913
rect 5814 3839 5870 3848
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5644 2689 5672 3334
rect 5736 3194 5764 3402
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5828 3058 5856 3839
rect 5920 3194 5948 4519
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 5630 2680 5686 2689
rect 5630 2615 5686 2624
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5644 800 5672 2382
rect 5736 800 5764 2858
rect 5828 800 5856 2858
rect 5920 2650 5948 2994
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6104 2446 6132 5222
rect 6276 5170 6328 5176
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6196 2774 6224 4966
rect 6276 4616 6328 4622
rect 6380 4604 6408 5306
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6472 4826 6500 5238
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6328 4576 6408 4604
rect 6276 4558 6328 4564
rect 6564 4146 6592 6598
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6288 3058 6316 3878
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6196 2746 6316 2774
rect 6182 2680 6238 2689
rect 6182 2615 6238 2624
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 5920 1562 5948 2246
rect 5908 1556 5960 1562
rect 5908 1498 5960 1504
rect 5908 1420 5960 1426
rect 5908 1362 5960 1368
rect 5920 800 5948 1362
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 6012 800 6040 1294
rect 6104 800 6132 2382
rect 6196 800 6224 2615
rect 6288 800 6316 2746
rect 6380 800 6408 4014
rect 6656 4010 6684 5102
rect 6748 4622 6776 5850
rect 6840 5710 6868 7534
rect 7116 5710 7144 14350
rect 7208 12434 7236 14418
rect 7760 14414 7788 14758
rect 8220 14414 8248 15506
rect 8312 15502 8340 16662
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13870 7328 14214
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7208 12406 7328 12434
rect 7300 11694 7328 12406
rect 7392 11898 7420 12786
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8128 12374 8156 12718
rect 8496 12434 8524 19110
rect 8588 18358 8616 19110
rect 9048 18970 9076 25230
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 9232 17882 9260 27814
rect 9600 26874 9628 33798
rect 9876 32910 9904 34002
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 10232 33992 10284 33998
rect 10232 33934 10284 33940
rect 10152 33590 10180 33934
rect 10140 33584 10192 33590
rect 10140 33526 10192 33532
rect 10048 32972 10100 32978
rect 10048 32914 10100 32920
rect 9864 32904 9916 32910
rect 9864 32846 9916 32852
rect 9956 32904 10008 32910
rect 9956 32846 10008 32852
rect 9968 32502 9996 32846
rect 9956 32496 10008 32502
rect 9956 32438 10008 32444
rect 9968 32026 9996 32438
rect 9956 32020 10008 32026
rect 9956 31962 10008 31968
rect 9680 31748 9732 31754
rect 9680 31690 9732 31696
rect 9692 31482 9720 31690
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 10060 31346 10088 32914
rect 10140 32224 10192 32230
rect 10140 32166 10192 32172
rect 10152 31346 10180 32166
rect 9864 31340 9916 31346
rect 9864 31282 9916 31288
rect 10029 31340 10088 31346
rect 10081 31288 10088 31340
rect 10029 31282 10088 31288
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 9876 31210 9904 31282
rect 9864 31204 9916 31210
rect 9864 31146 9916 31152
rect 9680 30728 9732 30734
rect 9680 30670 9732 30676
rect 9692 29102 9720 30670
rect 10060 30122 10088 31282
rect 10244 31278 10272 33934
rect 10336 33658 10364 35702
rect 10428 34066 10456 35974
rect 10520 35154 10548 35974
rect 10888 35766 10916 36110
rect 10980 35766 11008 40938
rect 11532 40934 11560 41386
rect 11428 40928 11480 40934
rect 11428 40870 11480 40876
rect 11520 40928 11572 40934
rect 11520 40870 11572 40876
rect 11704 40928 11756 40934
rect 11704 40870 11756 40876
rect 11440 40118 11468 40870
rect 11428 40112 11480 40118
rect 11428 40054 11480 40060
rect 11612 40044 11664 40050
rect 11612 39986 11664 39992
rect 11624 39846 11652 39986
rect 11612 39840 11664 39846
rect 11612 39782 11664 39788
rect 11624 38758 11652 39782
rect 11612 38752 11664 38758
rect 11612 38694 11664 38700
rect 11716 36922 11744 40870
rect 12084 39098 12112 41550
rect 12176 41206 12204 42298
rect 12728 42226 12756 42638
rect 14648 42628 14700 42634
rect 14648 42570 14700 42576
rect 16304 42628 16356 42634
rect 16304 42570 16356 42576
rect 14660 42294 14688 42570
rect 14924 42560 14976 42566
rect 14924 42502 14976 42508
rect 15936 42560 15988 42566
rect 15936 42502 15988 42508
rect 14648 42288 14700 42294
rect 14648 42230 14700 42236
rect 12716 42220 12768 42226
rect 12716 42162 12768 42168
rect 12900 42220 12952 42226
rect 12900 42162 12952 42168
rect 13912 42220 13964 42226
rect 13912 42162 13964 42168
rect 12716 42084 12768 42090
rect 12716 42026 12768 42032
rect 12440 42016 12492 42022
rect 12440 41958 12492 41964
rect 12452 41206 12480 41958
rect 12728 41682 12756 42026
rect 12912 41818 12940 42162
rect 12992 42084 13044 42090
rect 12992 42026 13044 42032
rect 12900 41812 12952 41818
rect 12900 41754 12952 41760
rect 12716 41676 12768 41682
rect 12716 41618 12768 41624
rect 12532 41268 12584 41274
rect 12532 41210 12584 41216
rect 12164 41200 12216 41206
rect 12164 41142 12216 41148
rect 12440 41200 12492 41206
rect 12440 41142 12492 41148
rect 12072 39092 12124 39098
rect 12072 39034 12124 39040
rect 11980 37936 12032 37942
rect 11980 37878 12032 37884
rect 11992 37330 12020 37878
rect 11980 37324 12032 37330
rect 11980 37266 12032 37272
rect 11704 36916 11756 36922
rect 11704 36858 11756 36864
rect 10876 35760 10928 35766
rect 10876 35702 10928 35708
rect 10968 35760 11020 35766
rect 10968 35702 11020 35708
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 10692 35488 10744 35494
rect 10692 35430 10744 35436
rect 10508 35148 10560 35154
rect 10508 35090 10560 35096
rect 10600 34536 10652 34542
rect 10600 34478 10652 34484
rect 10416 34060 10468 34066
rect 10416 34002 10468 34008
rect 10612 33930 10640 34478
rect 10704 33998 10732 35430
rect 11900 35290 11928 35634
rect 11888 35284 11940 35290
rect 11888 35226 11940 35232
rect 11152 35012 11204 35018
rect 11152 34954 11204 34960
rect 11164 34202 11192 34954
rect 12084 34746 12112 39034
rect 12176 38486 12204 41142
rect 12544 41018 12572 41210
rect 12452 40990 12572 41018
rect 12452 40390 12480 40990
rect 12532 40452 12584 40458
rect 12532 40394 12584 40400
rect 12440 40384 12492 40390
rect 12440 40326 12492 40332
rect 12452 39794 12480 40326
rect 12544 39982 12572 40394
rect 12532 39976 12584 39982
rect 12728 39964 12756 41618
rect 13004 41614 13032 42026
rect 12992 41608 13044 41614
rect 12992 41550 13044 41556
rect 12900 41064 12952 41070
rect 12900 41006 12952 41012
rect 12912 40526 12940 41006
rect 12900 40520 12952 40526
rect 12900 40462 12952 40468
rect 13004 40050 13032 41550
rect 13924 41414 13952 42162
rect 14556 42016 14608 42022
rect 14556 41958 14608 41964
rect 14568 41614 14596 41958
rect 14556 41608 14608 41614
rect 14556 41550 14608 41556
rect 14936 41546 14964 42502
rect 15384 42220 15436 42226
rect 15384 42162 15436 42168
rect 15476 42220 15528 42226
rect 15476 42162 15528 42168
rect 15752 42220 15804 42226
rect 15752 42162 15804 42168
rect 15396 41818 15424 42162
rect 15488 42090 15516 42162
rect 15476 42084 15528 42090
rect 15476 42026 15528 42032
rect 15384 41812 15436 41818
rect 15384 41754 15436 41760
rect 14924 41540 14976 41546
rect 14924 41482 14976 41488
rect 14096 41472 14148 41478
rect 14096 41414 14148 41420
rect 13832 41386 13952 41414
rect 13832 40934 13860 41386
rect 14108 41206 14136 41414
rect 14096 41200 14148 41206
rect 14096 41142 14148 41148
rect 14924 41132 14976 41138
rect 14924 41074 14976 41080
rect 13820 40928 13872 40934
rect 13820 40870 13872 40876
rect 12992 40044 13044 40050
rect 12992 39986 13044 39992
rect 12900 39976 12952 39982
rect 12728 39936 12900 39964
rect 12532 39918 12584 39924
rect 12900 39918 12952 39924
rect 13360 39976 13412 39982
rect 13360 39918 13412 39924
rect 12452 39766 12572 39794
rect 12164 38480 12216 38486
rect 12164 38422 12216 38428
rect 12440 38344 12492 38350
rect 12440 38286 12492 38292
rect 12452 36854 12480 38286
rect 12256 36848 12308 36854
rect 12256 36790 12308 36796
rect 12440 36848 12492 36854
rect 12440 36790 12492 36796
rect 12268 36582 12296 36790
rect 12256 36576 12308 36582
rect 12256 36518 12308 36524
rect 12440 36100 12492 36106
rect 12440 36042 12492 36048
rect 12452 35834 12480 36042
rect 12440 35828 12492 35834
rect 12440 35770 12492 35776
rect 12544 35154 12572 39766
rect 13372 38894 13400 39918
rect 13360 38888 13412 38894
rect 13360 38830 13412 38836
rect 13268 38820 13320 38826
rect 13268 38762 13320 38768
rect 13280 38554 13308 38762
rect 13268 38548 13320 38554
rect 13268 38490 13320 38496
rect 13544 38548 13596 38554
rect 13544 38490 13596 38496
rect 12624 38344 12676 38350
rect 12624 38286 12676 38292
rect 12992 38344 13044 38350
rect 12992 38286 13044 38292
rect 12636 38214 12664 38286
rect 12808 38276 12860 38282
rect 12808 38218 12860 38224
rect 12624 38208 12676 38214
rect 12624 38150 12676 38156
rect 12820 37942 12848 38218
rect 12808 37936 12860 37942
rect 12808 37878 12860 37884
rect 13004 37874 13032 38286
rect 12992 37868 13044 37874
rect 12992 37810 13044 37816
rect 12808 37800 12860 37806
rect 12808 37742 12860 37748
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 12636 36718 12664 37198
rect 12716 36848 12768 36854
rect 12716 36790 12768 36796
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12532 35148 12584 35154
rect 12532 35090 12584 35096
rect 12440 35012 12492 35018
rect 12636 35000 12664 36654
rect 12492 34972 12664 35000
rect 12440 34954 12492 34960
rect 12072 34740 12124 34746
rect 12072 34682 12124 34688
rect 12084 34610 12112 34682
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 11152 34196 11204 34202
rect 11152 34138 11204 34144
rect 10692 33992 10744 33998
rect 10692 33934 10744 33940
rect 10600 33924 10652 33930
rect 10600 33866 10652 33872
rect 10324 33652 10376 33658
rect 10324 33594 10376 33600
rect 10612 33522 10640 33866
rect 10600 33516 10652 33522
rect 10600 33458 10652 33464
rect 10508 31340 10560 31346
rect 10508 31282 10560 31288
rect 10232 31272 10284 31278
rect 10232 31214 10284 31220
rect 10140 30252 10192 30258
rect 10140 30194 10192 30200
rect 10048 30116 10100 30122
rect 10048 30058 10100 30064
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9692 28626 9720 29038
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9968 28558 9996 29446
rect 10060 28694 10088 30058
rect 10152 28762 10180 30194
rect 10244 30190 10272 31214
rect 10520 31210 10548 31282
rect 10508 31204 10560 31210
rect 10508 31146 10560 31152
rect 10232 30184 10284 30190
rect 10232 30126 10284 30132
rect 10140 28756 10192 28762
rect 10140 28698 10192 28704
rect 10048 28688 10100 28694
rect 10048 28630 10100 28636
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9772 28416 9824 28422
rect 9772 28358 9824 28364
rect 9784 27878 9812 28358
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9784 27470 9812 27814
rect 9772 27464 9824 27470
rect 9772 27406 9824 27412
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9968 26994 9996 27406
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 9508 26846 9628 26874
rect 9312 22704 9364 22710
rect 9312 22646 9364 22652
rect 9324 22030 9352 22646
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9416 21690 9444 22578
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9508 19242 9536 26846
rect 9680 25900 9732 25906
rect 9680 25842 9732 25848
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9600 24886 9628 25094
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9588 24064 9640 24070
rect 9692 24052 9720 25842
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9784 24070 9812 25774
rect 10140 25424 10192 25430
rect 10140 25366 10192 25372
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9864 24608 9916 24614
rect 9864 24550 9916 24556
rect 9876 24138 9904 24550
rect 10060 24274 10088 25230
rect 10152 24886 10180 25366
rect 10140 24880 10192 24886
rect 10140 24822 10192 24828
rect 10048 24268 10100 24274
rect 10048 24210 10100 24216
rect 9864 24132 9916 24138
rect 9864 24074 9916 24080
rect 9640 24024 9720 24052
rect 9588 24006 9640 24012
rect 9692 21962 9720 24024
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 22642 9812 23054
rect 9876 22710 9904 24074
rect 9864 22704 9916 22710
rect 9864 22646 9916 22652
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9784 22030 9812 22578
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9680 20936 9732 20942
rect 9680 20878 9732 20884
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9220 17876 9272 17882
rect 9220 17818 9272 17824
rect 9324 17678 9352 18226
rect 9600 18222 9628 18702
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9600 17746 9628 18158
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9324 17338 9352 17614
rect 9416 17338 9444 17614
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9692 17066 9720 20878
rect 9784 17202 9812 21830
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9680 17060 9732 17066
rect 9680 17002 9732 17008
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 16114 9444 16934
rect 9692 16794 9720 17002
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9968 16590 9996 22374
rect 10152 21672 10180 24822
rect 10060 21644 10180 21672
rect 10060 18426 10088 21644
rect 10140 21548 10192 21554
rect 10140 21490 10192 21496
rect 10152 21146 10180 21490
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 10244 21010 10272 30126
rect 10416 27328 10468 27334
rect 10416 27270 10468 27276
rect 10428 26314 10456 27270
rect 10416 26308 10468 26314
rect 10416 26250 10468 26256
rect 10324 24608 10376 24614
rect 10324 24550 10376 24556
rect 10336 24206 10364 24550
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10336 22778 10364 23666
rect 10428 23662 10456 26250
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10520 22094 10548 31146
rect 10612 26382 10640 33458
rect 10692 33380 10744 33386
rect 10692 33322 10744 33328
rect 10704 28082 10732 33322
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11992 32570 12020 32778
rect 11980 32564 12032 32570
rect 11980 32506 12032 32512
rect 11060 31816 11112 31822
rect 11060 31758 11112 31764
rect 10784 30728 10836 30734
rect 10784 30670 10836 30676
rect 10796 30394 10824 30670
rect 11072 30598 11100 31758
rect 11704 31204 11756 31210
rect 11704 31146 11756 31152
rect 11060 30592 11112 30598
rect 11060 30534 11112 30540
rect 10784 30388 10836 30394
rect 10784 30330 10836 30336
rect 10796 30122 10824 30330
rect 10784 30116 10836 30122
rect 10784 30058 10836 30064
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 10876 26920 10928 26926
rect 10876 26862 10928 26868
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10796 24818 10824 25638
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10428 22066 10548 22094
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10428 20806 10456 22066
rect 10508 21072 10560 21078
rect 10508 21014 10560 21020
rect 10520 20942 10548 21014
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10416 20800 10468 20806
rect 10416 20742 10468 20748
rect 10520 20602 10548 20878
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10796 20466 10824 20878
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10140 20256 10192 20262
rect 10140 20198 10192 20204
rect 10152 19786 10180 20198
rect 10336 19854 10364 20402
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10612 20058 10640 20266
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 10060 17202 10088 17546
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 10152 16590 10180 19722
rect 10428 19514 10456 19722
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 10244 18970 10272 19178
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10244 17542 10272 17682
rect 10508 17672 10560 17678
rect 10506 17640 10508 17649
rect 10560 17640 10562 17649
rect 10506 17575 10562 17584
rect 10520 17542 10548 17575
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10244 16114 10272 17478
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10428 16590 10456 17070
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10336 16182 10364 16458
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 10232 16108 10284 16114
rect 10520 16096 10548 17478
rect 10692 17264 10744 17270
rect 10692 17206 10744 17212
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10232 16050 10284 16056
rect 10428 16068 10548 16096
rect 10060 15910 10088 16050
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9416 13938 9444 15438
rect 9956 15360 10008 15366
rect 9956 15302 10008 15308
rect 9588 14272 9640 14278
rect 9586 14240 9588 14249
rect 9640 14240 9642 14249
rect 9586 14175 9642 14184
rect 9600 13954 9628 14175
rect 9600 13938 9904 13954
rect 9404 13932 9456 13938
rect 9600 13932 9916 13938
rect 9600 13926 9864 13932
rect 9404 13874 9456 13880
rect 9864 13874 9916 13880
rect 8576 13320 8628 13326
rect 8576 13262 8628 13268
rect 8588 12782 8616 13262
rect 9128 12844 9180 12850
rect 9128 12786 9180 12792
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8496 12406 8616 12434
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7208 10062 7236 10950
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7208 8974 7236 9998
rect 7300 9926 7328 11630
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 11082 7420 11562
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7208 8566 7236 8910
rect 7196 8560 7248 8566
rect 7196 8502 7248 8508
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 6866 7236 7686
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6840 4468 6868 5510
rect 6932 5234 6960 5646
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6748 4440 6868 4468
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6472 800 6500 3470
rect 6564 800 6592 3606
rect 6656 3466 6684 3946
rect 6748 3602 6776 4440
rect 6826 4312 6882 4321
rect 6826 4247 6828 4256
rect 6880 4247 6882 4256
rect 6828 4218 6880 4224
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6644 3460 6696 3466
rect 6644 3402 6696 3408
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6642 2680 6698 2689
rect 6642 2615 6644 2624
rect 6696 2615 6698 2624
rect 6644 2586 6696 2592
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6656 800 6684 2042
rect 6840 800 6868 2994
rect 6932 800 6960 4150
rect 7024 2836 7052 5510
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7116 4758 7144 5034
rect 7104 4752 7156 4758
rect 7104 4694 7156 4700
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7116 3126 7144 4558
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 7024 2808 7144 2836
rect 7116 1170 7144 2808
rect 7208 2446 7236 6666
rect 7300 6390 7328 9862
rect 7392 8974 7420 11018
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7852 9654 7880 10610
rect 7944 9654 7972 11494
rect 8128 9674 8156 12310
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11762 8432 12174
rect 8496 11830 8524 12242
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8496 9674 8524 11766
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7932 9648 7984 9654
rect 8128 9646 8248 9674
rect 7932 9590 7984 9596
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7392 5817 7420 8910
rect 7852 8634 7880 9590
rect 8220 9586 8248 9646
rect 8404 9646 8524 9674
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7484 6866 7512 8502
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7576 6644 7604 8366
rect 8404 8362 8432 9646
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8404 7818 8432 8298
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6798 7696 7142
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7576 6616 7696 6644
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 7576 5914 7604 6190
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7378 5808 7434 5817
rect 7378 5743 7434 5752
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7024 1142 7144 1170
rect 7024 800 7052 1142
rect 7208 800 7236 2382
rect 7300 800 7328 4082
rect 7392 2990 7420 5578
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7576 4282 7604 5170
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7668 4162 7696 6616
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7576 4134 7696 4162
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7484 2514 7512 4082
rect 7576 3738 7604 4134
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7380 2304 7432 2310
rect 7380 2246 7432 2252
rect 7392 800 7420 2246
rect 7472 1896 7524 1902
rect 7472 1838 7524 1844
rect 7484 1426 7512 1838
rect 7472 1420 7524 1426
rect 7472 1362 7524 1368
rect 7576 800 7604 3130
rect 7668 800 7696 3674
rect 7760 3058 7788 7686
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 6866 7880 7346
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7852 5409 7880 6326
rect 7838 5400 7894 5409
rect 7838 5335 7894 5344
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7748 1556 7800 1562
rect 7748 1498 7800 1504
rect 7760 800 7788 1498
rect 7852 1442 7880 3130
rect 7944 2378 7972 7482
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8036 6458 8064 6802
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 8024 6316 8076 6322
rect 8076 6276 8156 6304
rect 8024 6258 8076 6264
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 8036 5234 8064 5782
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8036 4622 8064 5170
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8022 4040 8078 4049
rect 8022 3975 8078 3984
rect 8036 3398 8064 3975
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7932 2372 7984 2378
rect 7932 2314 7984 2320
rect 7944 1766 7972 2314
rect 7932 1760 7984 1766
rect 7932 1702 7984 1708
rect 7852 1414 7972 1442
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 7852 800 7880 1294
rect 7944 800 7972 1414
rect 8036 800 8064 2790
rect 8128 800 8156 6276
rect 8220 2378 8248 6734
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8312 4826 8340 6258
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8404 5710 8432 6122
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8312 4146 8340 4762
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8312 3670 8340 4082
rect 8404 4078 8432 4558
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8404 3942 8432 4014
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8300 3664 8352 3670
rect 8300 3606 8352 3612
rect 8496 3534 8524 7686
rect 8588 5370 8616 12406
rect 9140 11898 9168 12786
rect 9416 12238 9444 13874
rect 9772 13864 9824 13870
rect 9772 13806 9824 13812
rect 9784 12374 9812 13806
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8680 11354 8708 11630
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 9926 9352 10406
rect 9600 10130 9628 10542
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9128 9920 9180 9926
rect 9312 9920 9364 9926
rect 9128 9862 9180 9868
rect 9310 9888 9312 9897
rect 9680 9920 9732 9926
rect 9364 9888 9366 9897
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8956 9178 8984 9522
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9140 8974 9168 9862
rect 9680 9862 9732 9868
rect 9310 9823 9366 9832
rect 9692 9722 9720 9862
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8680 5234 8708 6666
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 6322 8892 6598
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8772 5545 8800 6258
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8758 5536 8814 5545
rect 8758 5471 8814 5480
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8404 3074 8432 3402
rect 8312 3046 8432 3074
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8208 1760 8260 1766
rect 8208 1702 8260 1708
rect 8220 800 8248 1702
rect 8312 800 8340 3046
rect 8390 2952 8446 2961
rect 8390 2887 8446 2896
rect 8404 800 8432 2887
rect 8496 800 8524 3470
rect 8588 3058 8616 3878
rect 8680 3738 8708 5170
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8864 3942 8892 4490
rect 8956 4146 8984 4626
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 9140 3738 9168 5646
rect 9232 4554 9260 8230
rect 9968 8090 9996 15302
rect 10060 13954 10088 15846
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10152 14074 10180 14282
rect 10244 14074 10272 14350
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10060 13926 10180 13954
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 9654 10088 12174
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9324 4690 9352 6054
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9310 4040 9366 4049
rect 9310 3975 9312 3984
rect 9364 3975 9366 3984
rect 9312 3946 9364 3952
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8680 2854 8708 3538
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8850 3224 8906 3233
rect 8850 3159 8906 3168
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8588 800 8616 2586
rect 8772 800 8800 3062
rect 8864 3058 8892 3159
rect 8852 3052 8904 3058
rect 8852 2994 8904 3000
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8864 800 8892 2858
rect 9048 800 9076 3470
rect 9140 2990 9168 3674
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 9232 2774 9260 3878
rect 9416 3126 9444 7142
rect 9508 6934 9536 7822
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9508 5817 9536 6734
rect 9494 5808 9550 5817
rect 9494 5743 9550 5752
rect 9494 5536 9550 5545
rect 9494 5471 9550 5480
rect 9508 3602 9536 5471
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9494 3088 9550 3097
rect 9494 3023 9496 3032
rect 9548 3023 9550 3032
rect 9496 2994 9548 3000
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9140 2746 9260 2774
rect 9140 800 9168 2746
rect 9324 800 9352 2926
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9416 2446 9444 2518
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9508 2378 9536 2450
rect 9600 2378 9628 7142
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 2774 9720 5646
rect 9784 3738 9812 5850
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9876 5030 9904 5578
rect 10060 5098 10088 5646
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 10060 4758 10088 5034
rect 10152 4826 10180 13926
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10336 9042 10364 9454
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10428 8362 10456 16068
rect 10612 15502 10640 16390
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10704 13530 10732 17206
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10796 16658 10824 17002
rect 10784 16652 10836 16658
rect 10784 16594 10836 16600
rect 10796 16454 10824 16594
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10888 16250 10916 26862
rect 10980 25294 11008 27610
rect 11072 26586 11100 30534
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 11164 29034 11192 29582
rect 11716 29170 11744 31146
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11428 29096 11480 29102
rect 11428 29038 11480 29044
rect 11152 29028 11204 29034
rect 11152 28970 11204 28976
rect 11440 28558 11468 29038
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11060 26580 11112 26586
rect 11060 26522 11112 26528
rect 11072 25362 11100 26522
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10980 24818 11008 25230
rect 11060 25152 11112 25158
rect 11060 25094 11112 25100
rect 11072 24886 11100 25094
rect 11060 24880 11112 24886
rect 11060 24822 11112 24828
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11072 24206 11100 24550
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 11334 24168 11390 24177
rect 11072 22001 11100 24142
rect 11152 24132 11204 24138
rect 11334 24103 11336 24112
rect 11152 24074 11204 24080
rect 11388 24103 11390 24112
rect 11336 24074 11388 24080
rect 11164 23866 11192 24074
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 11244 22976 11296 22982
rect 11244 22918 11296 22924
rect 11058 21992 11114 22001
rect 11058 21927 11114 21936
rect 11152 20868 11204 20874
rect 11152 20810 11204 20816
rect 11164 20602 11192 20810
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 10980 18086 11008 19382
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 16522 11008 18022
rect 10968 16516 11020 16522
rect 10968 16458 11020 16464
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 11072 16046 11100 18566
rect 11060 16040 11112 16046
rect 11060 15982 11112 15988
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 10888 14414 10916 15506
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12442 10548 13194
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10980 11762 11008 12582
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 10784 9512 10836 9518
rect 10784 9454 10836 9460
rect 10796 9042 10824 9454
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10980 6882 11008 11698
rect 11072 10266 11100 12038
rect 11164 11286 11192 19994
rect 11256 16590 11284 22918
rect 11336 21344 11388 21350
rect 11336 21286 11388 21292
rect 11348 20534 11376 21286
rect 11336 20528 11388 20534
rect 11336 20470 11388 20476
rect 11348 17610 11376 20470
rect 11440 17882 11468 28494
rect 11716 27946 11744 29106
rect 11888 29028 11940 29034
rect 11888 28970 11940 28976
rect 11704 27940 11756 27946
rect 11704 27882 11756 27888
rect 11716 27606 11744 27882
rect 11704 27600 11756 27606
rect 11704 27542 11756 27548
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11716 25906 11744 26318
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11624 23118 11652 23802
rect 11808 23798 11836 24006
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11612 23112 11664 23118
rect 11716 23089 11744 23666
rect 11796 23112 11848 23118
rect 11612 23054 11664 23060
rect 11702 23080 11758 23089
rect 11796 23054 11848 23060
rect 11702 23015 11704 23024
rect 11756 23015 11758 23024
rect 11704 22986 11756 22992
rect 11520 22636 11572 22642
rect 11520 22578 11572 22584
rect 11532 19378 11560 22578
rect 11612 21412 11664 21418
rect 11612 21354 11664 21360
rect 11624 20942 11652 21354
rect 11808 21146 11836 23054
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 11612 20936 11664 20942
rect 11612 20878 11664 20884
rect 11624 20058 11652 20878
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 18358 11560 19110
rect 11808 18630 11836 19314
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11716 17610 11744 18022
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11900 17270 11928 28970
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 11992 27402 12020 27814
rect 11980 27396 12032 27402
rect 11980 27338 12032 27344
rect 11888 17264 11940 17270
rect 11888 17206 11940 17212
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11348 16114 11376 17138
rect 11612 16516 11664 16522
rect 11612 16458 11664 16464
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11256 12322 11284 15642
rect 11348 12434 11376 16050
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11532 14346 11560 15370
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11624 13802 11652 16458
rect 11716 15910 11744 17138
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11808 16590 11836 17070
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11888 16516 11940 16522
rect 11888 16458 11940 16464
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11348 12406 11560 12434
rect 11256 12294 11376 12322
rect 11348 12050 11376 12294
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11440 12102 11468 12174
rect 11256 12022 11376 12050
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11072 7546 11100 10202
rect 11256 9058 11284 12022
rect 11532 11914 11560 12406
rect 11164 9030 11284 9058
rect 11348 11886 11560 11914
rect 11164 8838 11192 9030
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11164 7750 11192 7890
rect 11256 7818 11284 8774
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11152 7744 11204 7750
rect 11152 7686 11204 7692
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 10980 6854 11192 6882
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10048 4752 10100 4758
rect 10048 4694 10100 4700
rect 10060 4078 10088 4694
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9692 2746 9996 2774
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9496 2372 9548 2378
rect 9496 2314 9548 2320
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9416 800 9444 2246
rect 9600 800 9628 2314
rect 9692 800 9720 2518
rect 9862 2408 9918 2417
rect 9862 2343 9918 2352
rect 9876 2310 9904 2343
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9968 800 9996 2746
rect 10244 800 10272 5578
rect 10336 3534 10364 6054
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10428 5166 10456 5782
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 10428 4622 10456 4966
rect 10416 4616 10468 4622
rect 10416 4558 10468 4564
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10414 3224 10470 3233
rect 10414 3159 10470 3168
rect 10428 3126 10456 3159
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10520 800 10548 6054
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 5166 10640 5714
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10612 4758 10640 4966
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10796 800 10824 5170
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10888 4690 10916 5102
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10966 3768 11022 3777
rect 10966 3703 10968 3712
rect 11020 3703 11022 3712
rect 10968 3674 11020 3680
rect 10966 3224 11022 3233
rect 10966 3159 11022 3168
rect 10980 3126 11008 3159
rect 10968 3120 11020 3126
rect 10968 3062 11020 3068
rect 11072 800 11100 5102
rect 11164 3534 11192 6854
rect 11256 6798 11284 7278
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11348 5794 11376 11886
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 11082 11560 11698
rect 11520 11076 11572 11082
rect 11520 11018 11572 11024
rect 11612 11008 11664 11014
rect 11612 10950 11664 10956
rect 11624 10674 11652 10950
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11612 8016 11664 8022
rect 11612 7958 11664 7964
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 11532 6730 11560 7686
rect 11624 7585 11652 7958
rect 11610 7576 11666 7585
rect 11610 7511 11666 7520
rect 11624 7478 11652 7511
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11256 5766 11376 5794
rect 11256 4049 11284 5766
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11242 4040 11298 4049
rect 11242 3975 11298 3984
rect 11244 3664 11296 3670
rect 11244 3606 11296 3612
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11152 3392 11204 3398
rect 11256 3380 11284 3606
rect 11204 3352 11284 3380
rect 11152 3334 11204 3340
rect 11348 800 11376 5646
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11532 4622 11560 4762
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11624 4146 11652 6054
rect 11716 5302 11744 15846
rect 11808 12986 11836 16118
rect 11900 15366 11928 16458
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11888 15360 11940 15366
rect 11888 15302 11940 15308
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11808 12238 11836 12922
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11900 9092 11928 15302
rect 11808 9064 11928 9092
rect 11808 8498 11836 9064
rect 11992 9024 12020 16186
rect 12084 15706 12112 34546
rect 12452 32824 12480 34954
rect 12532 34400 12584 34406
rect 12532 34342 12584 34348
rect 12544 34202 12572 34342
rect 12532 34196 12584 34202
rect 12532 34138 12584 34144
rect 12532 32836 12584 32842
rect 12452 32796 12532 32824
rect 12532 32778 12584 32784
rect 12624 32836 12676 32842
rect 12728 32824 12756 36790
rect 12820 36786 12848 37742
rect 12808 36780 12860 36786
rect 12808 36722 12860 36728
rect 12820 35086 12848 36722
rect 13084 36644 13136 36650
rect 13084 36586 13136 36592
rect 12900 36576 12952 36582
rect 12900 36518 12952 36524
rect 12912 35698 12940 36518
rect 13096 36378 13124 36586
rect 13084 36372 13136 36378
rect 13084 36314 13136 36320
rect 12900 35692 12952 35698
rect 12900 35634 12952 35640
rect 12808 35080 12860 35086
rect 12808 35022 12860 35028
rect 12820 32978 12848 35022
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 12808 32972 12860 32978
rect 12808 32914 12860 32920
rect 12676 32796 12756 32824
rect 12624 32778 12676 32784
rect 12256 31136 12308 31142
rect 12256 31078 12308 31084
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 12268 30666 12296 31078
rect 12256 30660 12308 30666
rect 12256 30602 12308 30608
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 12176 28626 12204 30194
rect 12164 28620 12216 28626
rect 12164 28562 12216 28568
rect 12164 27396 12216 27402
rect 12164 27338 12216 27344
rect 12176 25362 12204 27338
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 12164 25152 12216 25158
rect 12164 25094 12216 25100
rect 12176 24070 12204 25094
rect 12164 24064 12216 24070
rect 12164 24006 12216 24012
rect 12164 23248 12216 23254
rect 12164 23190 12216 23196
rect 12176 23050 12204 23190
rect 12164 23044 12216 23050
rect 12164 22986 12216 22992
rect 12268 22574 12296 30602
rect 12452 30190 12480 31078
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 12452 29034 12480 30126
rect 12544 29714 12572 32778
rect 12636 30648 12664 32778
rect 12716 32428 12768 32434
rect 12716 32370 12768 32376
rect 12728 32026 12756 32370
rect 12716 32020 12768 32026
rect 12716 31962 12768 31968
rect 12716 31816 12768 31822
rect 12716 31758 12768 31764
rect 12728 31414 12756 31758
rect 12716 31408 12768 31414
rect 12716 31350 12768 31356
rect 12716 30660 12768 30666
rect 12636 30620 12716 30648
rect 12636 30326 12664 30620
rect 12716 30602 12768 30608
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 12532 29708 12584 29714
rect 12532 29650 12584 29656
rect 12820 29646 12848 32914
rect 12992 32904 13044 32910
rect 12992 32846 13044 32852
rect 13004 32434 13032 32846
rect 13084 32768 13136 32774
rect 13084 32710 13136 32716
rect 12992 32428 13044 32434
rect 12992 32370 13044 32376
rect 12992 31816 13044 31822
rect 13096 31804 13124 32710
rect 13188 31822 13216 34478
rect 13044 31776 13124 31804
rect 13176 31816 13228 31822
rect 12992 31758 13044 31764
rect 13176 31758 13228 31764
rect 13188 31482 13216 31758
rect 13280 31686 13308 38490
rect 13360 38208 13412 38214
rect 13360 38150 13412 38156
rect 13372 37874 13400 38150
rect 13360 37868 13412 37874
rect 13360 37810 13412 37816
rect 13452 37868 13504 37874
rect 13452 37810 13504 37816
rect 13464 36854 13492 37810
rect 13556 37806 13584 38490
rect 13636 38480 13688 38486
rect 13636 38422 13688 38428
rect 13648 37874 13676 38422
rect 13832 38282 13860 40870
rect 14936 40526 14964 41074
rect 14924 40520 14976 40526
rect 14924 40462 14976 40468
rect 14372 39296 14424 39302
rect 14372 39238 14424 39244
rect 13820 38276 13872 38282
rect 13820 38218 13872 38224
rect 13636 37868 13688 37874
rect 13636 37810 13688 37816
rect 14004 37868 14056 37874
rect 14004 37810 14056 37816
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13452 36848 13504 36854
rect 13452 36790 13504 36796
rect 13464 36378 13492 36790
rect 13648 36530 13676 37810
rect 14016 37754 14044 37810
rect 13924 37738 14044 37754
rect 14096 37800 14148 37806
rect 14096 37742 14148 37748
rect 13912 37732 14044 37738
rect 13964 37726 14044 37732
rect 13912 37674 13964 37680
rect 14108 37330 14136 37742
rect 14096 37324 14148 37330
rect 14096 37266 14148 37272
rect 14096 37188 14148 37194
rect 14096 37130 14148 37136
rect 13648 36502 13768 36530
rect 13452 36372 13504 36378
rect 13452 36314 13504 36320
rect 13740 34134 13768 36502
rect 14108 36378 14136 37130
rect 14096 36372 14148 36378
rect 14096 36314 14148 36320
rect 14384 36174 14412 39238
rect 14936 37806 14964 40462
rect 15396 38418 15424 41754
rect 15488 41614 15516 42026
rect 15764 41682 15792 42162
rect 15752 41676 15804 41682
rect 15752 41618 15804 41624
rect 15476 41608 15528 41614
rect 15476 41550 15528 41556
rect 15488 41070 15516 41550
rect 15764 41274 15792 41618
rect 15752 41268 15804 41274
rect 15752 41210 15804 41216
rect 15948 41138 15976 42502
rect 16120 42016 16172 42022
rect 16120 41958 16172 41964
rect 16132 41614 16160 41958
rect 16120 41608 16172 41614
rect 16120 41550 16172 41556
rect 15936 41132 15988 41138
rect 15936 41074 15988 41080
rect 16120 41132 16172 41138
rect 16120 41074 16172 41080
rect 15476 41064 15528 41070
rect 15476 41006 15528 41012
rect 16132 41002 16160 41074
rect 16120 40996 16172 41002
rect 16120 40938 16172 40944
rect 15476 40928 15528 40934
rect 15476 40870 15528 40876
rect 15488 40458 15516 40870
rect 15476 40452 15528 40458
rect 15476 40394 15528 40400
rect 16316 40390 16344 42570
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19892 42152 19944 42158
rect 19892 42094 19944 42100
rect 19524 42016 19576 42022
rect 19524 41958 19576 41964
rect 19536 41614 19564 41958
rect 19904 41614 19932 42094
rect 20352 41812 20404 41818
rect 20352 41754 20404 41760
rect 16856 41608 16908 41614
rect 16856 41550 16908 41556
rect 18696 41608 18748 41614
rect 18696 41550 18748 41556
rect 19524 41608 19576 41614
rect 19524 41550 19576 41556
rect 19892 41608 19944 41614
rect 19944 41568 20024 41596
rect 19892 41550 19944 41556
rect 16868 40526 16896 41550
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 17972 41274 18000 41414
rect 17960 41268 18012 41274
rect 17960 41210 18012 41216
rect 17972 41138 18000 41210
rect 17960 41132 18012 41138
rect 17960 41074 18012 41080
rect 18420 41064 18472 41070
rect 18420 41006 18472 41012
rect 17960 40996 18012 41002
rect 17960 40938 18012 40944
rect 16856 40520 16908 40526
rect 16856 40462 16908 40468
rect 15568 40384 15620 40390
rect 15568 40326 15620 40332
rect 16304 40384 16356 40390
rect 16304 40326 16356 40332
rect 15384 38412 15436 38418
rect 15384 38354 15436 38360
rect 15108 38276 15160 38282
rect 15108 38218 15160 38224
rect 15120 38010 15148 38218
rect 15476 38208 15528 38214
rect 15476 38150 15528 38156
rect 15108 38004 15160 38010
rect 15108 37946 15160 37952
rect 15488 37874 15516 38150
rect 15580 37942 15608 40326
rect 16672 39840 16724 39846
rect 16672 39782 16724 39788
rect 16684 38962 16712 39782
rect 17972 39302 18000 40938
rect 18432 40050 18460 41006
rect 18708 40934 18736 41550
rect 18972 41540 19024 41546
rect 18972 41482 19024 41488
rect 19340 41540 19392 41546
rect 19340 41482 19392 41488
rect 18604 40928 18656 40934
rect 18604 40870 18656 40876
rect 18696 40928 18748 40934
rect 18696 40870 18748 40876
rect 18616 40458 18644 40870
rect 18512 40452 18564 40458
rect 18512 40394 18564 40400
rect 18604 40452 18656 40458
rect 18604 40394 18656 40400
rect 18420 40044 18472 40050
rect 18420 39986 18472 39992
rect 18524 39846 18552 40394
rect 18512 39840 18564 39846
rect 18512 39782 18564 39788
rect 17960 39296 18012 39302
rect 17960 39238 18012 39244
rect 16672 38956 16724 38962
rect 16672 38898 16724 38904
rect 16396 38752 16448 38758
rect 16396 38694 16448 38700
rect 15844 38276 15896 38282
rect 15844 38218 15896 38224
rect 15568 37936 15620 37942
rect 15568 37878 15620 37884
rect 15476 37868 15528 37874
rect 15476 37810 15528 37816
rect 14924 37800 14976 37806
rect 14924 37742 14976 37748
rect 15200 37732 15252 37738
rect 15200 37674 15252 37680
rect 14464 37664 14516 37670
rect 14464 37606 14516 37612
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 13912 36100 13964 36106
rect 13912 36042 13964 36048
rect 13728 34128 13780 34134
rect 13728 34070 13780 34076
rect 13740 33998 13768 34070
rect 13728 33992 13780 33998
rect 13728 33934 13780 33940
rect 13924 33930 13952 36042
rect 14384 36038 14412 36110
rect 14372 36032 14424 36038
rect 14372 35974 14424 35980
rect 14188 33992 14240 33998
rect 14188 33934 14240 33940
rect 13912 33924 13964 33930
rect 13912 33866 13964 33872
rect 13924 32434 13952 33866
rect 14200 32434 14228 33934
rect 13912 32428 13964 32434
rect 13912 32370 13964 32376
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 13268 31680 13320 31686
rect 13268 31622 13320 31628
rect 13176 31476 13228 31482
rect 13176 31418 13228 31424
rect 12992 30592 13044 30598
rect 12992 30534 13044 30540
rect 13004 30258 13032 30534
rect 13188 30258 13216 31418
rect 13280 30394 13308 31622
rect 14200 31210 14228 32370
rect 14384 31686 14412 32370
rect 14372 31680 14424 31686
rect 14372 31622 14424 31628
rect 14384 31346 14412 31622
rect 14372 31340 14424 31346
rect 14372 31282 14424 31288
rect 14188 31204 14240 31210
rect 14188 31146 14240 31152
rect 13360 30660 13412 30666
rect 13360 30602 13412 30608
rect 13268 30388 13320 30394
rect 13268 30330 13320 30336
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 13176 30252 13228 30258
rect 13176 30194 13228 30200
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12912 29714 12940 29990
rect 13188 29850 13216 30194
rect 13176 29844 13228 29850
rect 13176 29786 13228 29792
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 12808 29640 12860 29646
rect 12808 29582 12860 29588
rect 12820 29170 12848 29582
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12440 29028 12492 29034
rect 12440 28970 12492 28976
rect 12912 28762 12940 29650
rect 13372 29578 13400 30602
rect 13728 30592 13780 30598
rect 13728 30534 13780 30540
rect 13740 30258 13768 30534
rect 13728 30252 13780 30258
rect 13728 30194 13780 30200
rect 13452 30184 13504 30190
rect 13452 30126 13504 30132
rect 13360 29572 13412 29578
rect 13360 29514 13412 29520
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12544 28014 12572 28154
rect 12532 28008 12584 28014
rect 12532 27950 12584 27956
rect 12912 27946 12940 28698
rect 13464 28422 13492 30126
rect 14372 30116 14424 30122
rect 14372 30058 14424 30064
rect 14384 28966 14412 30058
rect 14372 28960 14424 28966
rect 14372 28902 14424 28908
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13452 28416 13504 28422
rect 13452 28358 13504 28364
rect 13084 28144 13136 28150
rect 13084 28086 13136 28092
rect 12900 27940 12952 27946
rect 12900 27882 12952 27888
rect 12912 27614 12940 27882
rect 13096 27674 13124 28086
rect 13464 28082 13492 28358
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 12820 27586 12940 27614
rect 13084 27668 13136 27674
rect 13084 27610 13136 27616
rect 12348 27056 12400 27062
rect 12348 26998 12400 27004
rect 12360 26586 12388 26998
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12624 25220 12676 25226
rect 12624 25162 12676 25168
rect 12636 24954 12664 25162
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12728 24886 12756 25094
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12348 24200 12400 24206
rect 12346 24168 12348 24177
rect 12400 24168 12402 24177
rect 12346 24103 12402 24112
rect 12544 24070 12572 24346
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12636 23322 12664 24142
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 12256 22568 12308 22574
rect 12256 22510 12308 22516
rect 12820 21622 12848 27586
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13464 26382 13492 27406
rect 13740 26994 13768 28426
rect 13832 28218 13860 28698
rect 14384 28626 14412 28902
rect 14372 28620 14424 28626
rect 14372 28562 14424 28568
rect 14188 28416 14240 28422
rect 14188 28358 14240 28364
rect 14200 28218 14228 28358
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 13728 26988 13780 26994
rect 13728 26930 13780 26936
rect 14384 26450 14412 27950
rect 14372 26444 14424 26450
rect 14372 26386 14424 26392
rect 13452 26376 13504 26382
rect 13452 26318 13504 26324
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 12898 24848 12954 24857
rect 12898 24783 12900 24792
rect 12952 24783 12954 24792
rect 12900 24754 12952 24760
rect 12912 24682 12940 24754
rect 12900 24676 12952 24682
rect 12900 24618 12952 24624
rect 13004 24138 13032 25774
rect 13084 25696 13136 25702
rect 13084 25638 13136 25644
rect 13096 24818 13124 25638
rect 13084 24812 13136 24818
rect 13084 24754 13136 24760
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 13280 24342 13308 24754
rect 13268 24336 13320 24342
rect 13268 24278 13320 24284
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23798 13032 24074
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12176 21350 12204 21558
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12164 21344 12216 21350
rect 12162 21312 12164 21321
rect 12216 21312 12218 21321
rect 12162 21247 12218 21256
rect 12820 20641 12848 21354
rect 12806 20632 12862 20641
rect 12806 20567 12862 20576
rect 12820 20534 12848 20567
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12176 19378 12204 19994
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12268 19446 12296 19858
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12452 18698 12480 19654
rect 12820 19378 12848 20266
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 12912 19514 12940 19790
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12268 17610 12296 18362
rect 12256 17604 12308 17610
rect 12256 17546 12308 17552
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12176 16046 12204 16526
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 12084 13326 12112 13738
rect 12268 13462 12296 17546
rect 12728 16794 12756 17546
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12716 16448 12768 16454
rect 12716 16390 12768 16396
rect 12728 16114 12756 16390
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12452 14822 12480 16050
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12268 12170 12296 13398
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12360 12102 12388 13126
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12176 9722 12204 9930
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 11900 8996 12020 9024
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11808 5846 11836 8434
rect 11900 5914 11928 8996
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 11992 8294 12020 8842
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11992 6118 12020 7822
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 12084 5681 12112 8842
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12176 7274 12204 7482
rect 12164 7268 12216 7274
rect 12164 7210 12216 7216
rect 12070 5672 12126 5681
rect 12070 5607 12126 5616
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 11808 4826 11836 4966
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11520 2576 11572 2582
rect 11518 2544 11520 2553
rect 11572 2544 11574 2553
rect 11518 2479 11574 2488
rect 11532 2038 11560 2479
rect 11520 2032 11572 2038
rect 11520 1974 11572 1980
rect 11624 800 11652 3878
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11716 2446 11744 2926
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11900 800 11928 4966
rect 12084 3194 12112 4966
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12176 800 12204 3878
rect 12268 3670 12296 4626
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12360 2774 12388 12038
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12452 10810 12480 11086
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12452 9586 12480 10406
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12544 9110 12572 10542
rect 12636 10130 12664 11086
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12728 10577 12756 10610
rect 12714 10568 12770 10577
rect 12714 10503 12770 10512
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12820 9194 12848 14758
rect 13004 12102 13032 23734
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13176 21004 13228 21010
rect 13176 20946 13228 20952
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 13096 20058 13124 20470
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13096 19854 13124 19994
rect 13188 19922 13216 20946
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13096 18970 13124 19314
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13280 17270 13308 20402
rect 13372 19990 13400 21286
rect 13360 19984 13412 19990
rect 13360 19926 13412 19932
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13188 14618 13216 17138
rect 13280 16114 13308 17206
rect 13372 17202 13400 18906
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13464 16794 13492 26318
rect 14372 26036 14424 26042
rect 14372 25978 14424 25984
rect 13912 25968 13964 25974
rect 13912 25910 13964 25916
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13832 23730 13860 25230
rect 13924 25158 13952 25910
rect 14280 25900 14332 25906
rect 14280 25842 14332 25848
rect 14292 25158 14320 25842
rect 13912 25152 13964 25158
rect 13912 25094 13964 25100
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 13924 24070 13952 25094
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14200 24614 14228 24754
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 14108 23866 14136 24074
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13832 22098 13860 23666
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 13912 22500 13964 22506
rect 13912 22442 13964 22448
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 13924 21554 13952 22442
rect 14108 21706 14136 23462
rect 14200 23050 14228 24550
rect 14188 23044 14240 23050
rect 14188 22986 14240 22992
rect 14016 21678 14136 21706
rect 14292 21690 14320 25094
rect 14384 24206 14412 25978
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23798 14412 24006
rect 14372 23792 14424 23798
rect 14372 23734 14424 23740
rect 14280 21684 14332 21690
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 13924 20534 13952 21490
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13832 19378 13860 19722
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13556 17746 13584 18702
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13556 15570 13584 17682
rect 14016 17202 14044 21678
rect 14280 21626 14332 21632
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14108 21146 14136 21490
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14200 21010 14228 21490
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20602 14136 20878
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14200 20058 14228 20402
rect 14476 20262 14504 37606
rect 14832 36780 14884 36786
rect 14832 36722 14884 36728
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14568 36174 14596 36518
rect 14648 36236 14700 36242
rect 14648 36178 14700 36184
rect 14556 36168 14608 36174
rect 14556 36110 14608 36116
rect 14660 35630 14688 36178
rect 14648 35624 14700 35630
rect 14648 35566 14700 35572
rect 14660 34066 14688 35566
rect 14648 34060 14700 34066
rect 14648 34002 14700 34008
rect 14844 33658 14872 36722
rect 14832 33652 14884 33658
rect 14832 33594 14884 33600
rect 15212 33590 15240 37674
rect 15856 37466 15884 38218
rect 15844 37460 15896 37466
rect 15844 37402 15896 37408
rect 15856 36854 15884 37402
rect 16212 37120 16264 37126
rect 16212 37062 16264 37068
rect 15844 36848 15896 36854
rect 15844 36790 15896 36796
rect 16224 36174 16252 37062
rect 16408 36174 16436 38694
rect 18708 38486 18736 40870
rect 18788 40384 18840 40390
rect 18788 40326 18840 40332
rect 18800 40118 18828 40326
rect 18788 40112 18840 40118
rect 18788 40054 18840 40060
rect 17408 38480 17460 38486
rect 17408 38422 17460 38428
rect 18696 38480 18748 38486
rect 18696 38422 18748 38428
rect 17420 38282 17448 38422
rect 18328 38412 18380 38418
rect 18328 38354 18380 38360
rect 17408 38276 17460 38282
rect 17408 38218 17460 38224
rect 16488 38208 16540 38214
rect 16488 38150 16540 38156
rect 16500 37738 16528 38150
rect 16764 37868 16816 37874
rect 16764 37810 16816 37816
rect 16488 37732 16540 37738
rect 16488 37674 16540 37680
rect 16672 36712 16724 36718
rect 16672 36654 16724 36660
rect 16684 36242 16712 36654
rect 16776 36378 16804 37810
rect 18340 37738 18368 38354
rect 18604 38276 18656 38282
rect 18604 38218 18656 38224
rect 18512 38208 18564 38214
rect 18512 38150 18564 38156
rect 18328 37732 18380 37738
rect 18328 37674 18380 37680
rect 17960 37664 18012 37670
rect 17960 37606 18012 37612
rect 17972 37330 18000 37606
rect 17960 37324 18012 37330
rect 17960 37266 18012 37272
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 16948 37188 17000 37194
rect 16948 37130 17000 37136
rect 16960 36786 16988 37130
rect 18064 36922 18092 37198
rect 18340 37194 18368 37674
rect 18328 37188 18380 37194
rect 18328 37130 18380 37136
rect 18052 36916 18104 36922
rect 18052 36858 18104 36864
rect 16948 36780 17000 36786
rect 16948 36722 17000 36728
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 17316 36780 17368 36786
rect 17316 36722 17368 36728
rect 16960 36394 16988 36722
rect 16764 36372 16816 36378
rect 16960 36366 17080 36394
rect 16764 36314 16816 36320
rect 16672 36236 16724 36242
rect 16672 36178 16724 36184
rect 16212 36168 16264 36174
rect 16212 36110 16264 36116
rect 16396 36168 16448 36174
rect 16448 36128 16620 36156
rect 16396 36110 16448 36116
rect 15568 36032 15620 36038
rect 15568 35974 15620 35980
rect 15200 33584 15252 33590
rect 15200 33526 15252 33532
rect 15016 33516 15068 33522
rect 15016 33458 15068 33464
rect 14556 32836 14608 32842
rect 14556 32778 14608 32784
rect 14568 32502 14596 32778
rect 15028 32502 15056 33458
rect 15580 32774 15608 35974
rect 16592 35834 16620 36128
rect 16580 35828 16632 35834
rect 16580 35770 16632 35776
rect 16684 35018 16712 36178
rect 17052 36174 17080 36366
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 17144 36106 17172 36722
rect 17328 36378 17356 36722
rect 17316 36372 17368 36378
rect 17316 36314 17368 36320
rect 17132 36100 17184 36106
rect 17132 36042 17184 36048
rect 17684 36100 17736 36106
rect 17684 36042 17736 36048
rect 16856 35488 16908 35494
rect 16856 35430 16908 35436
rect 16868 35086 16896 35430
rect 17144 35086 17172 36042
rect 17224 35284 17276 35290
rect 17224 35226 17276 35232
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 16672 35012 16724 35018
rect 16672 34954 16724 34960
rect 16764 34944 16816 34950
rect 16764 34886 16816 34892
rect 16776 34610 16804 34886
rect 16764 34604 16816 34610
rect 16764 34546 16816 34552
rect 16868 34134 16896 35022
rect 17236 34746 17264 35226
rect 17316 35216 17368 35222
rect 17316 35158 17368 35164
rect 17224 34740 17276 34746
rect 17224 34682 17276 34688
rect 16856 34128 16908 34134
rect 16856 34070 16908 34076
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 15108 32768 15160 32774
rect 15108 32710 15160 32716
rect 15476 32768 15528 32774
rect 15476 32710 15528 32716
rect 15568 32768 15620 32774
rect 15568 32710 15620 32716
rect 14556 32496 14608 32502
rect 14556 32438 14608 32444
rect 15016 32496 15068 32502
rect 15016 32438 15068 32444
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14660 25974 14688 29106
rect 14752 28082 14780 29446
rect 14844 29170 14872 29990
rect 15028 29782 15056 32438
rect 15120 32434 15148 32710
rect 15488 32502 15516 32710
rect 15476 32496 15528 32502
rect 15476 32438 15528 32444
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 16132 31890 16160 32846
rect 16592 32366 16620 33866
rect 16868 33046 16896 34070
rect 17328 33998 17356 35158
rect 17696 35086 17724 36042
rect 17684 35080 17736 35086
rect 17684 35022 17736 35028
rect 17868 35012 17920 35018
rect 17868 34954 17920 34960
rect 17880 34746 17908 34954
rect 17500 34740 17552 34746
rect 17500 34682 17552 34688
rect 17868 34740 17920 34746
rect 17868 34682 17920 34688
rect 17512 33998 17540 34682
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17500 33992 17552 33998
rect 17500 33934 17552 33940
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17788 33590 17816 33934
rect 16948 33584 17000 33590
rect 16948 33526 17000 33532
rect 17776 33584 17828 33590
rect 17776 33526 17828 33532
rect 16856 33040 16908 33046
rect 16856 32982 16908 32988
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16132 30802 16160 31826
rect 16592 31754 16620 32302
rect 16960 32298 16988 33526
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 16948 32292 17000 32298
rect 16948 32234 17000 32240
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 16776 31822 16804 31962
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16580 31748 16632 31754
rect 16580 31690 16632 31696
rect 16684 31482 16712 31758
rect 16672 31476 16724 31482
rect 16672 31418 16724 31424
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 15200 30660 15252 30666
rect 15200 30602 15252 30608
rect 15844 30660 15896 30666
rect 15844 30602 15896 30608
rect 15212 30326 15240 30602
rect 15856 30394 15884 30602
rect 15844 30388 15896 30394
rect 15844 30330 15896 30336
rect 16776 30326 16804 31758
rect 16856 31748 16908 31754
rect 16856 31690 16908 31696
rect 15200 30320 15252 30326
rect 15200 30262 15252 30268
rect 16764 30320 16816 30326
rect 16764 30262 16816 30268
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15016 29776 15068 29782
rect 15016 29718 15068 29724
rect 14832 29164 14884 29170
rect 14832 29106 14884 29112
rect 15028 28762 15056 29718
rect 15108 29096 15160 29102
rect 15108 29038 15160 29044
rect 15016 28756 15068 28762
rect 15016 28698 15068 28704
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 14832 28552 14884 28558
rect 14832 28494 14884 28500
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14844 27402 14872 28494
rect 14832 27396 14884 27402
rect 14832 27338 14884 27344
rect 14844 27062 14872 27338
rect 14832 27056 14884 27062
rect 14832 26998 14884 27004
rect 14648 25968 14700 25974
rect 14648 25910 14700 25916
rect 14740 25220 14792 25226
rect 14740 25162 14792 25168
rect 14752 24954 14780 25162
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14740 24064 14792 24070
rect 14740 24006 14792 24012
rect 14752 23866 14780 24006
rect 14740 23860 14792 23866
rect 14740 23802 14792 23808
rect 14648 22228 14700 22234
rect 14648 22170 14700 22176
rect 14660 22094 14688 22170
rect 14660 22066 14780 22094
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14568 21690 14596 21898
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 14752 20466 14780 22066
rect 14936 21486 14964 28562
rect 15016 28484 15068 28490
rect 15016 28426 15068 28432
rect 15028 28082 15056 28426
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 15120 27946 15148 29038
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15212 28150 15240 28358
rect 15200 28144 15252 28150
rect 15200 28086 15252 28092
rect 15304 28082 15332 30194
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 15752 29776 15804 29782
rect 15752 29718 15804 29724
rect 15764 29170 15792 29718
rect 15936 29572 15988 29578
rect 15936 29514 15988 29520
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 15488 28558 15516 28902
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15948 28422 15976 29514
rect 16684 29510 16712 30126
rect 16776 29646 16804 30262
rect 16764 29640 16816 29646
rect 16764 29582 16816 29588
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16672 29504 16724 29510
rect 16672 29446 16724 29452
rect 16040 29170 16068 29446
rect 16028 29164 16080 29170
rect 16028 29106 16080 29112
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 15936 28416 15988 28422
rect 15936 28358 15988 28364
rect 16132 28150 16160 29106
rect 16212 28688 16264 28694
rect 16212 28630 16264 28636
rect 16224 28218 16252 28630
rect 16212 28212 16264 28218
rect 16212 28154 16264 28160
rect 16120 28144 16172 28150
rect 16120 28086 16172 28092
rect 15292 28076 15344 28082
rect 15292 28018 15344 28024
rect 15108 27940 15160 27946
rect 15108 27882 15160 27888
rect 15304 27538 15332 28018
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15292 27532 15344 27538
rect 15292 27474 15344 27480
rect 15396 27418 15424 27814
rect 16132 27674 16160 28086
rect 16120 27668 16172 27674
rect 16120 27610 16172 27616
rect 16224 27554 16252 28154
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 15304 27390 15424 27418
rect 16132 27526 16252 27554
rect 15016 27328 15068 27334
rect 15016 27270 15068 27276
rect 15028 25974 15056 27270
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15016 25968 15068 25974
rect 15016 25910 15068 25916
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 15028 24070 15056 24346
rect 15016 24064 15068 24070
rect 15016 24006 15068 24012
rect 15016 23656 15068 23662
rect 15016 23598 15068 23604
rect 15028 23322 15056 23598
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14740 20460 14792 20466
rect 14740 20402 14792 20408
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14464 20256 14516 20262
rect 14464 20198 14516 20204
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 13648 16697 13676 16934
rect 14108 16726 14136 16934
rect 14096 16720 14148 16726
rect 13634 16688 13690 16697
rect 14096 16662 14148 16668
rect 13634 16623 13690 16632
rect 13648 16590 13676 16623
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13740 16046 13768 16390
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13556 14482 13584 15506
rect 14200 15162 14228 15914
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 14292 14006 14320 20198
rect 15120 20058 15148 26250
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15212 24410 15240 24754
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15304 24138 15332 27390
rect 16132 27130 16160 27526
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 16132 26994 16160 27066
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 15948 26518 15976 26930
rect 15936 26512 15988 26518
rect 15936 26454 15988 26460
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15580 24954 15608 25638
rect 15568 24948 15620 24954
rect 15568 24890 15620 24896
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15396 24410 15424 24754
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15476 24200 15528 24206
rect 15476 24142 15528 24148
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 15488 23798 15516 24142
rect 15672 24138 15700 25638
rect 15660 24132 15712 24138
rect 15660 24074 15712 24080
rect 15476 23792 15528 23798
rect 15476 23734 15528 23740
rect 15660 23792 15712 23798
rect 15660 23734 15712 23740
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 15212 23254 15240 23666
rect 15672 23610 15700 23734
rect 15304 23582 15700 23610
rect 15200 23248 15252 23254
rect 15200 23190 15252 23196
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15212 21554 15240 22714
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15212 18737 15240 21490
rect 15304 20874 15332 23582
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15488 23118 15516 23462
rect 15948 23254 15976 26454
rect 16120 26376 16172 26382
rect 16120 26318 16172 26324
rect 16028 24948 16080 24954
rect 16028 24890 16080 24896
rect 15936 23248 15988 23254
rect 15936 23190 15988 23196
rect 15476 23112 15528 23118
rect 15476 23054 15528 23060
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15672 22234 15700 23054
rect 15844 23044 15896 23050
rect 15844 22986 15896 22992
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 15672 20942 15700 22170
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15764 20942 15792 21286
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15292 20868 15344 20874
rect 15292 20810 15344 20816
rect 15764 20330 15792 20878
rect 15752 20324 15804 20330
rect 15752 20266 15804 20272
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15198 18728 15254 18737
rect 15198 18663 15254 18672
rect 15212 16590 15240 18663
rect 15304 16658 15332 19722
rect 15580 19514 15608 19790
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15396 18766 15424 19110
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15580 18358 15608 19314
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15200 16584 15252 16590
rect 15200 16526 15252 16532
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14568 16114 14596 16458
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14384 15502 14412 15846
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14844 15162 14872 16050
rect 15396 15978 15424 16186
rect 15384 15972 15436 15978
rect 15384 15914 15436 15920
rect 15292 15360 15344 15366
rect 15292 15302 15344 15308
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 15304 15026 15332 15302
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15304 14346 15332 14962
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13544 13252 13596 13258
rect 13544 13194 13596 13200
rect 13280 12986 13308 13194
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13280 12238 13308 12922
rect 13556 12889 13584 13194
rect 13542 12880 13598 12889
rect 13542 12815 13598 12824
rect 14016 12714 14044 13874
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 14108 12782 14136 13806
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12918 14228 13126
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14384 12850 14412 13670
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14669 13317 14721 13323
rect 14721 13280 14780 13308
rect 14669 13259 14721 13265
rect 14646 12880 14702 12889
rect 14372 12844 14424 12850
rect 14646 12815 14648 12824
rect 14372 12786 14424 12792
rect 14700 12815 14702 12824
rect 14648 12786 14700 12792
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 14108 12238 14136 12718
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 14096 12232 14148 12238
rect 14096 12174 14148 12180
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13004 11898 13032 12038
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 14108 11354 14136 12174
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13188 9382 13216 10678
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 12728 9166 12848 9194
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8430 12572 8774
rect 12532 8424 12584 8430
rect 12530 8392 12532 8401
rect 12584 8392 12586 8401
rect 12530 8327 12586 8336
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12452 7954 12480 8230
rect 12530 8120 12586 8129
rect 12530 8055 12586 8064
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12544 7886 12572 8055
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12636 6662 12664 7754
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12268 2746 12388 2774
rect 12268 2446 12296 2746
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12346 2408 12402 2417
rect 12346 2343 12402 2352
rect 12360 1970 12388 2343
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12452 800 12480 3878
rect 12636 3058 12664 6598
rect 12728 4826 12756 9166
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8634 12848 8978
rect 13188 8974 13216 9318
rect 13280 9178 13308 9998
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13372 8974 13400 9862
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13464 8974 13492 9590
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 13556 8498 13584 8774
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13266 8120 13322 8129
rect 13266 8055 13268 8064
rect 13320 8055 13322 8064
rect 13268 8026 13320 8032
rect 13924 7886 13952 8366
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 14384 7750 14412 12786
rect 14752 12238 14780 13280
rect 14936 13258 14964 13330
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12714 15240 13194
rect 15304 12850 15332 13262
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14648 12164 14700 12170
rect 14648 12106 14700 12112
rect 14660 11898 14688 12106
rect 15028 11898 15056 12650
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 14740 11688 14792 11694
rect 15120 11676 15148 12582
rect 15212 11830 15240 12650
rect 15200 11824 15252 11830
rect 15200 11766 15252 11772
rect 15304 11762 15332 12786
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15200 11688 15252 11694
rect 15120 11648 15200 11676
rect 14792 11636 15056 11642
rect 14740 11630 15056 11636
rect 15200 11630 15252 11636
rect 14752 11626 15056 11630
rect 14752 11620 15068 11626
rect 14752 11614 15016 11620
rect 15016 11562 15068 11568
rect 15304 11286 15332 11698
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 9382 14596 9522
rect 15396 9382 15424 13126
rect 15488 12918 15516 13466
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15488 12442 15516 12854
rect 15476 12436 15528 12442
rect 15476 12378 15528 12384
rect 15856 12102 15884 22986
rect 16040 19854 16068 24890
rect 16132 24886 16160 26318
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16120 24880 16172 24886
rect 16120 24822 16172 24828
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 23798 16160 24550
rect 16224 24206 16252 25094
rect 16316 24410 16344 28018
rect 16684 27554 16712 29446
rect 16868 28014 16896 31690
rect 16960 30258 16988 32234
rect 17144 31482 17172 33390
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17420 32298 17448 33050
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17500 32496 17552 32502
rect 17500 32438 17552 32444
rect 17408 32292 17460 32298
rect 17408 32234 17460 32240
rect 17512 32026 17540 32438
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17604 31754 17632 32846
rect 17776 32768 17828 32774
rect 17776 32710 17828 32716
rect 17788 32230 17816 32710
rect 17684 32224 17736 32230
rect 17684 32166 17736 32172
rect 17776 32224 17828 32230
rect 17776 32166 17828 32172
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17316 31680 17368 31686
rect 17316 31622 17368 31628
rect 17132 31476 17184 31482
rect 17132 31418 17184 31424
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 17144 29238 17172 31418
rect 17328 29238 17356 31622
rect 17408 31136 17460 31142
rect 17408 31078 17460 31084
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 17316 29232 17368 29238
rect 17316 29174 17368 29180
rect 17132 29028 17184 29034
rect 17132 28970 17184 28976
rect 17040 28552 17092 28558
rect 17040 28494 17092 28500
rect 16948 28212 17000 28218
rect 16948 28154 17000 28160
rect 16856 28008 16908 28014
rect 16856 27950 16908 27956
rect 16592 27526 16712 27554
rect 16592 26926 16620 27526
rect 16580 26920 16632 26926
rect 16580 26862 16632 26868
rect 16396 26784 16448 26790
rect 16396 26726 16448 26732
rect 16408 26450 16436 26726
rect 16396 26444 16448 26450
rect 16396 26386 16448 26392
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16212 24200 16264 24206
rect 16212 24142 16264 24148
rect 16120 23792 16172 23798
rect 16120 23734 16172 23740
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 16132 22642 16160 22918
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16120 22432 16172 22438
rect 16120 22374 16172 22380
rect 16132 21962 16160 22374
rect 16120 21956 16172 21962
rect 16120 21898 16172 21904
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19378 16068 19790
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 16132 18426 16160 21898
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16500 18766 16528 19246
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15948 16114 15976 16594
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16132 15434 16160 15846
rect 16120 15428 16172 15434
rect 16120 15370 16172 15376
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11898 16528 12038
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 12820 6390 12848 7686
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 13096 6322 13124 6734
rect 14476 6322 14504 7346
rect 14568 6730 14596 9318
rect 15580 9178 15608 11494
rect 16592 10130 16620 26862
rect 16960 26314 16988 28154
rect 17052 27402 17080 28494
rect 17144 28490 17172 28970
rect 17132 28484 17184 28490
rect 17132 28426 17184 28432
rect 17144 28218 17172 28426
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 16960 25430 16988 26250
rect 16948 25424 17000 25430
rect 16948 25366 17000 25372
rect 16960 22234 16988 25366
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 16960 21078 16988 21490
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16960 20874 16988 21014
rect 16948 20868 17000 20874
rect 16948 20810 17000 20816
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16684 18426 16712 19722
rect 16764 19440 16816 19446
rect 16764 19382 16816 19388
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16776 16182 16804 19382
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16854 18592 16910 18601
rect 16854 18527 16910 18536
rect 16868 18290 16896 18527
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16960 18154 16988 18906
rect 17052 18426 17080 27338
rect 17132 27124 17184 27130
rect 17132 27066 17184 27072
rect 17144 25906 17172 27066
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 17236 25498 17264 25842
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 17420 24614 17448 31078
rect 17592 29640 17644 29646
rect 17592 29582 17644 29588
rect 17604 28558 17632 29582
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 17408 24608 17460 24614
rect 17408 24550 17460 24556
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17420 24206 17448 24346
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17144 22386 17172 24006
rect 17512 23866 17540 24006
rect 17604 23866 17632 24142
rect 17500 23860 17552 23866
rect 17500 23802 17552 23808
rect 17592 23860 17644 23866
rect 17592 23802 17644 23808
rect 17408 23112 17460 23118
rect 17604 23089 17632 23802
rect 17408 23054 17460 23060
rect 17590 23080 17646 23089
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17236 22574 17264 22918
rect 17420 22778 17448 23054
rect 17590 23015 17646 23024
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 17144 22358 17264 22386
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16948 18148 17000 18154
rect 16948 18090 17000 18096
rect 17052 17542 17080 18226
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16946 16688 17002 16697
rect 16946 16623 16948 16632
rect 17000 16623 17002 16632
rect 16948 16594 17000 16600
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16684 15162 16712 15982
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16672 14000 16724 14006
rect 16672 13942 16724 13948
rect 16684 12918 16712 13942
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16684 12170 16712 12854
rect 16672 12164 16724 12170
rect 16672 12106 16724 12112
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16580 10124 16632 10130
rect 16580 10066 16632 10072
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 15568 9172 15620 9178
rect 15568 9114 15620 9120
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14936 8430 14964 8910
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14936 7410 14964 8366
rect 15028 8090 15056 8570
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14648 7200 14700 7206
rect 15028 7154 15056 8026
rect 15120 7886 15148 8366
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15304 7206 15332 7822
rect 14648 7142 14700 7148
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 13084 6316 13136 6322
rect 13084 6258 13136 6264
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12728 800 12756 4558
rect 13372 4486 13400 5646
rect 14476 5234 14504 6258
rect 14660 6118 14688 7142
rect 14844 7126 15056 7154
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14844 5710 14872 7126
rect 14924 6928 14976 6934
rect 14924 6870 14976 6876
rect 14936 6254 14964 6870
rect 15488 6866 15516 8842
rect 15580 8634 15608 9114
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 16592 8430 16620 9930
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 8838 16896 9318
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16776 8566 16804 8774
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 7750 15608 8230
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 16776 7410 16804 8502
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15856 6798 15884 7142
rect 15844 6792 15896 6798
rect 15844 6734 15896 6740
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14936 5846 14964 6190
rect 14924 5840 14976 5846
rect 14922 5808 14924 5817
rect 14976 5808 14978 5817
rect 14922 5743 14978 5752
rect 15120 5710 15148 6598
rect 15198 6488 15254 6497
rect 15198 6423 15200 6432
rect 15252 6423 15254 6432
rect 15200 6394 15252 6400
rect 15200 6316 15252 6322
rect 15304 6304 15332 6666
rect 15566 6488 15622 6497
rect 15566 6423 15568 6432
rect 15620 6423 15622 6432
rect 15568 6394 15620 6400
rect 15252 6276 15332 6304
rect 15200 6258 15252 6264
rect 15304 5710 15332 6276
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15672 6118 15700 6258
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5710 15792 6054
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14568 5302 14596 5510
rect 14844 5370 14872 5646
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 15304 5234 15332 5646
rect 16684 5370 16712 6666
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 16960 5166 16988 11154
rect 17144 10674 17172 22170
rect 17236 19174 17264 22358
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17328 20602 17356 20742
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17420 18766 17448 19654
rect 17592 19440 17644 19446
rect 17512 19400 17592 19428
rect 17512 18970 17540 19400
rect 17592 19382 17644 19388
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 17590 18728 17646 18737
rect 17590 18663 17592 18672
rect 17644 18663 17646 18672
rect 17592 18634 17644 18640
rect 17224 18420 17276 18426
rect 17224 18362 17276 18368
rect 17236 16250 17264 18362
rect 17696 18086 17724 32166
rect 18328 31680 18380 31686
rect 18328 31622 18380 31628
rect 18340 31414 18368 31622
rect 18328 31408 18380 31414
rect 18328 31350 18380 31356
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17776 30796 17828 30802
rect 17776 30738 17828 30744
rect 17788 29170 17816 30738
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17880 28762 17908 29106
rect 17868 28756 17920 28762
rect 17868 28698 17920 28704
rect 17972 28150 18000 31282
rect 18420 29504 18472 29510
rect 18420 29446 18472 29452
rect 18144 29232 18196 29238
rect 18144 29174 18196 29180
rect 18156 28558 18184 29174
rect 18432 28694 18460 29446
rect 18420 28688 18472 28694
rect 18420 28630 18472 28636
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 17960 28144 18012 28150
rect 17960 28086 18012 28092
rect 18328 27940 18380 27946
rect 18328 27882 18380 27888
rect 18340 25242 18368 27882
rect 18432 27878 18460 28630
rect 18420 27872 18472 27878
rect 18420 27814 18472 27820
rect 18420 26240 18472 26246
rect 18420 26182 18472 26188
rect 18432 25498 18460 26182
rect 18420 25492 18472 25498
rect 18420 25434 18472 25440
rect 18340 25214 18460 25242
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 18340 24993 18368 25094
rect 18326 24984 18382 24993
rect 18326 24919 18382 24928
rect 18328 24268 18380 24274
rect 18328 24210 18380 24216
rect 18340 23526 18368 24210
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17788 21486 17816 23054
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 18032 21548 18084 21554
rect 18084 21496 18092 21536
rect 18032 21490 18092 21496
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17788 21010 17816 21422
rect 17776 21004 17828 21010
rect 17776 20946 17828 20952
rect 17880 20942 17908 21490
rect 17960 21344 18012 21350
rect 17960 21286 18012 21292
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17776 19508 17828 19514
rect 17776 19450 17828 19456
rect 17788 19310 17816 19450
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17788 18290 17816 18906
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17328 16114 17356 16730
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17328 13938 17356 14554
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17328 12646 17356 13874
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17236 11354 17264 11766
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17236 9042 17264 11290
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17132 7948 17184 7954
rect 17132 7890 17184 7896
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 17052 6662 17080 7346
rect 17144 6798 17172 7890
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17052 5914 17080 6190
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16960 4758 16988 5102
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 13004 800 13032 3470
rect 13280 800 13308 3878
rect 13464 3058 13492 4422
rect 14002 4312 14058 4321
rect 14002 4247 14058 4256
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13556 800 13584 3538
rect 13832 800 13860 3878
rect 14016 3670 14044 4247
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 2650 13952 3538
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14108 800 14136 4558
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 2310 14228 3470
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 3194 14320 3334
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 800 14228 2246
rect 14384 800 14412 3878
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14476 800 14504 2994
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 14660 800 14688 2790
rect 14752 800 14780 4082
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14844 3466 14872 3878
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 14936 800 14964 2858
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 15028 800 15056 2314
rect 15212 800 15240 3470
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15396 800 15424 2790
rect 15672 800 15700 2790
rect 15948 800 15976 3470
rect 16488 2848 16540 2854
rect 16488 2790 16540 2796
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16224 800 16252 2518
rect 16500 800 16528 2790
rect 16776 800 16804 3470
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17052 800 17080 2450
rect 17236 2038 17264 7686
rect 17420 7342 17448 18022
rect 17972 17678 18000 21286
rect 18064 21146 18092 21490
rect 18156 21146 18184 21966
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18248 21554 18276 21626
rect 18236 21548 18288 21554
rect 18236 21490 18288 21496
rect 18236 21412 18288 21418
rect 18236 21354 18288 21360
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18156 20466 18184 21082
rect 18248 20942 18276 21354
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18156 19394 18184 20402
rect 18236 20052 18288 20058
rect 18236 19994 18288 20000
rect 18064 19378 18184 19394
rect 18248 19378 18276 19994
rect 18052 19372 18184 19378
rect 18104 19366 18184 19372
rect 18236 19372 18288 19378
rect 18052 19314 18104 19320
rect 18236 19314 18288 19320
rect 18236 18624 18288 18630
rect 18234 18592 18236 18601
rect 18288 18592 18290 18601
rect 18234 18527 18290 18536
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 17500 17672 17552 17678
rect 17500 17614 17552 17620
rect 17960 17672 18012 17678
rect 18064 17649 18092 17682
rect 18236 17672 18288 17678
rect 17960 17614 18012 17620
rect 18050 17640 18106 17649
rect 17512 16794 17540 17614
rect 18236 17614 18288 17620
rect 18050 17575 18106 17584
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17512 16590 17540 16730
rect 17500 16584 17552 16590
rect 17500 16526 17552 16532
rect 17788 16114 17816 17478
rect 18248 16998 18276 17614
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18234 16688 18290 16697
rect 18234 16623 18290 16632
rect 18248 16590 18276 16623
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17788 15026 17816 16050
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17880 15026 17908 15438
rect 18064 15026 18092 15846
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 15162 18184 15302
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17880 13530 17908 14962
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17880 12918 17908 13466
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12442 17540 12786
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17604 12238 17632 12378
rect 17696 12306 17724 12582
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17696 11898 17724 12242
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17512 11354 17540 11698
rect 17500 11348 17552 11354
rect 17500 11290 17552 11296
rect 17696 11218 17724 11834
rect 17880 11830 17908 12854
rect 17972 12238 18000 13806
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18064 12306 18092 12786
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17972 11150 18000 12038
rect 18340 11558 18368 21830
rect 18432 18086 18460 25214
rect 18524 22234 18552 38150
rect 18616 37262 18644 38218
rect 18800 38010 18828 40054
rect 18984 40050 19012 41482
rect 19352 41206 19380 41482
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19444 41206 19472 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19340 41200 19392 41206
rect 19340 41142 19392 41148
rect 19432 41200 19484 41206
rect 19432 41142 19484 41148
rect 19352 41018 19380 41142
rect 19352 40990 19472 41018
rect 19340 40928 19392 40934
rect 19340 40870 19392 40876
rect 19352 40526 19380 40870
rect 19340 40520 19392 40526
rect 19340 40462 19392 40468
rect 19352 40050 19380 40462
rect 19444 40066 19472 40990
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 18972 40044 19024 40050
rect 18972 39986 19024 39992
rect 19156 40044 19208 40050
rect 19156 39986 19208 39992
rect 19340 40044 19392 40050
rect 19444 40038 19564 40066
rect 19340 39986 19392 39992
rect 19168 38962 19196 39986
rect 19432 39908 19484 39914
rect 19432 39850 19484 39856
rect 19340 39364 19392 39370
rect 19340 39306 19392 39312
rect 19248 39296 19300 39302
rect 19248 39238 19300 39244
rect 19156 38956 19208 38962
rect 19156 38898 19208 38904
rect 18972 38276 19024 38282
rect 18972 38218 19024 38224
rect 18788 38004 18840 38010
rect 18788 37946 18840 37952
rect 18984 37874 19012 38218
rect 18972 37868 19024 37874
rect 18972 37810 19024 37816
rect 18788 37664 18840 37670
rect 18788 37606 18840 37612
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18604 37120 18656 37126
rect 18604 37062 18656 37068
rect 18616 26246 18644 37062
rect 18708 36582 18736 37198
rect 18696 36576 18748 36582
rect 18696 36518 18748 36524
rect 18708 36174 18736 36518
rect 18696 36168 18748 36174
rect 18696 36110 18748 36116
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18708 26382 18736 26862
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18604 26240 18656 26246
rect 18604 26182 18656 26188
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18616 21593 18644 21966
rect 18602 21584 18658 21593
rect 18602 21519 18658 21528
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18524 20534 18552 21286
rect 18616 20641 18644 21422
rect 18602 20632 18658 20641
rect 18602 20567 18658 20576
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18524 17678 18552 19314
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18616 18086 18644 18294
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18524 17542 18552 17614
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18432 12374 18460 17206
rect 18708 16794 18736 26318
rect 18800 22234 18828 37606
rect 19168 37262 19196 38898
rect 19260 38434 19288 39238
rect 19352 39098 19380 39306
rect 19340 39092 19392 39098
rect 19340 39034 19392 39040
rect 19340 38956 19392 38962
rect 19340 38898 19392 38904
rect 19352 38554 19380 38898
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 19260 38406 19380 38434
rect 19352 38214 19380 38406
rect 19340 38208 19392 38214
rect 19340 38150 19392 38156
rect 19352 37874 19380 38150
rect 19340 37868 19392 37874
rect 19340 37810 19392 37816
rect 19156 37256 19208 37262
rect 19156 37198 19208 37204
rect 19168 34610 19196 37198
rect 19352 35834 19380 37810
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19340 35556 19392 35562
rect 19340 35498 19392 35504
rect 19352 35086 19380 35498
rect 19444 35086 19472 39850
rect 19536 39506 19564 40038
rect 19996 39574 20024 41568
rect 20168 40044 20220 40050
rect 20168 39986 20220 39992
rect 20180 39642 20208 39986
rect 20260 39840 20312 39846
rect 20260 39782 20312 39788
rect 20168 39636 20220 39642
rect 20168 39578 20220 39584
rect 19984 39568 20036 39574
rect 19984 39510 20036 39516
rect 19524 39500 19576 39506
rect 19524 39442 19576 39448
rect 19984 39364 20036 39370
rect 19984 39306 20036 39312
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19800 37868 19852 37874
rect 19800 37810 19852 37816
rect 19812 37466 19840 37810
rect 19996 37738 20024 39306
rect 19984 37732 20036 37738
rect 19984 37674 20036 37680
rect 19800 37460 19852 37466
rect 19800 37402 19852 37408
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19524 35828 19576 35834
rect 19524 35770 19576 35776
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19432 35080 19484 35086
rect 19432 35022 19484 35028
rect 19536 34950 19564 35770
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 19524 34944 19576 34950
rect 19524 34886 19576 34892
rect 19156 34604 19208 34610
rect 19156 34546 19208 34552
rect 19064 33516 19116 33522
rect 19064 33458 19116 33464
rect 19076 31346 19104 33458
rect 19168 33114 19196 34546
rect 19352 34490 19380 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19996 34626 20024 37674
rect 20076 35080 20128 35086
rect 20076 35022 20128 35028
rect 20088 34746 20116 35022
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19432 34604 19484 34610
rect 19996 34598 20116 34626
rect 19432 34546 19484 34552
rect 19260 34462 19380 34490
rect 19260 33862 19288 34462
rect 19340 34400 19392 34406
rect 19340 34342 19392 34348
rect 19248 33856 19300 33862
rect 19248 33798 19300 33804
rect 19352 33658 19380 34342
rect 19444 33930 19472 34546
rect 19432 33924 19484 33930
rect 19432 33866 19484 33872
rect 19984 33924 20036 33930
rect 19984 33866 20036 33872
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19996 33658 20024 33866
rect 19340 33652 19392 33658
rect 19340 33594 19392 33600
rect 19984 33652 20036 33658
rect 19984 33594 20036 33600
rect 20088 33454 20116 34598
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 20076 33448 20128 33454
rect 20076 33390 20128 33396
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19064 31340 19116 31346
rect 19064 31282 19116 31288
rect 19340 31136 19392 31142
rect 19340 31078 19392 31084
rect 19352 29578 19380 31078
rect 19444 30258 19472 31758
rect 20180 31754 20208 33934
rect 20272 33522 20300 39782
rect 20364 39642 20392 41754
rect 20352 39636 20404 39642
rect 20352 39578 20404 39584
rect 20364 39438 20392 39578
rect 20352 39432 20404 39438
rect 20352 39374 20404 39380
rect 20364 38894 20392 39374
rect 20352 38888 20404 38894
rect 20352 38830 20404 38836
rect 20456 38010 20484 42638
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 24768 42016 24820 42022
rect 24768 41958 24820 41964
rect 23940 41132 23992 41138
rect 23940 41074 23992 41080
rect 23112 40928 23164 40934
rect 23112 40870 23164 40876
rect 22652 40384 22704 40390
rect 22652 40326 22704 40332
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22560 40044 22612 40050
rect 22560 39986 22612 39992
rect 21272 39840 21324 39846
rect 21272 39782 21324 39788
rect 21284 38962 21312 39782
rect 22296 39438 22324 39986
rect 22572 39642 22600 39986
rect 22560 39636 22612 39642
rect 22560 39578 22612 39584
rect 22100 39432 22152 39438
rect 22100 39374 22152 39380
rect 22284 39432 22336 39438
rect 22284 39374 22336 39380
rect 21916 39024 21968 39030
rect 21916 38966 21968 38972
rect 21272 38956 21324 38962
rect 21272 38898 21324 38904
rect 21928 38758 21956 38966
rect 21916 38752 21968 38758
rect 21916 38694 21968 38700
rect 20444 38004 20496 38010
rect 20444 37946 20496 37952
rect 21180 37732 21232 37738
rect 21180 37674 21232 37680
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 20732 36718 20760 37198
rect 21192 37194 21220 37674
rect 21180 37188 21232 37194
rect 21180 37130 21232 37136
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 20732 34950 20760 36654
rect 20812 36576 20864 36582
rect 20812 36518 20864 36524
rect 20824 36378 20852 36518
rect 20812 36372 20864 36378
rect 20812 36314 20864 36320
rect 20824 36174 20852 36314
rect 20812 36168 20864 36174
rect 21824 36168 21876 36174
rect 20864 36128 20944 36156
rect 20812 36110 20864 36116
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20732 34678 20760 34886
rect 20720 34672 20772 34678
rect 20720 34614 20772 34620
rect 20732 34066 20760 34614
rect 20720 34060 20772 34066
rect 20772 34020 20852 34048
rect 20720 34002 20772 34008
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20352 33108 20404 33114
rect 20352 33050 20404 33056
rect 20088 31726 20208 31754
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19984 30660 20036 30666
rect 19984 30602 20036 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 19892 30252 19944 30258
rect 19892 30194 19944 30200
rect 19432 30048 19484 30054
rect 19432 29990 19484 29996
rect 19444 29646 19472 29990
rect 19432 29640 19484 29646
rect 19432 29582 19484 29588
rect 19340 29572 19392 29578
rect 19904 29560 19932 30194
rect 19996 29850 20024 30602
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19904 29532 20024 29560
rect 19340 29514 19392 29520
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19996 29170 20024 29532
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19628 28626 19656 28902
rect 19616 28620 19668 28626
rect 19616 28562 19668 28568
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19352 27606 19380 28018
rect 19996 27878 20024 29106
rect 19984 27872 20036 27878
rect 19984 27814 20036 27820
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 18972 26988 19024 26994
rect 18972 26930 19024 26936
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18892 23662 18920 24754
rect 18984 24274 19012 26930
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 19076 25922 19104 26386
rect 19168 26042 19196 26930
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19720 26382 19748 26726
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19156 26036 19208 26042
rect 19156 25978 19208 25984
rect 19260 25974 19288 26182
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19248 25968 19300 25974
rect 19076 25894 19196 25922
rect 19248 25910 19300 25916
rect 19168 24682 19196 25894
rect 19248 25696 19300 25702
rect 19248 25638 19300 25644
rect 19260 25362 19288 25638
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19444 24954 19472 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19432 24948 19484 24954
rect 19432 24890 19484 24896
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19156 24676 19208 24682
rect 19156 24618 19208 24624
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18880 23656 18932 23662
rect 18880 23598 18932 23604
rect 18892 22438 18920 23598
rect 18880 22432 18932 22438
rect 18880 22374 18932 22380
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18800 17270 18828 21830
rect 18984 21554 19012 23666
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18984 21078 19012 21490
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18892 18834 18920 19110
rect 18880 18828 18932 18834
rect 18880 18770 18932 18776
rect 19076 18578 19104 23734
rect 19168 23594 19196 24618
rect 19352 24342 19380 24754
rect 19996 24410 20024 27814
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19340 24336 19392 24342
rect 19340 24278 19392 24284
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19168 23186 19196 23530
rect 19156 23180 19208 23186
rect 19156 23122 19208 23128
rect 19248 22432 19300 22438
rect 19248 22374 19300 22380
rect 19260 22273 19288 22374
rect 19246 22264 19302 22273
rect 19246 22199 19302 22208
rect 19444 21962 19472 24006
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23050 20024 24142
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20088 22438 20116 31726
rect 20364 26518 20392 33050
rect 20824 32910 20852 34020
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20916 32722 20944 36128
rect 21824 36110 21876 36116
rect 21836 35834 21864 36110
rect 21824 35828 21876 35834
rect 21824 35770 21876 35776
rect 21928 35698 21956 38694
rect 22112 38282 22140 39374
rect 22296 38962 22324 39374
rect 22284 38956 22336 38962
rect 22284 38898 22336 38904
rect 22560 38956 22612 38962
rect 22560 38898 22612 38904
rect 22192 38888 22244 38894
rect 22192 38830 22244 38836
rect 22100 38276 22152 38282
rect 22100 38218 22152 38224
rect 22204 36106 22232 38830
rect 22296 36174 22324 38898
rect 22572 38554 22600 38898
rect 22560 38548 22612 38554
rect 22560 38490 22612 38496
rect 22664 38350 22692 40326
rect 23124 40118 23152 40870
rect 23480 40452 23532 40458
rect 23480 40394 23532 40400
rect 23756 40452 23808 40458
rect 23756 40394 23808 40400
rect 23112 40112 23164 40118
rect 23112 40054 23164 40060
rect 23204 40044 23256 40050
rect 23204 39986 23256 39992
rect 22836 39976 22888 39982
rect 22836 39918 22888 39924
rect 22848 39438 22876 39918
rect 23216 39642 23244 39986
rect 23204 39636 23256 39642
rect 23204 39578 23256 39584
rect 22836 39432 22888 39438
rect 22836 39374 22888 39380
rect 23112 39432 23164 39438
rect 23112 39374 23164 39380
rect 22848 38894 22876 39374
rect 22928 38956 22980 38962
rect 22928 38898 22980 38904
rect 22836 38888 22888 38894
rect 22836 38830 22888 38836
rect 22652 38344 22704 38350
rect 22652 38286 22704 38292
rect 22468 36576 22520 36582
rect 22468 36518 22520 36524
rect 22560 36576 22612 36582
rect 22560 36518 22612 36524
rect 22284 36168 22336 36174
rect 22284 36110 22336 36116
rect 22192 36100 22244 36106
rect 22192 36042 22244 36048
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 21916 35692 21968 35698
rect 21916 35634 21968 35640
rect 21824 32836 21876 32842
rect 21824 32778 21876 32784
rect 20824 32694 20944 32722
rect 21088 32768 21140 32774
rect 21088 32710 21140 32716
rect 20628 30592 20680 30598
rect 20628 30534 20680 30540
rect 20640 30326 20668 30534
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20640 29714 20668 30262
rect 20628 29708 20680 29714
rect 20628 29650 20680 29656
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20628 29232 20680 29238
rect 20732 29186 20760 29446
rect 20680 29180 20760 29186
rect 20628 29174 20760 29180
rect 20640 29158 20760 29174
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20444 28008 20496 28014
rect 20444 27950 20496 27956
rect 20352 26512 20404 26518
rect 20352 26454 20404 26460
rect 20364 26314 20392 26454
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20260 24812 20312 24818
rect 20260 24754 20312 24760
rect 20272 24274 20300 24754
rect 20260 24268 20312 24274
rect 20260 24210 20312 24216
rect 20272 23866 20300 24210
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19432 21956 19484 21962
rect 19432 21898 19484 21904
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21486 20024 21830
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19340 20800 19392 20806
rect 19340 20742 19392 20748
rect 19352 20602 19380 20742
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19168 18630 19196 19110
rect 19352 18834 19380 20538
rect 20076 19780 20128 19786
rect 20076 19722 20128 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19984 18896 20036 18902
rect 19984 18838 20036 18844
rect 19248 18828 19300 18834
rect 19248 18770 19300 18776
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 18892 18550 19104 18578
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 18788 17264 18840 17270
rect 18788 17206 18840 17212
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18708 12102 18736 12174
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18432 11370 18460 11494
rect 18340 11342 18460 11370
rect 18708 11354 18736 12038
rect 18696 11348 18748 11354
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 18144 9648 18196 9654
rect 18144 9590 18196 9596
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17408 7336 17460 7342
rect 17408 7278 17460 7284
rect 17868 6656 17920 6662
rect 17868 6598 17920 6604
rect 17880 6390 17908 6598
rect 17868 6384 17920 6390
rect 17868 6326 17920 6332
rect 17880 5642 17908 6326
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17880 4486 17908 5102
rect 17972 5030 18000 9454
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 18064 8634 18092 8842
rect 18156 8634 18184 9590
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 18156 8090 18184 8570
rect 18340 8498 18368 11342
rect 18696 11290 18748 11296
rect 18708 11150 18736 11290
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10470 18552 11018
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18524 9382 18552 10406
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 8906 18552 9318
rect 18616 9178 18644 10542
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18512 8900 18564 8906
rect 18512 8842 18564 8848
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18340 7818 18368 8434
rect 18524 8090 18552 8434
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18616 7886 18644 9114
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18708 8498 18736 8570
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18604 7880 18656 7886
rect 18604 7822 18656 7828
rect 18328 7812 18380 7818
rect 18328 7754 18380 7760
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 18064 6730 18092 7210
rect 18052 6724 18104 6730
rect 18052 6666 18104 6672
rect 18708 6662 18736 8434
rect 18800 8362 18828 16934
rect 18892 11762 18920 18550
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18892 9926 18920 10610
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18800 7818 18828 8298
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18984 6186 19012 18362
rect 19260 18290 19288 18770
rect 19996 18766 20024 18838
rect 19984 18760 20036 18766
rect 19890 18728 19946 18737
rect 19340 18692 19392 18698
rect 19984 18702 20036 18708
rect 19890 18663 19892 18672
rect 19340 18634 19392 18640
rect 19944 18663 19946 18672
rect 19892 18634 19944 18640
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 17066 19288 18226
rect 19352 18204 19380 18634
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19444 18358 19472 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18352 19484 18358
rect 19708 18352 19760 18358
rect 19432 18294 19484 18300
rect 19706 18320 19708 18329
rect 19760 18320 19762 18329
rect 19996 18290 20024 18702
rect 19706 18255 19762 18264
rect 19984 18284 20036 18290
rect 19720 18204 19748 18255
rect 19984 18226 20036 18232
rect 19352 18176 19748 18204
rect 19996 17746 20024 18226
rect 20088 17882 20116 19722
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19984 17740 20036 17746
rect 19984 17682 20036 17688
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19248 17060 19300 17066
rect 19168 17020 19248 17048
rect 19168 10198 19196 17020
rect 19248 17002 19300 17008
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19444 16114 19472 16730
rect 19536 16590 19564 16934
rect 19720 16794 19748 17070
rect 19996 17066 20024 17274
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19536 16454 19564 16526
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19260 15570 19288 16050
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19352 14890 19380 15982
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19996 14618 20024 17002
rect 20088 16794 20116 17614
rect 20180 17338 20208 23734
rect 20260 23180 20312 23186
rect 20260 23122 20312 23128
rect 20272 23050 20300 23122
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20364 22438 20392 26250
rect 20456 23798 20484 27950
rect 20548 24154 20576 28902
rect 20732 28082 20760 29158
rect 20824 28694 20852 32694
rect 21100 32502 21128 32710
rect 21836 32502 21864 32778
rect 21088 32496 21140 32502
rect 21088 32438 21140 32444
rect 21640 32496 21692 32502
rect 21640 32438 21692 32444
rect 21824 32496 21876 32502
rect 21824 32438 21876 32444
rect 20904 32428 20956 32434
rect 20904 32370 20956 32376
rect 20916 32026 20944 32370
rect 20904 32020 20956 32026
rect 20904 31962 20956 31968
rect 21652 30734 21680 32438
rect 21928 31482 21956 35634
rect 22112 34950 22140 35702
rect 22100 34944 22152 34950
rect 22100 34886 22152 34892
rect 22008 33108 22060 33114
rect 22008 33050 22060 33056
rect 22020 32434 22048 33050
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 21916 31476 21968 31482
rect 21916 31418 21968 31424
rect 20904 30728 20956 30734
rect 20904 30670 20956 30676
rect 21640 30728 21692 30734
rect 21640 30670 21692 30676
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 20916 30190 20944 30670
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 20904 30184 20956 30190
rect 20904 30126 20956 30132
rect 20916 29646 20944 30126
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 20916 29170 20944 29582
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20812 28688 20864 28694
rect 20812 28630 20864 28636
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20824 26382 20852 27406
rect 20916 26994 20944 29106
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20720 26036 20772 26042
rect 20720 25978 20772 25984
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 24886 20668 25094
rect 20628 24880 20680 24886
rect 20628 24822 20680 24828
rect 20640 24274 20668 24822
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20548 24126 20668 24154
rect 20444 23792 20496 23798
rect 20444 23734 20496 23740
rect 20444 23044 20496 23050
rect 20444 22986 20496 22992
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20456 22642 20484 22986
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20272 18465 20300 18634
rect 20258 18456 20314 18465
rect 20364 18426 20392 19314
rect 20456 18902 20484 22578
rect 20548 22574 20576 22986
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20536 22092 20588 22098
rect 20536 22034 20588 22040
rect 20548 21865 20576 22034
rect 20534 21856 20590 21865
rect 20534 21791 20590 21800
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20548 20806 20576 21490
rect 20536 20800 20588 20806
rect 20536 20742 20588 20748
rect 20444 18896 20496 18902
rect 20444 18838 20496 18844
rect 20442 18728 20498 18737
rect 20442 18663 20498 18672
rect 20258 18391 20314 18400
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20088 16590 20116 16730
rect 20166 16688 20222 16697
rect 20166 16623 20222 16632
rect 20180 16590 20208 16623
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20076 15360 20128 15366
rect 20180 15348 20208 16526
rect 20272 15910 20300 18226
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20364 15722 20392 18362
rect 20272 15694 20392 15722
rect 20272 15502 20300 15694
rect 20456 15502 20484 18663
rect 20548 18426 20576 20742
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20640 18290 20668 24126
rect 20732 22642 20760 25978
rect 20824 25974 20852 26318
rect 20812 25968 20864 25974
rect 20812 25910 20864 25916
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20824 21486 20852 25910
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 20916 21894 20944 22986
rect 21008 22642 21036 30534
rect 21836 29782 21864 30670
rect 21180 29776 21232 29782
rect 21180 29718 21232 29724
rect 21824 29776 21876 29782
rect 21824 29718 21876 29724
rect 21088 29572 21140 29578
rect 21088 29514 21140 29520
rect 21100 29238 21128 29514
rect 21088 29232 21140 29238
rect 21088 29174 21140 29180
rect 21088 28688 21140 28694
rect 21088 28630 21140 28636
rect 21100 26042 21128 28630
rect 21088 26036 21140 26042
rect 21088 25978 21140 25984
rect 21100 25945 21128 25978
rect 21086 25936 21142 25945
rect 21086 25871 21142 25880
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21192 22094 21220 29718
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21272 27532 21324 27538
rect 21272 27474 21324 27480
rect 21284 26450 21312 27474
rect 21468 26858 21496 29582
rect 21560 27526 21772 27554
rect 21560 27334 21588 27526
rect 21640 27464 21692 27470
rect 21640 27406 21692 27412
rect 21744 27418 21772 27526
rect 21836 27418 21864 29718
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21652 26926 21680 27406
rect 21744 27390 21864 27418
rect 21640 26920 21692 26926
rect 21640 26862 21692 26868
rect 21456 26852 21508 26858
rect 21456 26794 21508 26800
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21284 26042 21312 26386
rect 21652 26314 21680 26862
rect 21640 26308 21692 26314
rect 21640 26250 21692 26256
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21652 25838 21680 26250
rect 21640 25832 21692 25838
rect 21640 25774 21692 25780
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21468 23730 21496 24346
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21560 23730 21588 23802
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21548 23724 21600 23730
rect 21548 23666 21600 23672
rect 21272 23248 21324 23254
rect 21272 23190 21324 23196
rect 21284 22166 21312 23190
rect 21652 22642 21680 25774
rect 21744 23866 21772 27390
rect 21824 27328 21876 27334
rect 21824 27270 21876 27276
rect 21836 27062 21864 27270
rect 21824 27056 21876 27062
rect 21824 26998 21876 27004
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 21732 23860 21784 23866
rect 21732 23802 21784 23808
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 21272 22160 21324 22166
rect 21272 22102 21324 22108
rect 21008 22066 21220 22094
rect 21836 22094 21864 26522
rect 21928 24410 21956 31418
rect 22008 30660 22060 30666
rect 22008 30602 22060 30608
rect 22020 30326 22048 30602
rect 22008 30320 22060 30326
rect 22008 30262 22060 30268
rect 22020 29578 22048 30262
rect 22112 30258 22140 34886
rect 22204 32434 22232 36042
rect 22296 34898 22324 36110
rect 22480 36106 22508 36518
rect 22468 36100 22520 36106
rect 22468 36042 22520 36048
rect 22376 36032 22428 36038
rect 22376 35974 22428 35980
rect 22388 35018 22416 35974
rect 22376 35012 22428 35018
rect 22376 34954 22428 34960
rect 22296 34870 22508 34898
rect 22376 34060 22428 34066
rect 22376 34002 22428 34008
rect 22388 33862 22416 34002
rect 22376 33856 22428 33862
rect 22376 33798 22428 33804
rect 22192 32428 22244 32434
rect 22192 32370 22244 32376
rect 22204 31414 22232 32370
rect 22192 31408 22244 31414
rect 22192 31350 22244 31356
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 22008 29572 22060 29578
rect 22008 29514 22060 29520
rect 22388 29458 22416 33798
rect 22480 32434 22508 34870
rect 22468 32428 22520 32434
rect 22468 32370 22520 32376
rect 22480 30716 22508 32370
rect 22572 30818 22600 36518
rect 22664 36174 22692 38286
rect 22836 38276 22888 38282
rect 22940 38264 22968 38898
rect 22888 38236 22968 38264
rect 22836 38218 22888 38224
rect 22744 37120 22796 37126
rect 22744 37062 22796 37068
rect 22756 36786 22784 37062
rect 22744 36780 22796 36786
rect 22744 36722 22796 36728
rect 22652 36168 22704 36174
rect 22652 36110 22704 36116
rect 22652 36032 22704 36038
rect 22652 35974 22704 35980
rect 22664 34066 22692 35974
rect 22848 35698 22876 38218
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22756 31754 22784 33798
rect 22848 31890 22876 35634
rect 23020 34400 23072 34406
rect 23020 34342 23072 34348
rect 23032 33930 23060 34342
rect 23020 33924 23072 33930
rect 23020 33866 23072 33872
rect 23032 33590 23060 33866
rect 23020 33584 23072 33590
rect 23020 33526 23072 33532
rect 22928 33516 22980 33522
rect 22928 33458 22980 33464
rect 22940 32434 22968 33458
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 22940 32026 22968 32370
rect 23124 32298 23152 39374
rect 23492 39098 23520 40394
rect 23768 39982 23796 40394
rect 23756 39976 23808 39982
rect 23756 39918 23808 39924
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23480 39092 23532 39098
rect 23480 39034 23532 39040
rect 23676 38962 23704 39782
rect 23848 39364 23900 39370
rect 23848 39306 23900 39312
rect 23860 39098 23888 39306
rect 23848 39092 23900 39098
rect 23848 39034 23900 39040
rect 23664 38956 23716 38962
rect 23664 38898 23716 38904
rect 23572 38820 23624 38826
rect 23572 38762 23624 38768
rect 23584 38554 23612 38762
rect 23572 38548 23624 38554
rect 23572 38490 23624 38496
rect 23584 37262 23612 38490
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23400 36802 23428 37198
rect 23296 36780 23348 36786
rect 23400 36774 23520 36802
rect 23676 36786 23704 38898
rect 23296 36722 23348 36728
rect 23308 36106 23336 36722
rect 23388 36712 23440 36718
rect 23388 36654 23440 36660
rect 23400 36156 23428 36654
rect 23492 36582 23520 36774
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23480 36576 23532 36582
rect 23480 36518 23532 36524
rect 23480 36168 23532 36174
rect 23400 36128 23480 36156
rect 23296 36100 23348 36106
rect 23296 36042 23348 36048
rect 23400 35494 23428 36128
rect 23480 36110 23532 36116
rect 23664 36032 23716 36038
rect 23662 36000 23664 36009
rect 23716 36000 23718 36009
rect 23662 35935 23718 35944
rect 23664 35556 23716 35562
rect 23664 35498 23716 35504
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 23400 33998 23428 35430
rect 23388 33992 23440 33998
rect 23388 33934 23440 33940
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23112 32292 23164 32298
rect 23112 32234 23164 32240
rect 22928 32020 22980 32026
rect 22928 31962 22980 31968
rect 22836 31884 22888 31890
rect 22836 31826 22888 31832
rect 22756 31726 22876 31754
rect 22572 30790 22784 30818
rect 22560 30728 22612 30734
rect 22480 30688 22560 30716
rect 22560 30670 22612 30676
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22468 29504 22520 29510
rect 22388 29452 22468 29458
rect 22388 29446 22520 29452
rect 22388 29430 22508 29446
rect 22192 28620 22244 28626
rect 22192 28562 22244 28568
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 22020 27538 22048 27814
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22020 26450 22048 27474
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 22204 26194 22232 28562
rect 22204 26166 22324 26194
rect 22190 25936 22246 25945
rect 22190 25871 22192 25880
rect 22244 25871 22246 25880
rect 22192 25842 22244 25848
rect 22192 25696 22244 25702
rect 22192 25638 22244 25644
rect 21916 24404 21968 24410
rect 21916 24346 21968 24352
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22112 22710 22140 23530
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 22008 22094 22060 22098
rect 21836 22092 22060 22094
rect 21836 22066 22008 22092
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20824 17270 20852 18158
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 15978 20576 17138
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20640 16250 20668 16458
rect 20812 16448 20864 16454
rect 20812 16390 20864 16396
rect 20824 16250 20852 16390
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20536 15972 20588 15978
rect 20536 15914 20588 15920
rect 20548 15502 20576 15914
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20444 15496 20496 15502
rect 20444 15438 20496 15444
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20128 15320 20208 15348
rect 20076 15302 20128 15308
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19260 13530 19288 13942
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19352 9926 19380 14554
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20088 12730 20116 15302
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 12850 20208 13670
rect 20272 13326 20300 15438
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20364 14414 20392 15302
rect 20456 14822 20484 15438
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20548 14822 20576 14962
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20352 14408 20404 14414
rect 20536 14408 20588 14414
rect 20352 14350 20404 14356
rect 20456 14368 20536 14396
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20456 12850 20484 14368
rect 20640 14396 20668 16186
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20588 14368 20668 14396
rect 20536 14350 20588 14356
rect 20732 13326 20760 15846
rect 20812 15088 20864 15094
rect 20812 15030 20864 15036
rect 20824 14618 20852 15030
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 12850 20576 13126
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20444 12844 20496 12850
rect 20444 12786 20496 12792
rect 20536 12844 20588 12850
rect 20536 12786 20588 12792
rect 19996 12702 20116 12730
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19444 9994 19472 12106
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19432 9988 19484 9994
rect 19432 9930 19484 9936
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19260 8974 19288 9862
rect 19352 9586 19380 9862
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19444 9450 19472 9930
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9586 20024 12702
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 12238 20116 12582
rect 20076 12232 20128 12238
rect 20076 12174 20128 12180
rect 20180 11898 20208 12786
rect 20732 12442 20760 13262
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20548 12170 20576 12378
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20456 11830 20484 12038
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20916 11665 20944 21830
rect 21008 18766 21036 22066
rect 22008 22034 22060 22040
rect 22020 21622 22048 22034
rect 22204 22030 22232 25638
rect 22296 24138 22324 26166
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22388 23338 22416 25434
rect 22480 23526 22508 29430
rect 22560 27396 22612 27402
rect 22560 27338 22612 27344
rect 22572 26042 22600 27338
rect 22560 26036 22612 26042
rect 22560 25978 22612 25984
rect 22664 25362 22692 29990
rect 22652 25356 22704 25362
rect 22652 25298 22704 25304
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22664 24206 22692 24754
rect 22756 24342 22784 30790
rect 22848 28626 22876 31726
rect 22928 31748 22980 31754
rect 22928 31690 22980 31696
rect 22940 31346 22968 31690
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 23124 28558 23152 30194
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23020 27872 23072 27878
rect 23020 27814 23072 27820
rect 23032 27690 23060 27814
rect 23032 27674 23152 27690
rect 23032 27668 23164 27674
rect 23032 27662 23112 27668
rect 22928 26784 22980 26790
rect 22848 26732 22928 26738
rect 22848 26726 22980 26732
rect 22848 26710 22968 26726
rect 22744 24336 22796 24342
rect 22744 24278 22796 24284
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22468 23520 22520 23526
rect 22468 23462 22520 23468
rect 22388 23310 22508 23338
rect 22376 22976 22428 22982
rect 22376 22918 22428 22924
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 21272 21616 21324 21622
rect 21272 21558 21324 21564
rect 22008 21616 22060 21622
rect 22008 21558 22060 21564
rect 21284 20942 21312 21558
rect 21732 21480 21784 21486
rect 21732 21422 21784 21428
rect 21744 21010 21772 21422
rect 22284 21072 22336 21078
rect 22284 21014 22336 21020
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21100 20534 21128 20878
rect 21284 20602 21312 20878
rect 21272 20596 21324 20602
rect 21272 20538 21324 20544
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 21284 20058 21312 20538
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21744 19514 21772 20946
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22112 20262 22140 20878
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22204 20534 22232 20742
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 22100 20256 22152 20262
rect 22100 20198 22152 20204
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 21008 18290 21036 18566
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 21008 17202 21036 18226
rect 21732 18216 21784 18222
rect 21732 18158 21784 18164
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21192 17882 21220 18022
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21008 16454 21036 17138
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21100 15162 21128 17614
rect 21744 17202 21772 18158
rect 22112 17542 22140 20198
rect 22296 20058 22324 21014
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22100 17536 22152 17542
rect 22100 17478 22152 17484
rect 21732 17196 21784 17202
rect 21732 17138 21784 17144
rect 21916 17196 21968 17202
rect 21916 17138 21968 17144
rect 21744 16250 21772 17138
rect 21928 17066 21956 17138
rect 21916 17060 21968 17066
rect 21916 17002 21968 17008
rect 21928 16794 21956 17002
rect 21916 16788 21968 16794
rect 21916 16730 21968 16736
rect 21732 16244 21784 16250
rect 21732 16186 21784 16192
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 22008 15156 22060 15162
rect 22008 15098 22060 15104
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21100 14006 21128 14350
rect 21088 14000 21140 14006
rect 21088 13942 21140 13948
rect 20902 11656 20958 11665
rect 20902 11591 20958 11600
rect 21100 10742 21128 13942
rect 21468 13394 21496 14894
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21744 14385 21772 14486
rect 21730 14376 21786 14385
rect 22020 14346 22048 15098
rect 22112 14958 22140 17478
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 21730 14311 21732 14320
rect 21784 14311 21786 14320
rect 22008 14340 22060 14346
rect 21732 14282 21784 14288
rect 22008 14282 22060 14288
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21744 12986 21772 14282
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 22388 11354 22416 22918
rect 22480 22234 22508 23310
rect 22848 23100 22876 26710
rect 22928 24880 22980 24886
rect 22928 24822 22980 24828
rect 22940 24138 22968 24822
rect 22928 24132 22980 24138
rect 22928 24074 22980 24080
rect 22940 23322 22968 24074
rect 22928 23316 22980 23322
rect 22928 23258 22980 23264
rect 23032 23100 23060 27662
rect 23112 27610 23164 27616
rect 23216 27402 23244 33798
rect 23584 33590 23612 33798
rect 23572 33584 23624 33590
rect 23572 33526 23624 33532
rect 23676 33114 23704 35498
rect 23952 33590 23980 41074
rect 24308 40384 24360 40390
rect 24308 40326 24360 40332
rect 24320 39506 24348 40326
rect 24308 39500 24360 39506
rect 24308 39442 24360 39448
rect 24216 37868 24268 37874
rect 24216 37810 24268 37816
rect 24032 37664 24084 37670
rect 24032 37606 24084 37612
rect 24044 37126 24072 37606
rect 24032 37120 24084 37126
rect 24032 37062 24084 37068
rect 24044 36786 24072 37062
rect 24032 36780 24084 36786
rect 24032 36722 24084 36728
rect 23940 33584 23992 33590
rect 23940 33526 23992 33532
rect 23952 33114 23980 33526
rect 23664 33108 23716 33114
rect 23664 33050 23716 33056
rect 23940 33108 23992 33114
rect 23940 33050 23992 33056
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23584 32366 23612 32710
rect 23572 32360 23624 32366
rect 23572 32302 23624 32308
rect 23676 31754 23704 33050
rect 23848 32360 23900 32366
rect 23848 32302 23900 32308
rect 23584 31726 23704 31754
rect 23388 29096 23440 29102
rect 23388 29038 23440 29044
rect 23400 28762 23428 29038
rect 23388 28756 23440 28762
rect 23388 28698 23440 28704
rect 23584 28082 23612 31726
rect 23860 31482 23888 32302
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 23664 30728 23716 30734
rect 23664 30670 23716 30676
rect 23676 29170 23704 30670
rect 23664 29164 23716 29170
rect 23664 29106 23716 29112
rect 23860 28218 23888 31078
rect 23952 30818 23980 32166
rect 24044 31142 24072 36722
rect 24124 36712 24176 36718
rect 24124 36654 24176 36660
rect 24136 36378 24164 36654
rect 24124 36372 24176 36378
rect 24124 36314 24176 36320
rect 24124 34604 24176 34610
rect 24124 34546 24176 34552
rect 24136 33658 24164 34546
rect 24228 33930 24256 37810
rect 24320 33998 24348 39442
rect 24492 37664 24544 37670
rect 24492 37606 24544 37612
rect 24504 36922 24532 37606
rect 24676 37460 24728 37466
rect 24676 37402 24728 37408
rect 24688 36922 24716 37402
rect 24492 36916 24544 36922
rect 24492 36858 24544 36864
rect 24676 36916 24728 36922
rect 24676 36858 24728 36864
rect 24504 36174 24532 36858
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 24492 36032 24544 36038
rect 24492 35974 24544 35980
rect 24504 35494 24532 35974
rect 24688 35894 24716 36858
rect 24780 36768 24808 41958
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 58164 41608 58216 41614
rect 58162 41576 58164 41585
rect 58216 41576 58218 41585
rect 58162 41511 58218 41520
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 27804 41132 27856 41138
rect 27804 41074 27856 41080
rect 27712 41064 27764 41070
rect 27712 41006 27764 41012
rect 27724 40594 27752 41006
rect 27816 40730 27844 41074
rect 29276 40928 29328 40934
rect 29276 40870 29328 40876
rect 27804 40724 27856 40730
rect 27804 40666 27856 40672
rect 27712 40588 27764 40594
rect 27712 40530 27764 40536
rect 25964 40520 26016 40526
rect 25964 40462 26016 40468
rect 27252 40520 27304 40526
rect 27252 40462 27304 40468
rect 24952 40112 25004 40118
rect 24952 40054 25004 40060
rect 24860 36780 24912 36786
rect 24780 36740 24860 36768
rect 24780 36038 24808 36740
rect 24860 36722 24912 36728
rect 24860 36168 24912 36174
rect 24860 36110 24912 36116
rect 24768 36032 24820 36038
rect 24768 35974 24820 35980
rect 24688 35866 24808 35894
rect 24492 35488 24544 35494
rect 24492 35430 24544 35436
rect 24504 34474 24532 35430
rect 24492 34468 24544 34474
rect 24492 34410 24544 34416
rect 24308 33992 24360 33998
rect 24308 33934 24360 33940
rect 24216 33924 24268 33930
rect 24216 33866 24268 33872
rect 24124 33652 24176 33658
rect 24124 33594 24176 33600
rect 24032 31136 24084 31142
rect 24032 31078 24084 31084
rect 23952 30790 24072 30818
rect 23940 28688 23992 28694
rect 23940 28630 23992 28636
rect 23848 28212 23900 28218
rect 23848 28154 23900 28160
rect 23572 28076 23624 28082
rect 23572 28018 23624 28024
rect 23204 27396 23256 27402
rect 23204 27338 23256 27344
rect 23756 27396 23808 27402
rect 23756 27338 23808 27344
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 23204 26512 23256 26518
rect 23204 26454 23256 26460
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23124 25294 23152 25842
rect 23216 25838 23244 26454
rect 23400 26042 23428 27270
rect 23664 26784 23716 26790
rect 23664 26726 23716 26732
rect 23676 26314 23704 26726
rect 23664 26308 23716 26314
rect 23664 26250 23716 26256
rect 23480 26240 23532 26246
rect 23480 26182 23532 26188
rect 23388 26036 23440 26042
rect 23388 25978 23440 25984
rect 23204 25832 23256 25838
rect 23204 25774 23256 25780
rect 23388 25764 23440 25770
rect 23388 25706 23440 25712
rect 23296 25696 23348 25702
rect 23296 25638 23348 25644
rect 23308 25514 23336 25638
rect 23216 25486 23336 25514
rect 23400 25498 23428 25706
rect 23388 25492 23440 25498
rect 23216 25294 23244 25486
rect 23388 25434 23440 25440
rect 23492 25294 23520 26182
rect 23572 25968 23624 25974
rect 23572 25910 23624 25916
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23204 25288 23256 25294
rect 23204 25230 23256 25236
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23124 24818 23152 25230
rect 23584 25158 23612 25910
rect 23768 25888 23796 27338
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23860 26246 23888 27270
rect 23848 26240 23900 26246
rect 23848 26182 23900 26188
rect 23848 25900 23900 25906
rect 23768 25860 23848 25888
rect 23848 25842 23900 25848
rect 23204 25152 23256 25158
rect 23204 25094 23256 25100
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23216 24886 23244 25094
rect 23204 24880 23256 24886
rect 23204 24822 23256 24828
rect 23754 24848 23810 24857
rect 23112 24812 23164 24818
rect 23112 24754 23164 24760
rect 23572 24812 23624 24818
rect 23754 24783 23756 24792
rect 23572 24754 23624 24760
rect 23808 24783 23810 24792
rect 23756 24754 23808 24760
rect 23584 24698 23612 24754
rect 23400 24670 23612 24698
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23124 23254 23152 24550
rect 23400 23798 23428 24670
rect 23952 24426 23980 28630
rect 24044 25226 24072 30790
rect 24228 28422 24256 33866
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 24412 33525 24440 33594
rect 24387 33519 24440 33525
rect 24439 33476 24440 33519
rect 24387 33461 24439 33467
rect 24504 33318 24532 34410
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24596 33590 24624 33934
rect 24780 33658 24808 35866
rect 24872 34610 24900 36110
rect 24964 35834 24992 40054
rect 25976 39982 26004 40462
rect 25964 39976 26016 39982
rect 25964 39918 26016 39924
rect 25976 39302 26004 39918
rect 25964 39296 26016 39302
rect 25964 39238 26016 39244
rect 25976 38350 26004 39238
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 25964 38344 26016 38350
rect 25964 38286 26016 38292
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25148 36922 25176 37810
rect 25976 37806 26004 38286
rect 25964 37800 26016 37806
rect 25964 37742 26016 37748
rect 25976 37262 26004 37742
rect 25964 37256 26016 37262
rect 25964 37198 26016 37204
rect 25688 37120 25740 37126
rect 25688 37062 25740 37068
rect 25136 36916 25188 36922
rect 25136 36858 25188 36864
rect 25700 36786 25728 37062
rect 25504 36780 25556 36786
rect 25504 36722 25556 36728
rect 25688 36780 25740 36786
rect 25688 36722 25740 36728
rect 25516 36174 25544 36722
rect 25700 36242 25728 36722
rect 25688 36236 25740 36242
rect 25688 36178 25740 36184
rect 25504 36168 25556 36174
rect 25504 36110 25556 36116
rect 24952 35828 25004 35834
rect 24952 35770 25004 35776
rect 25688 35828 25740 35834
rect 25688 35770 25740 35776
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 24872 33862 24900 34546
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 24860 33856 24912 33862
rect 24860 33798 24912 33804
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24584 33584 24636 33590
rect 24584 33526 24636 33532
rect 24492 33312 24544 33318
rect 24492 33254 24544 33260
rect 24492 32904 24544 32910
rect 24596 32892 24624 33526
rect 24544 32864 24624 32892
rect 24492 32846 24544 32852
rect 24504 32570 24532 32846
rect 24492 32564 24544 32570
rect 24492 32506 24544 32512
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 24412 31346 24440 31622
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24412 30870 24440 31282
rect 24400 30864 24452 30870
rect 24400 30806 24452 30812
rect 24504 30734 24532 32506
rect 24676 32496 24728 32502
rect 24676 32438 24728 32444
rect 24688 31414 24716 32438
rect 24780 32348 24808 33594
rect 24872 32502 24900 33798
rect 24964 33658 24992 34002
rect 25056 33862 25084 34546
rect 25228 34400 25280 34406
rect 25228 34342 25280 34348
rect 25240 33998 25268 34342
rect 25207 33992 25268 33998
rect 25259 33952 25268 33992
rect 25207 33934 25259 33940
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 24952 33652 25004 33658
rect 24952 33594 25004 33600
rect 24860 32496 24912 32502
rect 24860 32438 24912 32444
rect 24860 32360 24912 32366
rect 24780 32320 24860 32348
rect 24860 32302 24912 32308
rect 24768 32224 24820 32230
rect 24768 32166 24820 32172
rect 24780 31822 24808 32166
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24688 30938 24716 31350
rect 24676 30932 24728 30938
rect 24676 30874 24728 30880
rect 24492 30728 24544 30734
rect 24492 30670 24544 30676
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24504 29646 24532 30670
rect 24584 30592 24636 30598
rect 24584 30534 24636 30540
rect 24596 30190 24624 30534
rect 24584 30184 24636 30190
rect 24584 30126 24636 30132
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24596 29578 24624 30126
rect 24584 29572 24636 29578
rect 24584 29514 24636 29520
rect 24688 28762 24716 30670
rect 24872 30258 24900 32302
rect 24952 31272 25004 31278
rect 24952 31214 25004 31220
rect 24964 30802 24992 31214
rect 24952 30796 25004 30802
rect 24952 30738 25004 30744
rect 25056 30326 25084 33798
rect 25136 33516 25188 33522
rect 25136 33458 25188 33464
rect 25148 33318 25176 33458
rect 25228 33380 25280 33386
rect 25228 33322 25280 33328
rect 25136 33312 25188 33318
rect 25136 33254 25188 33260
rect 25148 33114 25176 33254
rect 25136 33108 25188 33114
rect 25136 33050 25188 33056
rect 25148 31210 25176 33050
rect 25240 32978 25268 33322
rect 25228 32972 25280 32978
rect 25228 32914 25280 32920
rect 25240 32434 25268 32914
rect 25228 32428 25280 32434
rect 25228 32370 25280 32376
rect 25240 32337 25268 32370
rect 25226 32328 25282 32337
rect 25226 32263 25282 32272
rect 25700 31754 25728 35770
rect 26988 34950 27016 38694
rect 27264 36922 27292 40462
rect 27724 40186 27752 40530
rect 28448 40520 28500 40526
rect 28448 40462 28500 40468
rect 27712 40180 27764 40186
rect 27712 40122 27764 40128
rect 28460 40050 28488 40462
rect 29012 40446 29224 40474
rect 28908 40384 28960 40390
rect 29012 40372 29040 40446
rect 28960 40344 29040 40372
rect 29092 40384 29144 40390
rect 28908 40326 28960 40332
rect 29092 40326 29144 40332
rect 29000 40180 29052 40186
rect 29000 40122 29052 40128
rect 27712 40044 27764 40050
rect 27712 39986 27764 39992
rect 28448 40044 28500 40050
rect 28448 39986 28500 39992
rect 27724 39098 27752 39986
rect 27712 39092 27764 39098
rect 27712 39034 27764 39040
rect 28460 38962 28488 39986
rect 29012 38962 29040 40122
rect 28448 38956 28500 38962
rect 28448 38898 28500 38904
rect 29000 38956 29052 38962
rect 29000 38898 29052 38904
rect 28460 38758 28488 38898
rect 28448 38752 28500 38758
rect 29012 38740 29040 38898
rect 28448 38694 28500 38700
rect 28920 38712 29040 38740
rect 27712 38276 27764 38282
rect 27712 38218 27764 38224
rect 27724 36922 27752 38218
rect 27896 37188 27948 37194
rect 27896 37130 27948 37136
rect 27252 36916 27304 36922
rect 27252 36858 27304 36864
rect 27712 36916 27764 36922
rect 27712 36858 27764 36864
rect 27264 35894 27292 36858
rect 27908 36378 27936 37130
rect 28632 37120 28684 37126
rect 28632 37062 28684 37068
rect 28077 36780 28129 36786
rect 28077 36722 28129 36728
rect 27896 36372 27948 36378
rect 27896 36314 27948 36320
rect 28092 36310 28120 36722
rect 28264 36712 28316 36718
rect 28264 36654 28316 36660
rect 28172 36644 28224 36650
rect 28172 36586 28224 36592
rect 28080 36304 28132 36310
rect 28080 36246 28132 36252
rect 27804 36168 27856 36174
rect 27804 36110 27856 36116
rect 27620 36100 27672 36106
rect 27620 36042 27672 36048
rect 27172 35866 27292 35894
rect 27172 35290 27200 35866
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27344 35624 27396 35630
rect 27344 35566 27396 35572
rect 27160 35284 27212 35290
rect 27160 35226 27212 35232
rect 26976 34944 27028 34950
rect 26976 34886 27028 34892
rect 26240 34536 26292 34542
rect 26240 34478 26292 34484
rect 26252 31890 26280 34478
rect 26792 32224 26844 32230
rect 26792 32166 26844 32172
rect 26804 31890 26832 32166
rect 26240 31884 26292 31890
rect 26240 31826 26292 31832
rect 26792 31884 26844 31890
rect 26792 31826 26844 31832
rect 26516 31816 26568 31822
rect 26516 31758 26568 31764
rect 25700 31726 25820 31754
rect 25504 31476 25556 31482
rect 25504 31418 25556 31424
rect 25136 31204 25188 31210
rect 25136 31146 25188 31152
rect 25228 30728 25280 30734
rect 25228 30670 25280 30676
rect 25044 30320 25096 30326
rect 25044 30262 25096 30268
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24952 29640 25004 29646
rect 24952 29582 25004 29588
rect 24964 29306 24992 29582
rect 24952 29300 25004 29306
rect 24952 29242 25004 29248
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24676 28756 24728 28762
rect 24676 28698 24728 28704
rect 24780 28642 24808 29106
rect 25240 28694 25268 30670
rect 25516 29170 25544 31418
rect 25688 31204 25740 31210
rect 25688 31146 25740 31152
rect 25596 30592 25648 30598
rect 25596 30534 25648 30540
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 25516 28762 25544 29106
rect 25608 29034 25636 30534
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 24688 28614 24808 28642
rect 25228 28688 25280 28694
rect 25228 28630 25280 28636
rect 24688 28490 24716 28614
rect 25608 28558 25636 28970
rect 25596 28552 25648 28558
rect 25596 28494 25648 28500
rect 24676 28484 24728 28490
rect 24676 28426 24728 28432
rect 24216 28416 24268 28422
rect 24216 28358 24268 28364
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24124 27328 24176 27334
rect 24124 27270 24176 27276
rect 24136 27062 24164 27270
rect 24124 27056 24176 27062
rect 24124 26998 24176 27004
rect 24136 25945 24164 26998
rect 24216 26988 24268 26994
rect 24216 26930 24268 26936
rect 24228 26586 24256 26930
rect 24216 26580 24268 26586
rect 24216 26522 24268 26528
rect 24216 26308 24268 26314
rect 24216 26250 24268 26256
rect 24228 25974 24256 26250
rect 24216 25968 24268 25974
rect 24122 25936 24178 25945
rect 24216 25910 24268 25916
rect 24122 25871 24178 25880
rect 24032 25220 24084 25226
rect 24032 25162 24084 25168
rect 23584 24398 23980 24426
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23112 23248 23164 23254
rect 23112 23190 23164 23196
rect 22848 23072 22968 23100
rect 23032 23072 23152 23100
rect 22468 22228 22520 22234
rect 22468 22170 22520 22176
rect 22940 22094 22968 23072
rect 22940 22066 23060 22094
rect 22468 21344 22520 21350
rect 22468 21286 22520 21292
rect 22480 20942 22508 21286
rect 22468 20936 22520 20942
rect 22468 20878 22520 20884
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22480 17814 22508 18158
rect 22468 17808 22520 17814
rect 22468 17750 22520 17756
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22664 16590 22692 17138
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 16250 22692 16526
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22664 15502 22692 16186
rect 23032 15638 23060 22066
rect 23020 15632 23072 15638
rect 23020 15574 23072 15580
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 22928 15088 22980 15094
rect 22928 15030 22980 15036
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22664 14822 22692 14962
rect 22652 14816 22704 14822
rect 22652 14758 22704 14764
rect 22940 13530 22968 15030
rect 22928 13524 22980 13530
rect 23124 13512 23152 23072
rect 23400 22438 23428 23734
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23386 21992 23442 22001
rect 23386 21927 23442 21936
rect 23400 21894 23428 21927
rect 23388 21888 23440 21894
rect 23388 21830 23440 21836
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23492 20534 23520 21422
rect 23480 20528 23532 20534
rect 23480 20470 23532 20476
rect 23584 17490 23612 24398
rect 23848 22636 23900 22642
rect 23848 22578 23900 22584
rect 23860 21894 23888 22578
rect 24320 22094 24348 27814
rect 24688 27130 24716 28426
rect 25228 27668 25280 27674
rect 25228 27610 25280 27616
rect 24860 27396 24912 27402
rect 24860 27338 24912 27344
rect 24872 27130 24900 27338
rect 24676 27124 24728 27130
rect 24676 27066 24728 27072
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 24400 26988 24452 26994
rect 24768 26988 24820 26994
rect 24452 26948 24532 26976
rect 24400 26930 24452 26936
rect 24400 26308 24452 26314
rect 24400 26250 24452 26256
rect 24412 25906 24440 26250
rect 24400 25900 24452 25906
rect 24400 25842 24452 25848
rect 24412 23730 24440 25842
rect 24504 25838 24532 26948
rect 24768 26930 24820 26936
rect 24780 26330 24808 26930
rect 25044 26920 25096 26926
rect 25044 26862 25096 26868
rect 24596 26302 24808 26330
rect 24596 26234 24624 26302
rect 24596 26206 24808 26234
rect 24492 25832 24544 25838
rect 24492 25774 24544 25780
rect 24780 25294 24808 26206
rect 25056 25294 25084 26862
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 25044 25288 25096 25294
rect 25044 25230 25096 25236
rect 24584 25220 24636 25226
rect 24584 25162 24636 25168
rect 24596 24818 24624 25162
rect 24780 24954 24808 25230
rect 24964 24954 24992 25230
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24952 24948 25004 24954
rect 24952 24890 25004 24896
rect 24584 24812 24636 24818
rect 24584 24754 24636 24760
rect 24596 24410 24624 24754
rect 24584 24404 24636 24410
rect 24584 24346 24636 24352
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24504 23322 24532 23598
rect 24492 23316 24544 23322
rect 24492 23258 24544 23264
rect 24780 22710 24808 24890
rect 25056 24154 25084 25230
rect 24964 24126 25084 24154
rect 24768 22704 24820 22710
rect 24768 22646 24820 22652
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24228 22066 24348 22094
rect 23848 21888 23900 21894
rect 23848 21830 23900 21836
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23952 20466 23980 20742
rect 24136 20466 24164 20878
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23768 19854 23796 20198
rect 23756 19848 23808 19854
rect 23756 19790 23808 19796
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23676 17678 23704 18566
rect 23768 18290 23796 19790
rect 23952 18766 23980 20402
rect 24136 19786 24164 20402
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23940 18624 23992 18630
rect 23940 18566 23992 18572
rect 23952 18290 23980 18566
rect 24228 18426 24256 22066
rect 24872 21690 24900 22578
rect 24964 22506 24992 24126
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 25056 22642 25084 23258
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 24952 22500 25004 22506
rect 24952 22442 25004 22448
rect 25044 22500 25096 22506
rect 25044 22442 25096 22448
rect 24860 21684 24912 21690
rect 24860 21626 24912 21632
rect 24964 21486 24992 22442
rect 25056 21554 25084 22442
rect 25136 22432 25188 22438
rect 25136 22374 25188 22380
rect 25148 21570 25176 22374
rect 25240 21672 25268 27610
rect 25504 26988 25556 26994
rect 25504 26930 25556 26936
rect 25516 26586 25544 26930
rect 25504 26580 25556 26586
rect 25504 26522 25556 26528
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 25332 22001 25360 22374
rect 25318 21992 25374 22001
rect 25318 21927 25374 21936
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25516 21690 25544 21898
rect 25504 21684 25556 21690
rect 25240 21644 25360 21672
rect 25148 21554 25268 21570
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25148 21548 25280 21554
rect 25148 21542 25228 21548
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 25148 21146 25176 21542
rect 25228 21490 25280 21496
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 24308 18964 24360 18970
rect 24308 18906 24360 18912
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23940 18284 23992 18290
rect 23940 18226 23992 18232
rect 24216 17808 24268 17814
rect 24216 17750 24268 17756
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23584 17462 23704 17490
rect 23202 16688 23258 16697
rect 23202 16623 23204 16632
rect 23256 16623 23258 16632
rect 23204 16594 23256 16600
rect 23202 16144 23258 16153
rect 23202 16079 23258 16088
rect 23216 15706 23244 16079
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 23308 15586 23336 15642
rect 23216 15558 23336 15586
rect 23572 15564 23624 15570
rect 23216 15162 23244 15558
rect 23572 15506 23624 15512
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23388 15020 23440 15026
rect 23388 14962 23440 14968
rect 23204 14884 23256 14890
rect 23204 14826 23256 14832
rect 23216 14074 23244 14826
rect 23400 14550 23428 14962
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23308 14074 23336 14282
rect 23204 14068 23256 14074
rect 23204 14010 23256 14016
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 22928 13466 22980 13472
rect 23032 13484 23152 13512
rect 22468 13456 22520 13462
rect 22468 13398 22520 13404
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 21088 10736 21140 10742
rect 21088 10678 21140 10684
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19996 9042 20024 9522
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 8362 19196 8774
rect 19260 8401 19288 8910
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19352 8430 19380 8774
rect 19340 8424 19392 8430
rect 19246 8392 19302 8401
rect 19156 8356 19208 8362
rect 19340 8366 19392 8372
rect 19246 8327 19302 8336
rect 19156 8298 19208 8304
rect 19260 8022 19288 8327
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19248 7744 19300 7750
rect 19248 7686 19300 7692
rect 19260 6798 19288 7686
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19352 6254 19380 8366
rect 19444 7886 19472 8910
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19432 7880 19484 7886
rect 19536 7857 19564 8366
rect 19432 7822 19484 7828
rect 19522 7848 19578 7857
rect 19444 7546 19472 7822
rect 19522 7783 19578 7792
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19430 7440 19486 7449
rect 19430 7375 19486 7384
rect 19984 7404 20036 7410
rect 19444 7342 19472 7375
rect 19984 7346 20036 7352
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 18512 5840 18564 5846
rect 19076 5817 19104 6190
rect 19444 5914 19472 7278
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19996 6458 20024 7346
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 20088 6322 20116 10610
rect 20812 10056 20864 10062
rect 20812 9998 20864 10004
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 20088 6118 20116 6258
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 18512 5782 18564 5788
rect 19062 5808 19118 5817
rect 18524 5642 18552 5782
rect 19062 5743 19118 5752
rect 19340 5772 19392 5778
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18892 5030 18920 5170
rect 19076 5166 19104 5743
rect 19340 5714 19392 5720
rect 19352 5370 19380 5714
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5302 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19248 5296 19300 5302
rect 19248 5238 19300 5244
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19982 5264 20038 5273
rect 19064 5160 19116 5166
rect 19064 5102 19116 5108
rect 19260 5098 19288 5238
rect 19982 5199 19984 5208
rect 20036 5199 20038 5208
rect 19984 5170 20036 5176
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18880 5024 18932 5030
rect 18880 4966 18932 4972
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 18340 4758 18368 4966
rect 18328 4752 18380 4758
rect 18328 4694 18380 4700
rect 19168 4554 19196 4966
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19156 4548 19208 4554
rect 19156 4490 19208 4496
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 19352 4146 19380 4558
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 17316 2440 17368 2446
rect 17316 2382 17368 2388
rect 17224 2032 17276 2038
rect 17224 1974 17276 1980
rect 17328 800 17356 2382
rect 17604 800 17632 3470
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 17880 800 17908 2790
rect 18144 2508 18196 2514
rect 18144 2450 18196 2456
rect 18156 800 18184 2450
rect 18432 800 18460 3470
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18708 800 18736 2926
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 18984 800 19012 2314
rect 19260 800 19288 2790
rect 19444 1850 19472 3470
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19444 1822 19564 1850
rect 19536 800 19564 1822
rect 19996 1442 20024 2926
rect 20088 2774 20116 6054
rect 20180 5234 20208 9590
rect 20444 9512 20496 9518
rect 20444 9454 20496 9460
rect 20456 9042 20484 9454
rect 20444 9036 20496 9042
rect 20444 8978 20496 8984
rect 20720 8424 20772 8430
rect 20718 8392 20720 8401
rect 20772 8392 20774 8401
rect 20718 8327 20774 8336
rect 20824 7478 20852 9998
rect 21100 9926 21128 10678
rect 22008 10668 22060 10674
rect 22008 10610 22060 10616
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21928 10266 21956 10542
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21088 9920 21140 9926
rect 21088 9862 21140 9868
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8498 21220 8842
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 21284 7546 21312 8910
rect 22020 8906 22048 10610
rect 22296 10062 22324 10950
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 22112 8294 22140 9930
rect 22388 9722 22416 11290
rect 22480 10810 22508 13398
rect 23032 12374 23060 13484
rect 23020 12368 23072 12374
rect 23020 12310 23072 12316
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 22848 11898 22876 12242
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22572 10742 22600 11698
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 22560 10736 22612 10742
rect 22560 10678 22612 10684
rect 22572 10266 22600 10678
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22664 9976 22692 11154
rect 22848 11150 22876 11834
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 22928 11280 22980 11286
rect 22928 11222 22980 11228
rect 22836 11144 22888 11150
rect 22836 11086 22888 11092
rect 22940 10130 22968 11222
rect 23032 11150 23060 11494
rect 23020 11144 23072 11150
rect 23020 11086 23072 11092
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 22744 9988 22796 9994
rect 22664 9948 22744 9976
rect 22744 9930 22796 9936
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 23124 8634 23152 11834
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23388 11620 23440 11626
rect 23388 11562 23440 11568
rect 23400 11150 23428 11562
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23308 10538 23336 10610
rect 23296 10532 23348 10538
rect 23296 10474 23348 10480
rect 23204 9920 23256 9926
rect 23204 9862 23256 9868
rect 23216 9586 23244 9862
rect 23204 9580 23256 9586
rect 23204 9522 23256 9528
rect 23308 9382 23336 10474
rect 23400 9994 23428 11086
rect 23492 10810 23520 11698
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23216 8650 23244 9114
rect 23308 8974 23336 9318
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23112 8628 23164 8634
rect 23216 8622 23336 8650
rect 23112 8570 23164 8576
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22008 8288 22060 8294
rect 22008 8230 22060 8236
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20456 6322 20484 6598
rect 20732 6390 20760 7346
rect 20824 7002 20852 7414
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20456 5914 20484 6258
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20640 5710 20668 5741
rect 20628 5704 20680 5710
rect 20824 5658 20852 6938
rect 21284 6390 21312 7482
rect 22020 7002 22048 8230
rect 22572 7886 22600 8434
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 22560 7880 22612 7886
rect 22560 7822 22612 7828
rect 22572 7546 22600 7822
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 23216 7342 23244 8366
rect 23308 7750 23336 8622
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23492 7886 23520 8434
rect 23584 8090 23612 15506
rect 23676 15502 23704 17462
rect 24228 17338 24256 17750
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24124 17060 24176 17066
rect 24124 17002 24176 17008
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23664 15020 23716 15026
rect 23664 14962 23716 14968
rect 23676 14822 23704 14962
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23676 14414 23704 14758
rect 23860 14618 23888 14758
rect 23848 14612 23900 14618
rect 23848 14554 23900 14560
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 24044 10062 24072 10610
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23676 9722 23704 9998
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 24044 9466 24072 9998
rect 23952 9438 24072 9466
rect 23952 9110 23980 9438
rect 24032 9376 24084 9382
rect 24032 9318 24084 9324
rect 23940 9104 23992 9110
rect 23940 9046 23992 9052
rect 23952 8498 23980 9046
rect 24044 9042 24072 9318
rect 24136 9178 24164 17002
rect 24320 16454 24348 18906
rect 24768 18760 24820 18766
rect 24688 18720 24768 18748
rect 24688 18290 24716 18720
rect 24768 18702 24820 18708
rect 25044 18692 25096 18698
rect 25044 18634 25096 18640
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24412 17134 24440 17614
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24596 16794 24624 18022
rect 24688 17678 24716 18226
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 24964 16998 24992 18566
rect 25056 18426 25084 18634
rect 25044 18420 25096 18426
rect 25044 18362 25096 18368
rect 25332 17202 25360 21644
rect 25504 21626 25556 21632
rect 25596 21548 25648 21554
rect 25596 21490 25648 21496
rect 25608 21078 25636 21490
rect 25596 21072 25648 21078
rect 25596 21014 25648 21020
rect 25700 18442 25728 31146
rect 25792 29034 25820 31726
rect 26528 31686 26556 31758
rect 26516 31680 26568 31686
rect 26516 31622 26568 31628
rect 26528 31482 26556 31622
rect 26516 31476 26568 31482
rect 26516 31418 26568 31424
rect 26056 31272 26108 31278
rect 26056 31214 26108 31220
rect 26068 30938 26096 31214
rect 26056 30932 26108 30938
rect 26056 30874 26108 30880
rect 26804 30716 26832 31826
rect 26884 30728 26936 30734
rect 26804 30688 26884 30716
rect 26056 30320 26108 30326
rect 26056 30262 26108 30268
rect 25872 29504 25924 29510
rect 25872 29446 25924 29452
rect 25884 29238 25912 29446
rect 25872 29232 25924 29238
rect 25872 29174 25924 29180
rect 25780 29028 25832 29034
rect 25780 28970 25832 28976
rect 25792 26994 25820 28970
rect 25964 27396 26016 27402
rect 25964 27338 26016 27344
rect 25976 27130 26004 27338
rect 25964 27124 26016 27130
rect 25964 27066 26016 27072
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25792 26450 25820 26930
rect 25780 26444 25832 26450
rect 26068 26432 26096 30262
rect 26804 29578 26832 30688
rect 26884 30670 26936 30676
rect 26792 29572 26844 29578
rect 26792 29514 26844 29520
rect 26516 28620 26568 28626
rect 26516 28562 26568 28568
rect 26332 27328 26384 27334
rect 26332 27270 26384 27276
rect 25780 26386 25832 26392
rect 25976 26404 26096 26432
rect 25780 25152 25832 25158
rect 25780 25094 25832 25100
rect 25792 24886 25820 25094
rect 25780 24880 25832 24886
rect 25780 24822 25832 24828
rect 25792 21418 25820 24822
rect 25870 21992 25926 22001
rect 25870 21927 25926 21936
rect 25780 21412 25832 21418
rect 25780 21354 25832 21360
rect 25884 20874 25912 21927
rect 25872 20868 25924 20874
rect 25872 20810 25924 20816
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25792 18766 25820 19110
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25608 18414 25728 18442
rect 25320 17196 25372 17202
rect 25320 17138 25372 17144
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 24768 16992 24820 16998
rect 24768 16934 24820 16940
rect 24952 16992 25004 16998
rect 24952 16934 25004 16940
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24780 16658 24808 16934
rect 24492 16652 24544 16658
rect 24492 16594 24544 16600
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24308 16448 24360 16454
rect 24308 16390 24360 16396
rect 24504 16250 24532 16594
rect 24676 16584 24728 16590
rect 24676 16526 24728 16532
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 24492 16244 24544 16250
rect 24492 16186 24544 16192
rect 24584 14952 24636 14958
rect 24584 14894 24636 14900
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24504 14550 24532 14758
rect 24492 14544 24544 14550
rect 24492 14486 24544 14492
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24400 12368 24452 12374
rect 24400 12310 24452 12316
rect 24412 11354 24440 12310
rect 24504 11898 24532 14214
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24400 11348 24452 11354
rect 24400 11290 24452 11296
rect 24412 10674 24440 11290
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24032 9036 24084 9042
rect 24032 8978 24084 8984
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23308 7478 23336 7686
rect 23296 7472 23348 7478
rect 23492 7426 23520 7822
rect 24596 7546 24624 14894
rect 24688 13462 24716 16526
rect 25056 16046 25084 16526
rect 25044 16040 25096 16046
rect 25042 16008 25044 16017
rect 25096 16008 25098 16017
rect 25042 15943 25098 15952
rect 24952 15904 25004 15910
rect 24952 15846 25004 15852
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24676 13456 24728 13462
rect 24676 13398 24728 13404
rect 24780 12434 24808 15574
rect 24872 15026 24900 15642
rect 24964 15434 24992 15846
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 24688 12406 24808 12434
rect 24688 10470 24716 12406
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24676 10464 24728 10470
rect 24676 10406 24728 10412
rect 24688 10266 24716 10406
rect 24676 10260 24728 10266
rect 24676 10202 24728 10208
rect 24688 10062 24716 10202
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 24780 9586 24808 10746
rect 24964 10470 24992 15370
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25148 13258 25176 15030
rect 25240 14006 25268 17070
rect 25332 16794 25360 17138
rect 25320 16788 25372 16794
rect 25320 16730 25372 16736
rect 25608 15706 25636 18414
rect 25780 18352 25832 18358
rect 25780 18294 25832 18300
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25700 17882 25728 18226
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25792 17542 25820 18294
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25884 17134 25912 17614
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25688 15904 25740 15910
rect 25688 15846 25740 15852
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25700 15434 25728 15846
rect 25976 15706 26004 26404
rect 26148 26308 26200 26314
rect 26068 26268 26148 26296
rect 26068 25906 26096 26268
rect 26148 26250 26200 26256
rect 26344 25974 26372 27270
rect 26332 25968 26384 25974
rect 26332 25910 26384 25916
rect 26056 25900 26108 25906
rect 26056 25842 26108 25848
rect 26068 24818 26096 25842
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 26068 22642 26096 24754
rect 26528 24138 26556 28562
rect 26804 27538 26832 29514
rect 26792 27532 26844 27538
rect 26792 27474 26844 27480
rect 26988 25498 27016 34886
rect 27356 34542 27384 35566
rect 27448 35290 27476 35634
rect 27436 35284 27488 35290
rect 27436 35226 27488 35232
rect 27632 34678 27660 36042
rect 27816 36038 27844 36110
rect 27804 36032 27856 36038
rect 27724 35992 27804 36020
rect 27620 34672 27672 34678
rect 27620 34614 27672 34620
rect 27344 34536 27396 34542
rect 27344 34478 27396 34484
rect 27528 34536 27580 34542
rect 27528 34478 27580 34484
rect 27540 34066 27568 34478
rect 27528 34060 27580 34066
rect 27528 34002 27580 34008
rect 27344 33108 27396 33114
rect 27344 33050 27396 33056
rect 27356 32502 27384 33050
rect 27724 32774 27752 35992
rect 27804 35974 27856 35980
rect 28184 35834 28212 36586
rect 28276 36174 28304 36654
rect 28448 36236 28500 36242
rect 28448 36178 28500 36184
rect 28264 36168 28316 36174
rect 28264 36110 28316 36116
rect 28172 35828 28224 35834
rect 28172 35770 28224 35776
rect 28276 35714 28304 36110
rect 28092 35686 28304 35714
rect 28092 35086 28120 35686
rect 28264 35488 28316 35494
rect 28184 35436 28264 35442
rect 28184 35430 28316 35436
rect 28184 35414 28304 35430
rect 27988 35080 28040 35086
rect 27988 35022 28040 35028
rect 28080 35080 28132 35086
rect 28080 35022 28132 35028
rect 28000 34746 28028 35022
rect 27988 34740 28040 34746
rect 27988 34682 28040 34688
rect 28092 34678 28120 35022
rect 28080 34672 28132 34678
rect 28080 34614 28132 34620
rect 28184 34610 28212 35414
rect 28460 35154 28488 36178
rect 28540 36032 28592 36038
rect 28540 35974 28592 35980
rect 28552 35290 28580 35974
rect 28540 35284 28592 35290
rect 28540 35226 28592 35232
rect 28448 35148 28500 35154
rect 28448 35090 28500 35096
rect 28644 35018 28672 37062
rect 28632 35012 28684 35018
rect 28632 34954 28684 34960
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 27712 32768 27764 32774
rect 27712 32710 27764 32716
rect 27344 32496 27396 32502
rect 27344 32438 27396 32444
rect 27724 32026 27752 32710
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 27712 32020 27764 32026
rect 27712 31962 27764 31968
rect 26976 25492 27028 25498
rect 26976 25434 27028 25440
rect 26516 24132 26568 24138
rect 26516 24074 26568 24080
rect 27068 24132 27120 24138
rect 27068 24074 27120 24080
rect 26516 23588 26568 23594
rect 26516 23530 26568 23536
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26056 22636 26108 22642
rect 26056 22578 26108 22584
rect 26068 21622 26096 22578
rect 26344 22166 26372 22646
rect 26332 22160 26384 22166
rect 26332 22102 26384 22108
rect 26240 22024 26292 22030
rect 26240 21966 26292 21972
rect 26056 21616 26108 21622
rect 26056 21558 26108 21564
rect 26252 20942 26280 21966
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26252 19922 26280 20878
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 26068 17660 26096 18566
rect 26252 18306 26280 19858
rect 26252 18290 26372 18306
rect 26252 18284 26384 18290
rect 26252 18278 26332 18284
rect 26332 18226 26384 18232
rect 26528 17678 26556 23530
rect 27080 22506 27108 24074
rect 27068 22500 27120 22506
rect 27068 22442 27120 22448
rect 27068 22160 27120 22166
rect 27068 22102 27120 22108
rect 26700 21956 26752 21962
rect 26700 21898 26752 21904
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 26620 21554 26648 21830
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26240 17672 26292 17678
rect 26068 17632 26240 17660
rect 26240 17614 26292 17620
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26620 17490 26648 21490
rect 26528 17462 26648 17490
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26252 16114 26280 16730
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 25688 15428 25740 15434
rect 25688 15370 25740 15376
rect 25700 15026 25728 15370
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25332 14278 25360 14894
rect 25700 14346 25728 14962
rect 25976 14414 26004 15642
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 25964 14408 26016 14414
rect 25964 14350 26016 14356
rect 25688 14340 25740 14346
rect 25688 14282 25740 14288
rect 26056 14340 26108 14346
rect 26056 14282 26108 14288
rect 25320 14272 25372 14278
rect 25320 14214 25372 14220
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25148 12986 25176 13194
rect 25136 12980 25188 12986
rect 25136 12922 25188 12928
rect 25332 12434 25360 14214
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25608 13530 25636 13874
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25700 13258 25728 14282
rect 25964 14272 26016 14278
rect 25964 14214 26016 14220
rect 25976 13938 26004 14214
rect 26068 14074 26096 14282
rect 26056 14068 26108 14074
rect 26056 14010 26108 14016
rect 26344 13938 26372 14758
rect 25964 13932 26016 13938
rect 25964 13874 26016 13880
rect 26332 13932 26384 13938
rect 26332 13874 26384 13880
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25792 13326 25820 13670
rect 25780 13320 25832 13326
rect 25780 13262 25832 13268
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25872 13252 25924 13258
rect 25872 13194 25924 13200
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12918 25820 13126
rect 25780 12912 25832 12918
rect 25780 12854 25832 12860
rect 25148 12406 25360 12434
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 25044 9104 25096 9110
rect 25044 9046 25096 9052
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24688 8362 24716 8570
rect 25056 8566 25084 9046
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24780 7546 24808 8366
rect 24952 7812 25004 7818
rect 24952 7754 25004 7760
rect 24584 7540 24636 7546
rect 24584 7482 24636 7488
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 23296 7414 23348 7420
rect 23400 7410 23520 7426
rect 24860 7472 24912 7478
rect 24860 7414 24912 7420
rect 23388 7404 23520 7410
rect 23440 7398 23520 7404
rect 23664 7404 23716 7410
rect 23388 7346 23440 7352
rect 23664 7346 23716 7352
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24768 7404 24820 7410
rect 24768 7346 24820 7352
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23676 7274 23704 7346
rect 23480 7268 23532 7274
rect 23480 7210 23532 7216
rect 23664 7268 23716 7274
rect 23664 7210 23716 7216
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22204 6390 22232 6734
rect 21272 6384 21324 6390
rect 21272 6326 21324 6332
rect 22192 6384 22244 6390
rect 22192 6326 22244 6332
rect 20904 5840 20956 5846
rect 20904 5782 20956 5788
rect 20680 5652 20852 5658
rect 20628 5646 20852 5652
rect 20640 5630 20852 5646
rect 20168 5228 20220 5234
rect 20168 5170 20220 5176
rect 20260 5024 20312 5030
rect 20260 4966 20312 4972
rect 20272 4214 20300 4966
rect 20640 4622 20668 5630
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 20916 3942 20944 5782
rect 23492 5710 23520 7210
rect 24412 7206 24440 7346
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 24216 7200 24268 7206
rect 24216 7142 24268 7148
rect 24400 7200 24452 7206
rect 24400 7142 24452 7148
rect 23584 6322 23612 7142
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23480 5704 23532 5710
rect 23480 5646 23532 5652
rect 21272 5636 21324 5642
rect 21272 5578 21324 5584
rect 21284 4758 21312 5578
rect 23492 5370 23520 5646
rect 23480 5364 23532 5370
rect 23480 5306 23532 5312
rect 24228 5234 24256 7142
rect 24504 7002 24532 7346
rect 24492 6996 24544 7002
rect 24492 6938 24544 6944
rect 24780 5914 24808 7346
rect 24872 7274 24900 7414
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 24964 6458 24992 7754
rect 25148 7274 25176 12406
rect 25688 12096 25740 12102
rect 25884 12084 25912 13194
rect 25740 12056 25912 12084
rect 25688 12038 25740 12044
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25240 8498 25268 10542
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25332 9450 25360 9522
rect 25320 9444 25372 9450
rect 25320 9386 25372 9392
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25320 9172 25372 9178
rect 25320 9114 25372 9120
rect 25332 8838 25360 9114
rect 25320 8832 25372 8838
rect 25320 8774 25372 8780
rect 25424 8498 25452 9318
rect 25516 9110 25544 9522
rect 25504 9104 25556 9110
rect 25504 9046 25556 9052
rect 25516 8838 25544 9046
rect 25608 9042 25636 9590
rect 25596 9036 25648 9042
rect 25596 8978 25648 8984
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25240 8362 25268 8434
rect 25228 8356 25280 8362
rect 25228 8298 25280 8304
rect 25240 7410 25268 8298
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 25608 6662 25636 8978
rect 25700 8566 25728 12038
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25792 11150 25820 11698
rect 25780 11144 25832 11150
rect 25780 11086 25832 11092
rect 25872 8900 25924 8906
rect 25872 8842 25924 8848
rect 25884 8634 25912 8842
rect 25872 8628 25924 8634
rect 25872 8570 25924 8576
rect 25688 8560 25740 8566
rect 25688 8502 25740 8508
rect 25688 7812 25740 7818
rect 25688 7754 25740 7760
rect 25700 7478 25728 7754
rect 25976 7750 26004 13874
rect 26332 13728 26384 13734
rect 26332 13670 26384 13676
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 26252 13326 26280 13398
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 26344 12850 26372 13670
rect 26436 13462 26464 13874
rect 26424 13456 26476 13462
rect 26424 13398 26476 13404
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26148 9376 26200 9382
rect 26148 9318 26200 9324
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 25688 7472 25740 7478
rect 25688 7414 25740 7420
rect 26160 7410 26188 9318
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 26148 7404 26200 7410
rect 26148 7346 26200 7352
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 25608 6390 25636 6598
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 25596 6384 25648 6390
rect 25596 6326 25648 6332
rect 24768 5908 24820 5914
rect 24768 5850 24820 5856
rect 24872 5234 24900 6326
rect 25884 5710 25912 7346
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 26240 5704 26292 5710
rect 26240 5646 26292 5652
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 21272 4752 21324 4758
rect 21272 4694 21324 4700
rect 21284 4554 21312 4694
rect 21272 4548 21324 4554
rect 21272 4490 21324 4496
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 24872 3602 24900 5170
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24964 4622 24992 5102
rect 25780 5024 25832 5030
rect 25780 4966 25832 4972
rect 25792 4826 25820 4966
rect 25780 4820 25832 4826
rect 25780 4762 25832 4768
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 26056 4616 26108 4622
rect 26056 4558 26108 4564
rect 26068 3738 26096 4558
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 24860 3596 24912 3602
rect 24860 3538 24912 3544
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 21180 3528 21232 3534
rect 21180 3470 21232 3476
rect 22284 3528 22336 3534
rect 22284 3470 22336 3476
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 20088 2746 20208 2774
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 19812 1414 20024 1442
rect 19812 800 19840 1414
rect 20088 800 20116 2450
rect 20180 1970 20208 2746
rect 20168 1964 20220 1970
rect 20168 1906 20220 1912
rect 20364 800 20392 3470
rect 20536 2848 20588 2854
rect 20904 2848 20956 2854
rect 20588 2796 20668 2802
rect 20536 2790 20668 2796
rect 20904 2790 20956 2796
rect 20548 2774 20668 2790
rect 20640 800 20668 2774
rect 20916 800 20944 2790
rect 21192 800 21220 3470
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21468 800 21496 2586
rect 21744 800 21772 2790
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 22020 800 22048 2450
rect 22296 800 22324 3470
rect 22572 800 22600 3470
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 22836 2372 22888 2378
rect 22836 2314 22888 2320
rect 22848 800 22876 2314
rect 23124 800 23152 2790
rect 23400 800 23428 3470
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 24216 2848 24268 2854
rect 24216 2790 24268 2796
rect 23676 800 23704 2790
rect 23940 2372 23992 2378
rect 23940 2314 23992 2320
rect 23952 800 23980 2314
rect 24228 800 24256 2790
rect 24504 800 24532 3470
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24768 2440 24820 2446
rect 24768 2382 24820 2388
rect 24780 800 24808 2382
rect 25056 800 25084 2790
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 25332 800 25360 2450
rect 25608 800 25636 3470
rect 26252 3126 26280 5646
rect 26528 4622 26556 17462
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26620 16590 26648 17274
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26620 15502 26648 16526
rect 26608 15496 26660 15502
rect 26608 15438 26660 15444
rect 26620 14890 26648 15438
rect 26608 14884 26660 14890
rect 26608 14826 26660 14832
rect 26712 14385 26740 21898
rect 26976 21480 27028 21486
rect 26976 21422 27028 21428
rect 26988 21078 27016 21422
rect 26976 21072 27028 21078
rect 26976 21014 27028 21020
rect 27080 20942 27108 22102
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 26976 18692 27028 18698
rect 26976 18634 27028 18640
rect 26792 18624 26844 18630
rect 26792 18566 26844 18572
rect 26804 17660 26832 18566
rect 26988 18086 27016 18634
rect 27068 18284 27120 18290
rect 27068 18226 27120 18232
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 27080 17882 27108 18226
rect 27068 17876 27120 17882
rect 27068 17818 27120 17824
rect 26884 17672 26936 17678
rect 26804 17632 26884 17660
rect 26884 17614 26936 17620
rect 27172 17066 27200 31962
rect 27724 31822 27752 31962
rect 27712 31816 27764 31822
rect 27712 31758 27764 31764
rect 28184 30666 28212 34546
rect 28540 32836 28592 32842
rect 28540 32778 28592 32784
rect 28552 32570 28580 32778
rect 28540 32564 28592 32570
rect 28540 32506 28592 32512
rect 28264 32428 28316 32434
rect 28264 32370 28316 32376
rect 28276 32026 28304 32370
rect 28540 32292 28592 32298
rect 28540 32234 28592 32240
rect 28552 32026 28580 32234
rect 28264 32020 28316 32026
rect 28264 31962 28316 31968
rect 28540 32020 28592 32026
rect 28540 31962 28592 31968
rect 28448 31748 28500 31754
rect 28448 31690 28500 31696
rect 28172 30660 28224 30666
rect 28172 30602 28224 30608
rect 28460 27606 28488 31690
rect 28540 31340 28592 31346
rect 28540 31282 28592 31288
rect 28552 30734 28580 31282
rect 28540 30728 28592 30734
rect 28540 30670 28592 30676
rect 28552 30258 28580 30670
rect 28644 30326 28672 34954
rect 28724 32768 28776 32774
rect 28724 32710 28776 32716
rect 28736 31822 28764 32710
rect 28816 32564 28868 32570
rect 28816 32506 28868 32512
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 28724 31272 28776 31278
rect 28724 31214 28776 31220
rect 28736 30666 28764 31214
rect 28724 30660 28776 30666
rect 28724 30602 28776 30608
rect 28736 30326 28764 30602
rect 28632 30320 28684 30326
rect 28632 30262 28684 30268
rect 28724 30320 28776 30326
rect 28724 30262 28776 30268
rect 28828 30258 28856 32506
rect 28920 30734 28948 38712
rect 29000 38208 29052 38214
rect 29000 38150 29052 38156
rect 29012 35698 29040 38150
rect 29000 35692 29052 35698
rect 29000 35634 29052 35640
rect 29012 31482 29040 35634
rect 29104 33658 29132 40326
rect 29196 39914 29224 40446
rect 29184 39908 29236 39914
rect 29184 39850 29236 39856
rect 29288 39370 29316 40870
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 29920 40588 29972 40594
rect 29920 40530 29972 40536
rect 29552 40452 29604 40458
rect 29552 40394 29604 40400
rect 29564 39642 29592 40394
rect 29552 39636 29604 39642
rect 29552 39578 29604 39584
rect 29276 39364 29328 39370
rect 29276 39306 29328 39312
rect 29184 34740 29236 34746
rect 29184 34682 29236 34688
rect 29196 34202 29224 34682
rect 29184 34196 29236 34202
rect 29184 34138 29236 34144
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 29000 31136 29052 31142
rect 29000 31078 29052 31084
rect 28908 30728 28960 30734
rect 28908 30670 28960 30676
rect 28540 30252 28592 30258
rect 28540 30194 28592 30200
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 28448 27600 28500 27606
rect 28448 27542 28500 27548
rect 29012 27402 29040 31078
rect 29000 27396 29052 27402
rect 29000 27338 29052 27344
rect 29012 26994 29040 27338
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 28724 26784 28776 26790
rect 28724 26726 28776 26732
rect 27436 25968 27488 25974
rect 27436 25910 27488 25916
rect 27252 24608 27304 24614
rect 27252 24550 27304 24556
rect 27264 24274 27292 24550
rect 27252 24268 27304 24274
rect 27252 24210 27304 24216
rect 27344 23792 27396 23798
rect 27344 23734 27396 23740
rect 27356 22982 27384 23734
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27356 22778 27384 22918
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 27344 22432 27396 22438
rect 27344 22374 27396 22380
rect 27356 21690 27384 22374
rect 27344 21684 27396 21690
rect 27344 21626 27396 21632
rect 27448 21554 27476 25910
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 27632 24954 27660 25842
rect 27804 25764 27856 25770
rect 27804 25706 27856 25712
rect 27816 25226 27844 25706
rect 27896 25696 27948 25702
rect 27896 25638 27948 25644
rect 27804 25220 27856 25226
rect 27804 25162 27856 25168
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27804 24812 27856 24818
rect 27724 24772 27804 24800
rect 27724 24274 27752 24772
rect 27804 24754 27856 24760
rect 27804 24676 27856 24682
rect 27804 24618 27856 24624
rect 27712 24268 27764 24274
rect 27712 24210 27764 24216
rect 27816 24138 27844 24618
rect 27908 24206 27936 25638
rect 28540 25152 28592 25158
rect 28540 25094 28592 25100
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 28092 24410 28120 24754
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27620 24132 27672 24138
rect 27620 24074 27672 24080
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27632 23730 27660 24074
rect 27620 23724 27672 23730
rect 27620 23666 27672 23672
rect 27528 22500 27580 22506
rect 27528 22442 27580 22448
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27344 18352 27396 18358
rect 27344 18294 27396 18300
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 27264 17338 27292 17614
rect 27356 17542 27384 18294
rect 27448 17678 27476 18634
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27252 17332 27304 17338
rect 27304 17292 27384 17320
rect 27252 17274 27304 17280
rect 27160 17060 27212 17066
rect 27160 17002 27212 17008
rect 27160 14816 27212 14822
rect 27160 14758 27212 14764
rect 26698 14376 26754 14385
rect 26698 14311 26754 14320
rect 26712 11354 26740 14311
rect 27172 14006 27200 14758
rect 27160 14000 27212 14006
rect 27160 13942 27212 13948
rect 27172 13190 27200 13942
rect 27252 13296 27304 13302
rect 27252 13238 27304 13244
rect 27160 13184 27212 13190
rect 27160 13126 27212 13132
rect 27264 12646 27292 13238
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26712 10062 26740 11290
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 27160 8560 27212 8566
rect 27160 8502 27212 8508
rect 27172 8362 27200 8502
rect 27160 8356 27212 8362
rect 27160 8298 27212 8304
rect 27068 7880 27120 7886
rect 27068 7822 27120 7828
rect 26792 7472 26844 7478
rect 26792 7414 26844 7420
rect 26804 6798 26832 7414
rect 26792 6792 26844 6798
rect 26792 6734 26844 6740
rect 27080 6322 27108 7822
rect 27264 7002 27292 12582
rect 27356 12306 27384 17292
rect 27448 16794 27476 17614
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27448 14822 27476 15982
rect 27436 14816 27488 14822
rect 27436 14758 27488 14764
rect 27436 14340 27488 14346
rect 27436 14282 27488 14288
rect 27448 13326 27476 14282
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27344 9988 27396 9994
rect 27344 9930 27396 9936
rect 27356 9382 27384 9930
rect 27344 9376 27396 9382
rect 27344 9318 27396 9324
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 27448 8294 27476 8434
rect 27436 8288 27488 8294
rect 27436 8230 27488 8236
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 27540 6746 27568 22442
rect 27632 22094 27660 23666
rect 27712 23044 27764 23050
rect 27712 22986 27764 22992
rect 27724 22778 27752 22986
rect 27712 22772 27764 22778
rect 27712 22714 27764 22720
rect 27816 22574 27844 24074
rect 28172 23520 28224 23526
rect 28172 23462 28224 23468
rect 28184 22642 28212 23462
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 28276 22624 28304 24754
rect 28552 24138 28580 25094
rect 28632 24608 28684 24614
rect 28632 24550 28684 24556
rect 28644 24410 28672 24550
rect 28632 24404 28684 24410
rect 28632 24346 28684 24352
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28356 22636 28408 22642
rect 28276 22596 28356 22624
rect 27804 22568 27856 22574
rect 27804 22510 27856 22516
rect 27632 22066 27752 22094
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27632 17746 27660 19722
rect 27724 19514 27752 22066
rect 27712 19508 27764 19514
rect 27712 19450 27764 19456
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27632 14006 27660 17682
rect 27712 16788 27764 16794
rect 27712 16730 27764 16736
rect 27724 16590 27752 16730
rect 27816 16726 27844 22510
rect 28276 21962 28304 22596
rect 28356 22578 28408 22584
rect 28356 22228 28408 22234
rect 28356 22170 28408 22176
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28080 21888 28132 21894
rect 28080 21830 28132 21836
rect 28092 20942 28120 21830
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28184 20942 28212 21422
rect 28368 21146 28396 22170
rect 28540 21412 28592 21418
rect 28540 21354 28592 21360
rect 28552 21146 28580 21354
rect 28356 21140 28408 21146
rect 28356 21082 28408 21088
rect 28540 21140 28592 21146
rect 28540 21082 28592 21088
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 28172 20936 28224 20942
rect 28172 20878 28224 20884
rect 28184 20398 28212 20878
rect 28172 20392 28224 20398
rect 28172 20334 28224 20340
rect 28184 18834 28212 20334
rect 28172 18828 28224 18834
rect 28172 18770 28224 18776
rect 27896 18352 27948 18358
rect 27896 18294 27948 18300
rect 27804 16720 27856 16726
rect 27804 16662 27856 16668
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27908 16114 27936 18294
rect 27988 17604 28040 17610
rect 27988 17546 28040 17552
rect 28000 16697 28028 17546
rect 27986 16688 28042 16697
rect 27986 16623 28042 16632
rect 27896 16108 27948 16114
rect 27896 16050 27948 16056
rect 27908 15706 27936 16050
rect 27896 15700 27948 15706
rect 27896 15642 27948 15648
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27620 14000 27672 14006
rect 27620 13942 27672 13948
rect 27620 12232 27672 12238
rect 27620 12174 27672 12180
rect 27632 11898 27660 12174
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27632 10810 27660 11834
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27264 6718 27568 6746
rect 27068 6316 27120 6322
rect 27068 6258 27120 6264
rect 27160 6316 27212 6322
rect 27160 6258 27212 6264
rect 26976 6248 27028 6254
rect 26976 6190 27028 6196
rect 26988 5778 27016 6190
rect 27172 5914 27200 6258
rect 27160 5908 27212 5914
rect 27160 5850 27212 5856
rect 26976 5772 27028 5778
rect 26976 5714 27028 5720
rect 26988 5534 27016 5714
rect 27264 5710 27292 6718
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27448 5710 27476 6598
rect 27252 5704 27304 5710
rect 27252 5646 27304 5652
rect 27436 5704 27488 5710
rect 27436 5646 27488 5652
rect 27160 5636 27212 5642
rect 27160 5578 27212 5584
rect 26896 5506 27016 5534
rect 26896 4622 26924 5506
rect 27172 5166 27200 5578
rect 27160 5160 27212 5166
rect 27160 5102 27212 5108
rect 27172 4758 27200 5102
rect 27436 5092 27488 5098
rect 27436 5034 27488 5040
rect 27160 4752 27212 4758
rect 27160 4694 27212 4700
rect 27172 4622 27200 4694
rect 26516 4616 26568 4622
rect 26516 4558 26568 4564
rect 26884 4616 26936 4622
rect 26884 4558 26936 4564
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 26332 4480 26384 4486
rect 26332 4422 26384 4428
rect 26344 3534 26372 4422
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26240 3120 26292 3126
rect 26240 3062 26292 3068
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 25884 800 25912 2790
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26160 800 26188 2382
rect 26436 800 26464 2926
rect 26976 2848 27028 2854
rect 26976 2790 27028 2796
rect 26700 2508 26752 2514
rect 26700 2450 26752 2456
rect 26712 800 26740 2450
rect 26988 800 27016 2790
rect 27448 2582 27476 5034
rect 27632 4690 27660 10610
rect 27712 10124 27764 10130
rect 27712 10066 27764 10072
rect 27724 9042 27752 10066
rect 27816 9450 27844 14554
rect 28000 14414 28028 15302
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28356 14816 28408 14822
rect 28356 14758 28408 14764
rect 28080 14544 28132 14550
rect 28080 14486 28132 14492
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 28092 13326 28120 14486
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28276 14278 28304 14350
rect 28368 14346 28396 14758
rect 28356 14340 28408 14346
rect 28356 14282 28408 14288
rect 28264 14272 28316 14278
rect 28264 14214 28316 14220
rect 28276 13462 28304 14214
rect 28264 13456 28316 13462
rect 28264 13398 28316 13404
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 28080 12980 28132 12986
rect 28080 12922 28132 12928
rect 27896 10600 27948 10606
rect 27896 10542 27948 10548
rect 27908 9466 27936 10542
rect 28092 9722 28120 12922
rect 28080 9716 28132 9722
rect 28080 9658 28132 9664
rect 27988 9512 28040 9518
rect 27908 9460 27988 9466
rect 27908 9454 28040 9460
rect 27804 9444 27856 9450
rect 27804 9386 27856 9392
rect 27908 9438 28028 9454
rect 27908 9330 27936 9438
rect 27816 9302 27936 9330
rect 27712 9036 27764 9042
rect 27712 8978 27764 8984
rect 27816 8974 27844 9302
rect 27804 8968 27856 8974
rect 27804 8910 27856 8916
rect 27988 8968 28040 8974
rect 27988 8910 28040 8916
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27724 7818 27752 8298
rect 27712 7812 27764 7818
rect 27712 7754 27764 7760
rect 27816 7546 27844 8434
rect 27908 8362 27936 8570
rect 28000 8430 28028 8910
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 27896 8356 27948 8362
rect 27896 8298 27948 8304
rect 28092 8294 28120 9658
rect 28276 9178 28304 13398
rect 28368 13326 28396 14282
rect 28460 13734 28488 14894
rect 28552 14618 28580 14962
rect 28540 14612 28592 14618
rect 28540 14554 28592 14560
rect 28448 13728 28500 13734
rect 28448 13670 28500 13676
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28552 12986 28580 13262
rect 28540 12980 28592 12986
rect 28540 12922 28592 12928
rect 28644 11898 28672 24346
rect 28736 17814 28764 26726
rect 28816 25832 28868 25838
rect 28816 25774 28868 25780
rect 28828 25362 28856 25774
rect 28816 25356 28868 25362
rect 28816 25298 28868 25304
rect 28828 23186 28856 25298
rect 28908 25288 28960 25294
rect 28908 25230 28960 25236
rect 28920 24818 28948 25230
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28920 23730 28948 24754
rect 29104 24721 29132 33594
rect 29288 31346 29316 39306
rect 29932 38962 29960 40530
rect 58164 40520 58216 40526
rect 58164 40462 58216 40468
rect 30288 40452 30340 40458
rect 30288 40394 30340 40400
rect 30012 40384 30064 40390
rect 30012 40326 30064 40332
rect 30024 40050 30052 40326
rect 30300 40186 30328 40394
rect 31852 40384 31904 40390
rect 31852 40326 31904 40332
rect 30288 40180 30340 40186
rect 30288 40122 30340 40128
rect 31864 40118 31892 40326
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 58176 40225 58204 40462
rect 58162 40216 58218 40225
rect 58162 40151 58218 40160
rect 31852 40112 31904 40118
rect 31852 40054 31904 40060
rect 30012 40044 30064 40050
rect 30012 39986 30064 39992
rect 31208 40044 31260 40050
rect 31208 39986 31260 39992
rect 30104 39908 30156 39914
rect 30104 39850 30156 39856
rect 29920 38956 29972 38962
rect 29920 38898 29972 38904
rect 30116 38826 30144 39850
rect 30380 39296 30432 39302
rect 30380 39238 30432 39244
rect 30392 39030 30420 39238
rect 31220 39030 31248 39986
rect 31760 39432 31812 39438
rect 31760 39374 31812 39380
rect 31668 39296 31720 39302
rect 31668 39238 31720 39244
rect 30380 39024 30432 39030
rect 30380 38966 30432 38972
rect 31208 39024 31260 39030
rect 31208 38966 31260 38972
rect 30472 38956 30524 38962
rect 30472 38898 30524 38904
rect 30104 38820 30156 38826
rect 30104 38762 30156 38768
rect 30116 38282 30144 38762
rect 30484 38554 30512 38898
rect 31116 38752 31168 38758
rect 31116 38694 31168 38700
rect 30472 38548 30524 38554
rect 30472 38490 30524 38496
rect 31128 38350 31156 38694
rect 31116 38344 31168 38350
rect 31116 38286 31168 38292
rect 30104 38276 30156 38282
rect 30104 38218 30156 38224
rect 29920 38208 29972 38214
rect 29920 38150 29972 38156
rect 29828 37664 29880 37670
rect 29828 37606 29880 37612
rect 29552 35692 29604 35698
rect 29552 35634 29604 35640
rect 29564 35086 29592 35634
rect 29736 35148 29788 35154
rect 29736 35090 29788 35096
rect 29552 35080 29604 35086
rect 29552 35022 29604 35028
rect 29564 34678 29592 35022
rect 29552 34672 29604 34678
rect 29552 34614 29604 34620
rect 29644 33924 29696 33930
rect 29644 33866 29696 33872
rect 29656 33658 29684 33866
rect 29748 33658 29776 35090
rect 29840 34542 29868 37606
rect 29932 35086 29960 38150
rect 30116 36106 30144 38218
rect 31128 37874 31156 38286
rect 31220 38282 31248 38966
rect 31680 38962 31708 39238
rect 31668 38956 31720 38962
rect 31668 38898 31720 38904
rect 31680 38486 31708 38898
rect 31668 38480 31720 38486
rect 31668 38422 31720 38428
rect 31208 38276 31260 38282
rect 31208 38218 31260 38224
rect 31116 37868 31168 37874
rect 31116 37810 31168 37816
rect 30104 36100 30156 36106
rect 30104 36042 30156 36048
rect 30932 36100 30984 36106
rect 30932 36042 30984 36048
rect 31116 36100 31168 36106
rect 31116 36042 31168 36048
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29932 34746 29960 35022
rect 29920 34740 29972 34746
rect 29920 34682 29972 34688
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 29644 33652 29696 33658
rect 29644 33594 29696 33600
rect 29736 33652 29788 33658
rect 29736 33594 29788 33600
rect 29840 31754 29868 34478
rect 30116 31890 30144 36042
rect 30840 36032 30892 36038
rect 30840 35974 30892 35980
rect 30472 35624 30524 35630
rect 30472 35566 30524 35572
rect 30288 35216 30340 35222
rect 30288 35158 30340 35164
rect 30300 34066 30328 35158
rect 30288 34060 30340 34066
rect 30288 34002 30340 34008
rect 30484 32910 30512 35566
rect 30564 35080 30616 35086
rect 30564 35022 30616 35028
rect 30576 34542 30604 35022
rect 30852 35018 30880 35974
rect 30944 35290 30972 36042
rect 31128 35698 31156 36042
rect 31116 35692 31168 35698
rect 31116 35634 31168 35640
rect 30932 35284 30984 35290
rect 30932 35226 30984 35232
rect 30840 35012 30892 35018
rect 30840 34954 30892 34960
rect 30564 34536 30616 34542
rect 30564 34478 30616 34484
rect 30576 33522 30604 34478
rect 30564 33516 30616 33522
rect 30564 33458 30616 33464
rect 30472 32904 30524 32910
rect 30472 32846 30524 32852
rect 30564 32904 30616 32910
rect 30564 32846 30616 32852
rect 30380 32020 30432 32026
rect 30380 31962 30432 31968
rect 30104 31884 30156 31890
rect 30104 31826 30156 31832
rect 29828 31748 29880 31754
rect 29828 31690 29880 31696
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 29840 31142 29868 31690
rect 30392 31482 30420 31962
rect 30380 31476 30432 31482
rect 30380 31418 30432 31424
rect 29828 31136 29880 31142
rect 29828 31078 29880 31084
rect 30392 30734 30420 31418
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30380 30320 30432 30326
rect 30380 30262 30432 30268
rect 29920 30252 29972 30258
rect 29920 30194 29972 30200
rect 29828 30116 29880 30122
rect 29828 30058 29880 30064
rect 29552 30048 29604 30054
rect 29552 29990 29604 29996
rect 29564 29850 29592 29990
rect 29552 29844 29604 29850
rect 29552 29786 29604 29792
rect 29564 28762 29592 29786
rect 29840 29170 29868 30058
rect 29828 29164 29880 29170
rect 29828 29106 29880 29112
rect 29552 28756 29604 28762
rect 29552 28698 29604 28704
rect 29276 28688 29328 28694
rect 29276 28630 29328 28636
rect 29090 24712 29146 24721
rect 29090 24647 29146 24656
rect 28908 23724 28960 23730
rect 28908 23666 28960 23672
rect 28816 23180 28868 23186
rect 28816 23122 28868 23128
rect 29288 22778 29316 28630
rect 29840 28558 29868 29106
rect 29828 28552 29880 28558
rect 29828 28494 29880 28500
rect 29368 27328 29420 27334
rect 29368 27270 29420 27276
rect 29552 27328 29604 27334
rect 29552 27270 29604 27276
rect 29380 26314 29408 27270
rect 29368 26308 29420 26314
rect 29368 26250 29420 26256
rect 29380 25106 29408 26250
rect 29564 25226 29592 27270
rect 29840 26994 29868 28494
rect 29932 28082 29960 30194
rect 30392 29510 30420 30262
rect 30380 29504 30432 29510
rect 30380 29446 30432 29452
rect 30392 29170 30420 29446
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30104 28960 30156 28966
rect 30104 28902 30156 28908
rect 29920 28076 29972 28082
rect 29920 28018 29972 28024
rect 29828 26988 29880 26994
rect 29828 26930 29880 26936
rect 29644 26240 29696 26246
rect 29644 26182 29696 26188
rect 29656 25906 29684 26182
rect 29644 25900 29696 25906
rect 29644 25842 29696 25848
rect 29828 25900 29880 25906
rect 29828 25842 29880 25848
rect 29656 25378 29684 25842
rect 29840 25498 29868 25842
rect 29920 25764 29972 25770
rect 29920 25706 29972 25712
rect 29828 25492 29880 25498
rect 29828 25434 29880 25440
rect 29656 25350 29776 25378
rect 29932 25362 29960 25706
rect 29748 25294 29776 25350
rect 29920 25356 29972 25362
rect 29920 25298 29972 25304
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 30012 25288 30064 25294
rect 30012 25230 30064 25236
rect 29552 25220 29604 25226
rect 29552 25162 29604 25168
rect 29380 25078 29684 25106
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29276 22772 29328 22778
rect 29104 22732 29276 22760
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 29012 20874 29040 21626
rect 29000 20868 29052 20874
rect 29000 20810 29052 20816
rect 29012 20398 29040 20810
rect 29000 20392 29052 20398
rect 29000 20334 29052 20340
rect 29012 18902 29040 20334
rect 29000 18896 29052 18902
rect 29000 18838 29052 18844
rect 28724 17808 28776 17814
rect 28724 17750 28776 17756
rect 28724 15428 28776 15434
rect 28724 15370 28776 15376
rect 28736 14346 28764 15370
rect 28724 14340 28776 14346
rect 28724 14282 28776 14288
rect 28724 13728 28776 13734
rect 28724 13670 28776 13676
rect 28632 11892 28684 11898
rect 28632 11834 28684 11840
rect 28736 11762 28764 13670
rect 29104 12434 29132 22732
rect 29276 22714 29328 22720
rect 29276 22500 29328 22506
rect 29276 22442 29328 22448
rect 29184 21956 29236 21962
rect 29184 21898 29236 21904
rect 29012 12406 29132 12434
rect 28816 12164 28868 12170
rect 28816 12106 28868 12112
rect 28724 11756 28776 11762
rect 28724 11698 28776 11704
rect 28828 11694 28856 12106
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 28632 11280 28684 11286
rect 28632 11222 28684 11228
rect 28644 10742 28672 11222
rect 28724 11076 28776 11082
rect 28724 11018 28776 11024
rect 28632 10736 28684 10742
rect 28632 10678 28684 10684
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28552 8498 28580 9862
rect 28632 9172 28684 9178
rect 28632 9114 28684 9120
rect 28644 8634 28672 9114
rect 28632 8628 28684 8634
rect 28632 8570 28684 8576
rect 28540 8492 28592 8498
rect 28540 8434 28592 8440
rect 28080 8288 28132 8294
rect 28080 8230 28132 8236
rect 28736 8090 28764 11018
rect 29012 10690 29040 12406
rect 29196 10810 29224 21898
rect 29288 15706 29316 22442
rect 29564 22166 29592 23258
rect 29368 22160 29420 22166
rect 29368 22102 29420 22108
rect 29552 22160 29604 22166
rect 29552 22102 29604 22108
rect 29380 21690 29408 22102
rect 29656 22094 29684 25078
rect 29748 24410 29776 25230
rect 30024 24954 30052 25230
rect 30012 24948 30064 24954
rect 30012 24890 30064 24896
rect 29828 24608 29880 24614
rect 30116 24562 30144 28902
rect 30576 28762 30604 32846
rect 30944 30802 30972 35226
rect 31128 33930 31156 35634
rect 31220 35630 31248 38218
rect 31208 35624 31260 35630
rect 31208 35566 31260 35572
rect 31576 35624 31628 35630
rect 31576 35566 31628 35572
rect 31588 34610 31616 35566
rect 31576 34604 31628 34610
rect 31576 34546 31628 34552
rect 31116 33924 31168 33930
rect 31116 33866 31168 33872
rect 31128 33046 31156 33866
rect 31484 33856 31536 33862
rect 31484 33798 31536 33804
rect 31208 33652 31260 33658
rect 31208 33594 31260 33600
rect 31220 33318 31248 33594
rect 31208 33312 31260 33318
rect 31208 33254 31260 33260
rect 31116 33040 31168 33046
rect 31116 32982 31168 32988
rect 31300 31952 31352 31958
rect 31300 31894 31352 31900
rect 31116 31680 31168 31686
rect 31116 31622 31168 31628
rect 30932 30796 30984 30802
rect 30932 30738 30984 30744
rect 30944 30394 30972 30738
rect 30932 30388 30984 30394
rect 30932 30330 30984 30336
rect 30944 30122 30972 30330
rect 30932 30116 30984 30122
rect 30932 30058 30984 30064
rect 30654 28928 30710 28937
rect 30654 28863 30710 28872
rect 30564 28756 30616 28762
rect 30564 28698 30616 28704
rect 30564 28008 30616 28014
rect 30564 27950 30616 27956
rect 30380 27396 30432 27402
rect 30380 27338 30432 27344
rect 30392 26042 30420 27338
rect 30576 27130 30604 27950
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30380 26036 30432 26042
rect 30380 25978 30432 25984
rect 30196 25900 30248 25906
rect 30196 25842 30248 25848
rect 30208 25702 30236 25842
rect 30380 25764 30432 25770
rect 30380 25706 30432 25712
rect 30196 25696 30248 25702
rect 30196 25638 30248 25644
rect 29828 24550 29880 24556
rect 29736 24404 29788 24410
rect 29736 24346 29788 24352
rect 29840 24070 29868 24550
rect 30024 24534 30144 24562
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 29840 23798 29868 24006
rect 29828 23792 29880 23798
rect 29828 23734 29880 23740
rect 29656 22066 29776 22094
rect 29368 21684 29420 21690
rect 29368 21626 29420 21632
rect 29748 21554 29776 22066
rect 29920 22092 29972 22098
rect 30024 22094 30052 24534
rect 30104 24404 30156 24410
rect 30104 24346 30156 24352
rect 30116 24206 30144 24346
rect 30104 24200 30156 24206
rect 30104 24142 30156 24148
rect 30208 23746 30236 25638
rect 30392 25294 30420 25706
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30300 23866 30328 24142
rect 30288 23860 30340 23866
rect 30288 23802 30340 23808
rect 30208 23718 30328 23746
rect 30300 22982 30328 23718
rect 30288 22976 30340 22982
rect 30288 22918 30340 22924
rect 30300 22506 30328 22918
rect 30288 22500 30340 22506
rect 30288 22442 30340 22448
rect 30392 22098 30420 25230
rect 30564 25152 30616 25158
rect 30564 25094 30616 25100
rect 30576 24818 30604 25094
rect 30564 24812 30616 24818
rect 30564 24754 30616 24760
rect 30024 22066 30236 22094
rect 29920 22034 29972 22040
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 29736 20800 29788 20806
rect 29736 20742 29788 20748
rect 29552 20528 29604 20534
rect 29552 20470 29604 20476
rect 29564 19378 29592 20470
rect 29748 20466 29776 20742
rect 29736 20460 29788 20466
rect 29736 20402 29788 20408
rect 29748 19446 29776 20402
rect 29736 19440 29788 19446
rect 29736 19382 29788 19388
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29552 19372 29604 19378
rect 29552 19314 29604 19320
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29472 14414 29500 19314
rect 29564 18902 29592 19314
rect 29644 19168 29696 19174
rect 29644 19110 29696 19116
rect 29552 18896 29604 18902
rect 29552 18838 29604 18844
rect 29656 18086 29684 19110
rect 29748 18766 29776 19382
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 29828 18692 29880 18698
rect 29828 18634 29880 18640
rect 29736 18216 29788 18222
rect 29736 18158 29788 18164
rect 29644 18080 29696 18086
rect 29644 18022 29696 18028
rect 29552 17060 29604 17066
rect 29552 17002 29604 17008
rect 29564 16658 29592 17002
rect 29552 16652 29604 16658
rect 29552 16594 29604 16600
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 29552 14000 29604 14006
rect 29552 13942 29604 13948
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29288 13530 29316 13874
rect 29564 13530 29592 13942
rect 29276 13524 29328 13530
rect 29276 13466 29328 13472
rect 29552 13524 29604 13530
rect 29552 13466 29604 13472
rect 29368 12776 29420 12782
rect 29368 12718 29420 12724
rect 29184 10804 29236 10810
rect 29184 10746 29236 10752
rect 29012 10662 29224 10690
rect 28908 9512 28960 9518
rect 28908 9454 28960 9460
rect 28920 8566 28948 9454
rect 29000 8900 29052 8906
rect 29000 8842 29052 8848
rect 29012 8634 29040 8842
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 28908 8560 28960 8566
rect 28908 8502 28960 8508
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 28736 7410 28764 8026
rect 28724 7404 28776 7410
rect 28724 7346 28776 7352
rect 28828 6798 28856 8434
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28828 6458 28856 6734
rect 29196 6662 29224 10662
rect 29380 10198 29408 12718
rect 29460 12640 29512 12646
rect 29460 12582 29512 12588
rect 29472 11830 29500 12582
rect 29460 11824 29512 11830
rect 29460 11766 29512 11772
rect 29748 11354 29776 18158
rect 29840 15502 29868 18634
rect 29932 17542 29960 22034
rect 30208 21622 30236 22066
rect 30380 22092 30432 22098
rect 30668 22094 30696 28863
rect 30748 28484 30800 28490
rect 30748 28426 30800 28432
rect 30760 23118 30788 28426
rect 30840 24812 30892 24818
rect 30840 24754 30892 24760
rect 30852 24410 30880 24754
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 30748 23112 30800 23118
rect 30748 23054 30800 23060
rect 30668 22066 30788 22094
rect 30380 22034 30432 22040
rect 30656 22024 30708 22030
rect 30656 21966 30708 21972
rect 30196 21616 30248 21622
rect 30196 21558 30248 21564
rect 30288 21616 30340 21622
rect 30288 21558 30340 21564
rect 30012 21480 30064 21486
rect 30012 21422 30064 21428
rect 29920 17536 29972 17542
rect 29920 17478 29972 17484
rect 29920 16652 29972 16658
rect 29920 16594 29972 16600
rect 29828 15496 29880 15502
rect 29828 15438 29880 15444
rect 29840 15162 29868 15438
rect 29828 15156 29880 15162
rect 29828 15098 29880 15104
rect 29932 15042 29960 16594
rect 29840 15014 29960 15042
rect 29736 11348 29788 11354
rect 29736 11290 29788 11296
rect 29460 11144 29512 11150
rect 29460 11086 29512 11092
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29368 10192 29420 10198
rect 29368 10134 29420 10140
rect 29276 6724 29328 6730
rect 29276 6666 29328 6672
rect 29184 6656 29236 6662
rect 29184 6598 29236 6604
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 29288 6390 29316 6666
rect 29276 6384 29328 6390
rect 29276 6326 29328 6332
rect 29288 5710 29316 6326
rect 29276 5704 29328 5710
rect 29276 5646 29328 5652
rect 29288 4690 29316 5646
rect 27620 4684 27672 4690
rect 27620 4626 27672 4632
rect 29276 4684 29328 4690
rect 29276 4626 29328 4632
rect 27632 3738 27660 4626
rect 29288 4486 29316 4626
rect 29000 4480 29052 4486
rect 29000 4422 29052 4428
rect 29276 4480 29328 4486
rect 29276 4422 29328 4428
rect 29012 4282 29040 4422
rect 29000 4276 29052 4282
rect 29000 4218 29052 4224
rect 27620 3732 27672 3738
rect 27620 3674 27672 3680
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 27264 800 27292 2382
rect 27540 800 27568 3470
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27816 800 27844 2790
rect 28092 800 28120 2790
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28368 800 28396 2518
rect 28644 800 28672 3470
rect 29012 2961 29040 4218
rect 29472 3942 29500 11086
rect 29748 10674 29776 11086
rect 29552 10668 29604 10674
rect 29552 10610 29604 10616
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29564 10062 29592 10610
rect 29748 10130 29776 10610
rect 29736 10124 29788 10130
rect 29736 10066 29788 10072
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29564 8498 29592 9998
rect 29840 9058 29868 15014
rect 29920 14272 29972 14278
rect 29920 14214 29972 14220
rect 29932 13394 29960 14214
rect 29920 13388 29972 13394
rect 29920 13330 29972 13336
rect 29920 12844 29972 12850
rect 29920 12786 29972 12792
rect 29932 12442 29960 12786
rect 29920 12436 29972 12442
rect 29920 12378 29972 12384
rect 29748 9030 29868 9058
rect 29552 8492 29604 8498
rect 29552 8434 29604 8440
rect 29748 5098 29776 9030
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29840 7886 29868 8910
rect 30024 8634 30052 21422
rect 30196 21140 30248 21146
rect 30196 21082 30248 21088
rect 30104 21072 30156 21078
rect 30104 21014 30156 21020
rect 30116 20942 30144 21014
rect 30208 20942 30236 21082
rect 30300 21010 30328 21558
rect 30288 21004 30340 21010
rect 30288 20946 30340 20952
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 30196 20936 30248 20942
rect 30196 20878 30248 20884
rect 30116 20534 30144 20878
rect 30104 20528 30156 20534
rect 30104 20470 30156 20476
rect 30288 19236 30340 19242
rect 30288 19178 30340 19184
rect 30300 17882 30328 19178
rect 30472 18624 30524 18630
rect 30472 18566 30524 18572
rect 30484 17882 30512 18566
rect 30288 17876 30340 17882
rect 30288 17818 30340 17824
rect 30472 17876 30524 17882
rect 30472 17818 30524 17824
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 30380 16040 30432 16046
rect 30380 15982 30432 15988
rect 30392 15502 30420 15982
rect 30380 15496 30432 15502
rect 30380 15438 30432 15444
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30300 13938 30328 14350
rect 30288 13932 30340 13938
rect 30288 13874 30340 13880
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 30116 13258 30144 13466
rect 30104 13252 30156 13258
rect 30104 13194 30156 13200
rect 30116 10810 30144 13194
rect 30392 12850 30420 15438
rect 30484 15162 30512 15438
rect 30472 15156 30524 15162
rect 30472 15098 30524 15104
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 30392 12714 30420 12786
rect 30380 12708 30432 12714
rect 30380 12650 30432 12656
rect 30472 12164 30524 12170
rect 30472 12106 30524 12112
rect 30484 11082 30512 12106
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 30472 11076 30524 11082
rect 30472 11018 30524 11024
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30392 10742 30420 11018
rect 30380 10736 30432 10742
rect 30380 10678 30432 10684
rect 30392 9586 30420 10678
rect 30576 10538 30604 17614
rect 30564 10532 30616 10538
rect 30564 10474 30616 10480
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30012 8628 30064 8634
rect 30012 8570 30064 8576
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 29840 7206 29868 7822
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 30196 7200 30248 7206
rect 30196 7142 30248 7148
rect 30208 6798 30236 7142
rect 30196 6792 30248 6798
rect 30196 6734 30248 6740
rect 30012 6316 30064 6322
rect 30012 6258 30064 6264
rect 30024 5234 30052 6258
rect 30012 5228 30064 5234
rect 30012 5170 30064 5176
rect 29736 5092 29788 5098
rect 29736 5034 29788 5040
rect 30024 4622 30052 5170
rect 30012 4616 30064 4622
rect 30012 4558 30064 4564
rect 30208 4146 30236 6734
rect 30564 6656 30616 6662
rect 30564 6598 30616 6604
rect 30576 6322 30604 6598
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30472 6180 30524 6186
rect 30472 6122 30524 6128
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30392 5370 30420 5510
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 30288 5160 30340 5166
rect 30484 5148 30512 6122
rect 30340 5120 30512 5148
rect 30288 5102 30340 5108
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 30392 4282 30420 4558
rect 30484 4554 30512 5120
rect 30576 5030 30604 6258
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 30564 4752 30616 4758
rect 30564 4694 30616 4700
rect 30472 4548 30524 4554
rect 30472 4490 30524 4496
rect 30380 4276 30432 4282
rect 30380 4218 30432 4224
rect 30576 4214 30604 4694
rect 30668 4622 30696 21966
rect 30760 17678 30788 22066
rect 31024 22092 31076 22098
rect 31024 22034 31076 22040
rect 30840 20868 30892 20874
rect 30840 20810 30892 20816
rect 30852 19854 30880 20810
rect 30840 19848 30892 19854
rect 30892 19808 30972 19836
rect 30840 19790 30892 19796
rect 30840 19712 30892 19718
rect 30840 19654 30892 19660
rect 30852 19378 30880 19654
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 30944 18970 30972 19808
rect 31036 19378 31064 22034
rect 31128 22030 31156 31622
rect 31208 30728 31260 30734
rect 31208 30670 31260 30676
rect 31220 30394 31248 30670
rect 31208 30388 31260 30394
rect 31208 30330 31260 30336
rect 31312 22094 31340 31894
rect 31496 31822 31524 33798
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31484 30728 31536 30734
rect 31484 30670 31536 30676
rect 31496 29782 31524 30670
rect 31588 30666 31616 34546
rect 31680 32774 31708 38422
rect 31772 36650 31800 39374
rect 31760 36644 31812 36650
rect 31760 36586 31812 36592
rect 31864 36530 31892 40054
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 33324 39432 33376 39438
rect 33324 39374 33376 39380
rect 32128 39364 32180 39370
rect 32128 39306 32180 39312
rect 32140 39098 32168 39306
rect 33232 39296 33284 39302
rect 33232 39238 33284 39244
rect 32128 39092 32180 39098
rect 32128 39034 32180 39040
rect 33140 39024 33192 39030
rect 33140 38966 33192 38972
rect 32588 38956 32640 38962
rect 32588 38898 32640 38904
rect 31944 38752 31996 38758
rect 31944 38694 31996 38700
rect 31956 38282 31984 38694
rect 32600 38554 32628 38898
rect 32588 38548 32640 38554
rect 32588 38490 32640 38496
rect 33152 38418 33180 38966
rect 33140 38412 33192 38418
rect 33140 38354 33192 38360
rect 33244 38350 33272 39238
rect 33232 38344 33284 38350
rect 33232 38286 33284 38292
rect 31944 38276 31996 38282
rect 31944 38218 31996 38224
rect 32680 38276 32732 38282
rect 32680 38218 32732 38224
rect 32312 37800 32364 37806
rect 32312 37742 32364 37748
rect 32324 37466 32352 37742
rect 32312 37460 32364 37466
rect 32312 37402 32364 37408
rect 32036 36644 32088 36650
rect 32036 36586 32088 36592
rect 31772 36502 31892 36530
rect 31668 32768 31720 32774
rect 31668 32710 31720 32716
rect 31680 32026 31708 32710
rect 31772 32434 31800 36502
rect 32048 36106 32076 36586
rect 32036 36100 32088 36106
rect 32036 36042 32088 36048
rect 31852 33380 31904 33386
rect 31852 33322 31904 33328
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 31760 31952 31812 31958
rect 31760 31894 31812 31900
rect 31772 31793 31800 31894
rect 31758 31784 31814 31793
rect 31758 31719 31814 31728
rect 31864 30682 31892 33322
rect 32048 33114 32076 36042
rect 32404 36032 32456 36038
rect 32404 35974 32456 35980
rect 32416 34950 32444 35974
rect 32404 34944 32456 34950
rect 32404 34886 32456 34892
rect 32036 33108 32088 33114
rect 32036 33050 32088 33056
rect 31944 32768 31996 32774
rect 31944 32710 31996 32716
rect 31956 32570 31984 32710
rect 31944 32564 31996 32570
rect 31944 32506 31996 32512
rect 31944 32428 31996 32434
rect 31944 32370 31996 32376
rect 31956 31822 31984 32370
rect 31944 31816 31996 31822
rect 31944 31758 31996 31764
rect 31576 30660 31628 30666
rect 31576 30602 31628 30608
rect 31772 30654 31892 30682
rect 31588 30258 31616 30602
rect 31576 30252 31628 30258
rect 31576 30194 31628 30200
rect 31772 30054 31800 30654
rect 31852 30592 31904 30598
rect 31852 30534 31904 30540
rect 31760 30048 31812 30054
rect 31760 29990 31812 29996
rect 31484 29776 31536 29782
rect 31484 29718 31536 29724
rect 31392 27464 31444 27470
rect 31392 27406 31444 27412
rect 31404 26926 31432 27406
rect 31496 27130 31524 29718
rect 31576 29640 31628 29646
rect 31576 29582 31628 29588
rect 31588 27538 31616 29582
rect 31772 29306 31800 29990
rect 31864 29646 31892 30534
rect 31852 29640 31904 29646
rect 31852 29582 31904 29588
rect 31760 29300 31812 29306
rect 31760 29242 31812 29248
rect 31772 27606 31800 29242
rect 32048 28762 32076 33050
rect 32128 32768 32180 32774
rect 32128 32710 32180 32716
rect 32036 28756 32088 28762
rect 32036 28698 32088 28704
rect 31760 27600 31812 27606
rect 31760 27542 31812 27548
rect 31576 27532 31628 27538
rect 31576 27474 31628 27480
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31588 27062 31616 27474
rect 31576 27056 31628 27062
rect 31576 26998 31628 27004
rect 31392 26920 31444 26926
rect 31392 26862 31444 26868
rect 31588 26586 31616 26998
rect 32140 26874 32168 32710
rect 32220 32224 32272 32230
rect 32220 32166 32272 32172
rect 31864 26846 32168 26874
rect 31576 26580 31628 26586
rect 31576 26522 31628 26528
rect 31588 25974 31616 26522
rect 31576 25968 31628 25974
rect 31576 25910 31628 25916
rect 31588 25294 31616 25910
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 31588 24818 31616 25230
rect 31576 24812 31628 24818
rect 31576 24754 31628 24760
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31772 24206 31800 24346
rect 31760 24200 31812 24206
rect 31760 24142 31812 24148
rect 31668 23044 31720 23050
rect 31668 22986 31720 22992
rect 31680 22506 31708 22986
rect 31668 22500 31720 22506
rect 31668 22442 31720 22448
rect 31220 22066 31340 22094
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 31128 21078 31156 21490
rect 31116 21072 31168 21078
rect 31116 21014 31168 21020
rect 31128 20942 31156 21014
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31116 19780 31168 19786
rect 31116 19722 31168 19728
rect 31024 19372 31076 19378
rect 31024 19314 31076 19320
rect 30932 18964 30984 18970
rect 30932 18906 30984 18912
rect 31128 17814 31156 19722
rect 31220 18290 31248 22066
rect 31576 20528 31628 20534
rect 31576 20470 31628 20476
rect 31208 18284 31260 18290
rect 31208 18226 31260 18232
rect 31116 17808 31168 17814
rect 31116 17750 31168 17756
rect 30748 17672 30800 17678
rect 30748 17614 30800 17620
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30760 15094 30788 16050
rect 31300 15360 31352 15366
rect 31300 15302 31352 15308
rect 30748 15088 30800 15094
rect 30748 15030 30800 15036
rect 30760 12170 30788 15030
rect 31312 15026 31340 15302
rect 31300 15020 31352 15026
rect 31300 14962 31352 14968
rect 31116 13728 31168 13734
rect 31116 13670 31168 13676
rect 31128 12918 31156 13670
rect 31116 12912 31168 12918
rect 31116 12854 31168 12860
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 31208 12844 31260 12850
rect 31208 12786 31260 12792
rect 30840 12232 30892 12238
rect 30840 12174 30892 12180
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30748 6724 30800 6730
rect 30748 6666 30800 6672
rect 30760 6458 30788 6666
rect 30748 6452 30800 6458
rect 30748 6394 30800 6400
rect 30852 5914 30880 12174
rect 30840 5908 30892 5914
rect 30840 5850 30892 5856
rect 30840 5636 30892 5642
rect 30840 5578 30892 5584
rect 30852 5370 30880 5578
rect 30840 5364 30892 5370
rect 30840 5306 30892 5312
rect 30944 4622 30972 12786
rect 31220 12102 31248 12786
rect 31208 12096 31260 12102
rect 31208 12038 31260 12044
rect 31220 11762 31248 12038
rect 31312 11830 31340 14962
rect 31588 12986 31616 20470
rect 31680 19242 31708 22442
rect 31864 20874 31892 26846
rect 31944 24200 31996 24206
rect 31944 24142 31996 24148
rect 31956 23594 31984 24142
rect 31944 23588 31996 23594
rect 31944 23530 31996 23536
rect 31956 23118 31984 23530
rect 31944 23112 31996 23118
rect 31944 23054 31996 23060
rect 32128 23112 32180 23118
rect 32128 23054 32180 23060
rect 31956 22642 31984 23054
rect 32140 22778 32168 23054
rect 32128 22772 32180 22778
rect 32128 22714 32180 22720
rect 32036 22704 32088 22710
rect 32036 22646 32088 22652
rect 31944 22636 31996 22642
rect 31944 22578 31996 22584
rect 31944 21888 31996 21894
rect 31944 21830 31996 21836
rect 31956 21690 31984 21830
rect 31944 21684 31996 21690
rect 31944 21626 31996 21632
rect 32048 21622 32076 22646
rect 32126 21856 32182 21865
rect 32126 21791 32182 21800
rect 32140 21690 32168 21791
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 32232 21622 32260 32166
rect 32312 31816 32364 31822
rect 32416 31804 32444 34886
rect 32496 33856 32548 33862
rect 32496 33798 32548 33804
rect 32508 33590 32536 33798
rect 32496 33584 32548 33590
rect 32496 33526 32548 33532
rect 32588 32904 32640 32910
rect 32588 32846 32640 32852
rect 32600 32434 32628 32846
rect 32588 32428 32640 32434
rect 32588 32370 32640 32376
rect 32600 31890 32628 32370
rect 32692 31890 32720 38218
rect 33140 36100 33192 36106
rect 33140 36042 33192 36048
rect 33152 35834 33180 36042
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 33048 35692 33100 35698
rect 33048 35634 33100 35640
rect 33060 35494 33088 35634
rect 33140 35624 33192 35630
rect 33140 35566 33192 35572
rect 33048 35488 33100 35494
rect 33048 35430 33100 35436
rect 33060 32910 33088 35430
rect 33152 34746 33180 35566
rect 33140 34740 33192 34746
rect 33140 34682 33192 34688
rect 33048 32904 33100 32910
rect 33048 32846 33100 32852
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 32864 32836 32916 32842
rect 32864 32778 32916 32784
rect 32876 32450 32904 32778
rect 33152 32502 33180 32846
rect 32784 32434 32904 32450
rect 33140 32496 33192 32502
rect 33140 32438 33192 32444
rect 32772 32428 32904 32434
rect 32824 32422 32904 32428
rect 32772 32370 32824 32376
rect 32588 31884 32640 31890
rect 32588 31826 32640 31832
rect 32680 31884 32732 31890
rect 32680 31826 32732 31832
rect 32496 31816 32548 31822
rect 32416 31776 32496 31804
rect 32312 31758 32364 31764
rect 32496 31758 32548 31764
rect 32324 31346 32352 31758
rect 32784 31754 32812 32370
rect 32680 31748 32812 31754
rect 32732 31726 32812 31748
rect 32680 31690 32732 31696
rect 32692 31346 32720 31690
rect 33244 31346 33272 38286
rect 33336 36378 33364 39374
rect 34520 39296 34572 39302
rect 34520 39238 34572 39244
rect 34532 38962 34560 39238
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 33508 38956 33560 38962
rect 34520 38956 34572 38962
rect 33560 38916 33640 38944
rect 33508 38898 33560 38904
rect 33508 38480 33560 38486
rect 33508 38422 33560 38428
rect 33416 38276 33468 38282
rect 33416 38218 33468 38224
rect 33428 37942 33456 38218
rect 33416 37936 33468 37942
rect 33416 37878 33468 37884
rect 33428 36786 33456 37878
rect 33416 36780 33468 36786
rect 33416 36722 33468 36728
rect 33324 36372 33376 36378
rect 33324 36314 33376 36320
rect 33336 35766 33364 36314
rect 33324 35760 33376 35766
rect 33324 35702 33376 35708
rect 33336 35154 33364 35702
rect 33428 35630 33456 36722
rect 33520 36242 33548 38422
rect 33612 38282 33640 38916
rect 34520 38898 34572 38904
rect 35348 38956 35400 38962
rect 35400 38916 35480 38944
rect 35348 38898 35400 38904
rect 34796 38888 34848 38894
rect 34796 38830 34848 38836
rect 34704 38752 34756 38758
rect 34704 38694 34756 38700
rect 33692 38344 33744 38350
rect 33692 38286 33744 38292
rect 34520 38344 34572 38350
rect 34520 38286 34572 38292
rect 33600 38276 33652 38282
rect 33600 38218 33652 38224
rect 33612 37738 33640 38218
rect 33704 38010 33732 38286
rect 34060 38208 34112 38214
rect 34060 38150 34112 38156
rect 33692 38004 33744 38010
rect 33692 37946 33744 37952
rect 34072 37874 34100 38150
rect 34060 37868 34112 37874
rect 34060 37810 34112 37816
rect 33600 37732 33652 37738
rect 33600 37674 33652 37680
rect 33508 36236 33560 36242
rect 33508 36178 33560 36184
rect 33416 35624 33468 35630
rect 33416 35566 33468 35572
rect 33520 35154 33548 36178
rect 33612 36174 33640 37674
rect 33784 36576 33836 36582
rect 33784 36518 33836 36524
rect 33600 36168 33652 36174
rect 33600 36110 33652 36116
rect 33324 35148 33376 35154
rect 33324 35090 33376 35096
rect 33508 35148 33560 35154
rect 33508 35090 33560 35096
rect 33520 34678 33548 35090
rect 33508 34672 33560 34678
rect 33508 34614 33560 34620
rect 33612 34610 33640 36110
rect 33796 34610 33824 36518
rect 33600 34604 33652 34610
rect 33600 34546 33652 34552
rect 33784 34604 33836 34610
rect 33784 34546 33836 34552
rect 33416 34536 33468 34542
rect 33416 34478 33468 34484
rect 33428 33862 33456 34478
rect 33416 33856 33468 33862
rect 33416 33798 33468 33804
rect 33428 33658 33456 33798
rect 33416 33652 33468 33658
rect 33416 33594 33468 33600
rect 32312 31340 32364 31346
rect 32312 31282 32364 31288
rect 32680 31340 32732 31346
rect 32680 31282 32732 31288
rect 33232 31340 33284 31346
rect 33232 31282 33284 31288
rect 32324 30802 32352 31282
rect 32312 30796 32364 30802
rect 32312 30738 32364 30744
rect 32496 30728 32548 30734
rect 32496 30670 32548 30676
rect 32508 29170 32536 30670
rect 32692 30258 32720 31282
rect 32864 31136 32916 31142
rect 32864 31078 32916 31084
rect 32680 30252 32732 30258
rect 32680 30194 32732 30200
rect 32496 29164 32548 29170
rect 32496 29106 32548 29112
rect 32508 28558 32536 29106
rect 32588 28756 32640 28762
rect 32588 28698 32640 28704
rect 32496 28552 32548 28558
rect 32496 28494 32548 28500
rect 32508 28082 32536 28494
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32416 27674 32444 27814
rect 32404 27668 32456 27674
rect 32404 27610 32456 27616
rect 32508 27538 32536 28018
rect 32600 27946 32628 28698
rect 32588 27940 32640 27946
rect 32588 27882 32640 27888
rect 32496 27532 32548 27538
rect 32496 27474 32548 27480
rect 32600 26586 32628 27882
rect 32772 27532 32824 27538
rect 32772 27474 32824 27480
rect 32784 27441 32812 27474
rect 32770 27432 32826 27441
rect 32770 27367 32826 27376
rect 32588 26580 32640 26586
rect 32588 26522 32640 26528
rect 32600 26382 32628 26522
rect 32588 26376 32640 26382
rect 32588 26318 32640 26324
rect 32772 24268 32824 24274
rect 32772 24210 32824 24216
rect 32312 23520 32364 23526
rect 32312 23462 32364 23468
rect 32324 22710 32352 23462
rect 32784 23186 32812 24210
rect 32772 23180 32824 23186
rect 32772 23122 32824 23128
rect 32496 23044 32548 23050
rect 32496 22986 32548 22992
rect 32508 22710 32536 22986
rect 32312 22704 32364 22710
rect 32312 22646 32364 22652
rect 32496 22704 32548 22710
rect 32496 22646 32548 22652
rect 32508 22094 32536 22646
rect 32508 22066 32628 22094
rect 32600 21962 32628 22066
rect 32588 21956 32640 21962
rect 32588 21898 32640 21904
rect 32036 21616 32088 21622
rect 31942 21584 31998 21593
rect 32036 21558 32088 21564
rect 32220 21616 32272 21622
rect 32220 21558 32272 21564
rect 31942 21519 31998 21528
rect 32312 21548 32364 21554
rect 31956 21078 31984 21519
rect 32312 21490 32364 21496
rect 32036 21480 32088 21486
rect 32036 21422 32088 21428
rect 31944 21072 31996 21078
rect 31944 21014 31996 21020
rect 31760 20868 31812 20874
rect 31760 20810 31812 20816
rect 31852 20868 31904 20874
rect 31852 20810 31904 20816
rect 31772 19854 31800 20810
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31944 19440 31996 19446
rect 31944 19382 31996 19388
rect 31668 19236 31720 19242
rect 31668 19178 31720 19184
rect 31680 18698 31708 19178
rect 31956 18766 31984 19382
rect 31944 18760 31996 18766
rect 31944 18702 31996 18708
rect 31668 18692 31720 18698
rect 31668 18634 31720 18640
rect 31680 18222 31708 18634
rect 31668 18216 31720 18222
rect 31668 18158 31720 18164
rect 32048 16946 32076 21422
rect 32220 21344 32272 21350
rect 32220 21286 32272 21292
rect 32232 21078 32260 21286
rect 32324 21146 32352 21490
rect 32312 21140 32364 21146
rect 32312 21082 32364 21088
rect 32220 21072 32272 21078
rect 32220 21014 32272 21020
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32128 19304 32180 19310
rect 32128 19246 32180 19252
rect 31772 16918 32076 16946
rect 31576 12980 31628 12986
rect 31576 12922 31628 12928
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 31404 12238 31432 12786
rect 31392 12232 31444 12238
rect 31392 12174 31444 12180
rect 31300 11824 31352 11830
rect 31300 11766 31352 11772
rect 31404 11762 31432 12174
rect 31772 11898 31800 16918
rect 32036 16108 32088 16114
rect 32036 16050 32088 16056
rect 31852 15972 31904 15978
rect 31852 15914 31904 15920
rect 31864 15570 31892 15914
rect 31852 15564 31904 15570
rect 31852 15506 31904 15512
rect 31864 13002 31892 15506
rect 32048 14822 32076 16050
rect 32036 14816 32088 14822
rect 32036 14758 32088 14764
rect 31864 12974 31984 13002
rect 31956 12918 31984 12974
rect 31852 12912 31904 12918
rect 31852 12854 31904 12860
rect 31944 12912 31996 12918
rect 31944 12854 31996 12860
rect 31864 12102 31892 12854
rect 32048 12170 32076 14758
rect 32140 13530 32168 19246
rect 32128 13524 32180 13530
rect 32128 13466 32180 13472
rect 32140 12850 32168 13466
rect 32128 12844 32180 12850
rect 32128 12786 32180 12792
rect 32232 12374 32260 20878
rect 32312 20800 32364 20806
rect 32312 20742 32364 20748
rect 32324 20262 32352 20742
rect 32312 20256 32364 20262
rect 32312 20198 32364 20204
rect 32600 19786 32628 21898
rect 32680 19848 32732 19854
rect 32680 19790 32732 19796
rect 32784 19802 32812 23122
rect 32876 20534 32904 31078
rect 32956 30320 33008 30326
rect 32956 30262 33008 30268
rect 32968 29850 32996 30262
rect 33612 30258 33640 34546
rect 33692 30932 33744 30938
rect 33692 30874 33744 30880
rect 33704 30326 33732 30874
rect 33968 30660 34020 30666
rect 33968 30602 34020 30608
rect 33692 30320 33744 30326
rect 33692 30262 33744 30268
rect 33600 30252 33652 30258
rect 33600 30194 33652 30200
rect 33048 30184 33100 30190
rect 33048 30126 33100 30132
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32968 28082 32996 29786
rect 33060 29102 33088 30126
rect 33876 29572 33928 29578
rect 33876 29514 33928 29520
rect 33888 29238 33916 29514
rect 33876 29232 33928 29238
rect 33876 29174 33928 29180
rect 33048 29096 33100 29102
rect 33048 29038 33100 29044
rect 33980 29050 34008 30602
rect 34072 29170 34100 37810
rect 34532 37670 34560 38286
rect 34716 37874 34744 38694
rect 34808 38010 34836 38830
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 34796 38004 34848 38010
rect 34796 37946 34848 37952
rect 34704 37868 34756 37874
rect 34704 37810 34756 37816
rect 34520 37664 34572 37670
rect 34520 37606 34572 37612
rect 34520 36780 34572 36786
rect 34520 36722 34572 36728
rect 34532 35494 34560 36722
rect 34612 36032 34664 36038
rect 34612 35974 34664 35980
rect 34624 35698 34652 35974
rect 34612 35692 34664 35698
rect 34612 35634 34664 35640
rect 34520 35488 34572 35494
rect 34520 35430 34572 35436
rect 34532 32434 34560 35430
rect 34520 32428 34572 32434
rect 34520 32370 34572 32376
rect 34520 30728 34572 30734
rect 34520 30670 34572 30676
rect 34336 30592 34388 30598
rect 34336 30534 34388 30540
rect 34244 30320 34296 30326
rect 34244 30262 34296 30268
rect 34060 29164 34112 29170
rect 34060 29106 34112 29112
rect 33784 29028 33836 29034
rect 33980 29022 34100 29050
rect 34256 29034 34284 30262
rect 34348 30258 34376 30534
rect 34336 30252 34388 30258
rect 34336 30194 34388 30200
rect 33784 28970 33836 28976
rect 33416 28688 33468 28694
rect 33692 28688 33744 28694
rect 33468 28636 33692 28642
rect 33416 28630 33744 28636
rect 33428 28614 33732 28630
rect 33796 28490 33824 28970
rect 33784 28484 33836 28490
rect 33784 28426 33836 28432
rect 33692 28416 33744 28422
rect 33692 28358 33744 28364
rect 33416 28144 33468 28150
rect 33416 28086 33468 28092
rect 32956 28076 33008 28082
rect 32956 28018 33008 28024
rect 33232 27532 33284 27538
rect 33232 27474 33284 27480
rect 33140 27464 33192 27470
rect 33140 27406 33192 27412
rect 33152 27130 33180 27406
rect 33244 27334 33272 27474
rect 33428 27470 33456 28086
rect 33508 27872 33560 27878
rect 33508 27814 33560 27820
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 33232 27328 33284 27334
rect 33232 27270 33284 27276
rect 33416 27328 33468 27334
rect 33416 27270 33468 27276
rect 33140 27124 33192 27130
rect 33140 27066 33192 27072
rect 33428 26994 33456 27270
rect 33416 26988 33468 26994
rect 33416 26930 33468 26936
rect 33520 24970 33548 27814
rect 33428 24942 33548 24970
rect 33048 24676 33100 24682
rect 33048 24618 33100 24624
rect 33060 24138 33088 24618
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33048 24132 33100 24138
rect 33048 24074 33100 24080
rect 32864 20528 32916 20534
rect 32864 20470 32916 20476
rect 32588 19780 32640 19786
rect 32588 19722 32640 19728
rect 32692 19514 32720 19790
rect 32784 19774 32996 19802
rect 32864 19712 32916 19718
rect 32864 19654 32916 19660
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32324 18766 32352 19314
rect 32772 18828 32824 18834
rect 32772 18770 32824 18776
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 32324 14550 32352 18702
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 32600 16658 32628 18362
rect 32588 16652 32640 16658
rect 32588 16594 32640 16600
rect 32600 16114 32628 16594
rect 32588 16108 32640 16114
rect 32588 16050 32640 16056
rect 32784 15502 32812 18770
rect 32876 18766 32904 19654
rect 32864 18760 32916 18766
rect 32864 18702 32916 18708
rect 32864 16992 32916 16998
rect 32864 16934 32916 16940
rect 32876 16658 32904 16934
rect 32864 16652 32916 16658
rect 32864 16594 32916 16600
rect 32772 15496 32824 15502
rect 32772 15438 32824 15444
rect 32784 15094 32812 15438
rect 32772 15088 32824 15094
rect 32772 15030 32824 15036
rect 32312 14544 32364 14550
rect 32312 14486 32364 14492
rect 32324 14006 32352 14486
rect 32312 14000 32364 14006
rect 32312 13942 32364 13948
rect 32772 13320 32824 13326
rect 32772 13262 32824 13268
rect 32784 12986 32812 13262
rect 32772 12980 32824 12986
rect 32772 12922 32824 12928
rect 32312 12912 32364 12918
rect 32312 12854 32364 12860
rect 32220 12368 32272 12374
rect 32220 12310 32272 12316
rect 32036 12164 32088 12170
rect 32036 12106 32088 12112
rect 31852 12096 31904 12102
rect 31852 12038 31904 12044
rect 31484 11892 31536 11898
rect 31484 11834 31536 11840
rect 31760 11892 31812 11898
rect 31760 11834 31812 11840
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31024 10804 31076 10810
rect 31024 10746 31076 10752
rect 31036 7478 31064 10746
rect 31220 10742 31248 11698
rect 31208 10736 31260 10742
rect 31208 10678 31260 10684
rect 31116 10668 31168 10674
rect 31116 10610 31168 10616
rect 31128 9994 31156 10610
rect 31300 10600 31352 10606
rect 31404 10588 31432 11698
rect 31352 10560 31432 10588
rect 31300 10542 31352 10548
rect 31208 10532 31260 10538
rect 31208 10474 31260 10480
rect 31116 9988 31168 9994
rect 31116 9930 31168 9936
rect 31128 9178 31156 9930
rect 31116 9172 31168 9178
rect 31116 9114 31168 9120
rect 31024 7472 31076 7478
rect 31024 7414 31076 7420
rect 31220 4826 31248 10474
rect 31496 6662 31524 11834
rect 31864 11150 31892 12038
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31576 11076 31628 11082
rect 31576 11018 31628 11024
rect 31588 9994 31616 11018
rect 32324 10810 32352 12854
rect 32588 12844 32640 12850
rect 32508 12804 32588 12832
rect 32508 11354 32536 12804
rect 32588 12786 32640 12792
rect 32864 12844 32916 12850
rect 32864 12786 32916 12792
rect 32588 12640 32640 12646
rect 32588 12582 32640 12588
rect 32600 12238 32628 12582
rect 32588 12232 32640 12238
rect 32588 12174 32640 12180
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 32496 11348 32548 11354
rect 32496 11290 32548 11296
rect 32784 11218 32812 11698
rect 32876 11218 32904 12786
rect 32772 11212 32824 11218
rect 32772 11154 32824 11160
rect 32864 11212 32916 11218
rect 32864 11154 32916 11160
rect 32312 10804 32364 10810
rect 32312 10746 32364 10752
rect 32220 10668 32272 10674
rect 32220 10610 32272 10616
rect 32232 10266 32260 10610
rect 32220 10260 32272 10266
rect 32220 10202 32272 10208
rect 32324 10198 32352 10746
rect 32496 10668 32548 10674
rect 32496 10610 32548 10616
rect 32508 10266 32536 10610
rect 32876 10606 32904 11154
rect 32968 10674 32996 19774
rect 33060 18766 33088 24074
rect 33152 23322 33180 24142
rect 33232 23724 33284 23730
rect 33232 23666 33284 23672
rect 33140 23316 33192 23322
rect 33140 23258 33192 23264
rect 33244 23254 33272 23666
rect 33232 23248 33284 23254
rect 33232 23190 33284 23196
rect 33324 23112 33376 23118
rect 33324 23054 33376 23060
rect 33140 22704 33192 22710
rect 33140 22646 33192 22652
rect 33152 22506 33180 22646
rect 33232 22636 33284 22642
rect 33232 22578 33284 22584
rect 33140 22500 33192 22506
rect 33140 22442 33192 22448
rect 33244 22098 33272 22578
rect 33232 22092 33284 22098
rect 33232 22034 33284 22040
rect 33336 21894 33364 23054
rect 33324 21888 33376 21894
rect 33324 21830 33376 21836
rect 33324 19372 33376 19378
rect 33324 19314 33376 19320
rect 33336 18970 33364 19314
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 33048 18760 33100 18766
rect 33048 18702 33100 18708
rect 33060 18426 33088 18702
rect 33048 18420 33100 18426
rect 33048 18362 33100 18368
rect 33428 16017 33456 24942
rect 33600 24812 33652 24818
rect 33600 24754 33652 24760
rect 33612 24410 33640 24754
rect 33600 24404 33652 24410
rect 33600 24346 33652 24352
rect 33508 24132 33560 24138
rect 33508 24074 33560 24080
rect 33520 22710 33548 24074
rect 33704 23202 33732 28358
rect 33796 28082 33824 28426
rect 34072 28082 34100 29022
rect 34244 29028 34296 29034
rect 34244 28970 34296 28976
rect 34532 28694 34560 30670
rect 34612 29504 34664 29510
rect 34612 29446 34664 29452
rect 34624 28762 34652 29446
rect 34612 28756 34664 28762
rect 34612 28698 34664 28704
rect 34520 28688 34572 28694
rect 34520 28630 34572 28636
rect 34532 28082 34560 28630
rect 34716 28558 34744 37810
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35348 36576 35400 36582
rect 35348 36518 35400 36524
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35360 36174 35388 36518
rect 35348 36168 35400 36174
rect 35348 36110 35400 36116
rect 34796 35692 34848 35698
rect 34796 35634 34848 35640
rect 34808 34746 34836 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 34740 34848 34746
rect 34796 34682 34848 34688
rect 35360 34474 35388 36110
rect 35348 34468 35400 34474
rect 35348 34410 35400 34416
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35360 34202 35388 34410
rect 35348 34196 35400 34202
rect 35348 34138 35400 34144
rect 35452 34082 35480 38916
rect 36084 38888 36136 38894
rect 36084 38830 36136 38836
rect 58162 38856 58218 38865
rect 36096 38418 36124 38830
rect 58162 38791 58164 38800
rect 58216 38791 58218 38800
rect 58164 38762 58216 38768
rect 36084 38412 36136 38418
rect 36084 38354 36136 38360
rect 35532 37664 35584 37670
rect 35532 37606 35584 37612
rect 35360 34054 35480 34082
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 33046 35388 34054
rect 35348 33040 35400 33046
rect 35348 32982 35400 32988
rect 34796 32972 34848 32978
rect 34796 32914 34848 32920
rect 34808 29306 34836 32914
rect 35072 32836 35124 32842
rect 35072 32778 35124 32784
rect 35084 32502 35112 32778
rect 35072 32496 35124 32502
rect 35072 32438 35124 32444
rect 35348 32496 35400 32502
rect 35348 32438 35400 32444
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35360 31754 35388 32438
rect 35348 31748 35400 31754
rect 35348 31690 35400 31696
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30598 35388 31690
rect 35348 30592 35400 30598
rect 35348 30534 35400 30540
rect 35360 30190 35388 30534
rect 35348 30184 35400 30190
rect 35348 30126 35400 30132
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 34980 29164 35032 29170
rect 34980 29106 35032 29112
rect 34992 29050 35020 29106
rect 34808 29022 35020 29050
rect 34704 28552 34756 28558
rect 34704 28494 34756 28500
rect 34808 28370 34836 29022
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28558 35388 30126
rect 35440 29640 35492 29646
rect 35440 29582 35492 29588
rect 35452 29170 35480 29582
rect 35544 29510 35572 37606
rect 36096 36106 36124 38354
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 58164 37664 58216 37670
rect 58164 37606 58216 37612
rect 58176 37505 58204 37606
rect 58162 37496 58218 37505
rect 58162 37431 58218 37440
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 36636 36644 36688 36650
rect 36636 36586 36688 36592
rect 36648 36378 36676 36586
rect 36636 36372 36688 36378
rect 36636 36314 36688 36320
rect 58164 36168 58216 36174
rect 58162 36136 58164 36145
rect 58216 36136 58218 36145
rect 36084 36100 36136 36106
rect 36084 36042 36136 36048
rect 38568 36100 38620 36106
rect 58162 36071 58218 36080
rect 38568 36042 38620 36048
rect 36096 35766 36124 36042
rect 36084 35760 36136 35766
rect 36084 35702 36136 35708
rect 35900 33992 35952 33998
rect 35900 33934 35952 33940
rect 36084 33992 36136 33998
rect 36084 33934 36136 33940
rect 35912 33590 35940 33934
rect 35900 33584 35952 33590
rect 35900 33526 35952 33532
rect 35808 33040 35860 33046
rect 35808 32982 35860 32988
rect 35820 32774 35848 32982
rect 35912 32910 35940 33526
rect 35992 33516 36044 33522
rect 35992 33458 36044 33464
rect 36004 33114 36032 33458
rect 35992 33108 36044 33114
rect 35992 33050 36044 33056
rect 36096 32994 36124 33934
rect 36452 33924 36504 33930
rect 36452 33866 36504 33872
rect 36464 33454 36492 33866
rect 38200 33856 38252 33862
rect 38200 33798 38252 33804
rect 36452 33448 36504 33454
rect 36452 33390 36504 33396
rect 36004 32966 36124 32994
rect 35900 32904 35952 32910
rect 35900 32846 35952 32852
rect 35808 32768 35860 32774
rect 35808 32710 35860 32716
rect 35820 31822 35848 32710
rect 36004 32026 36032 32966
rect 36084 32904 36136 32910
rect 36084 32846 36136 32852
rect 36268 32904 36320 32910
rect 36268 32846 36320 32852
rect 36096 32570 36124 32846
rect 36084 32564 36136 32570
rect 36084 32506 36136 32512
rect 36280 32502 36308 32846
rect 36464 32842 36492 33390
rect 37280 33312 37332 33318
rect 37280 33254 37332 33260
rect 37292 32978 37320 33254
rect 37280 32972 37332 32978
rect 37280 32914 37332 32920
rect 38212 32910 38240 33798
rect 38580 33522 38608 36042
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 58164 35080 58216 35086
rect 58164 35022 58216 35028
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 58176 34785 58204 35022
rect 58162 34776 58218 34785
rect 58162 34711 58218 34720
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 38568 33516 38620 33522
rect 38568 33458 38620 33464
rect 38580 32978 38608 33458
rect 58162 33416 58218 33425
rect 58162 33351 58164 33360
rect 58216 33351 58218 33360
rect 58164 33322 58216 33328
rect 38568 32972 38620 32978
rect 38568 32914 38620 32920
rect 38200 32904 38252 32910
rect 38200 32846 38252 32852
rect 36452 32836 36504 32842
rect 36452 32778 36504 32784
rect 36268 32496 36320 32502
rect 36268 32438 36320 32444
rect 36084 32428 36136 32434
rect 36084 32370 36136 32376
rect 36096 32026 36124 32370
rect 35992 32020 36044 32026
rect 35992 31962 36044 31968
rect 36084 32020 36136 32026
rect 36084 31962 36136 31968
rect 35808 31816 35860 31822
rect 35808 31758 35860 31764
rect 36096 31414 36124 31962
rect 36084 31408 36136 31414
rect 36084 31350 36136 31356
rect 35900 30660 35952 30666
rect 35900 30602 35952 30608
rect 35912 30326 35940 30602
rect 35900 30320 35952 30326
rect 35900 30262 35952 30268
rect 36464 30258 36492 32778
rect 36544 32768 36596 32774
rect 36544 32710 36596 32716
rect 36556 31822 36584 32710
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 58164 32224 58216 32230
rect 58164 32166 58216 32172
rect 58176 32065 58204 32166
rect 58162 32056 58218 32065
rect 58162 31991 58218 32000
rect 36544 31816 36596 31822
rect 36544 31758 36596 31764
rect 38568 31816 38620 31822
rect 38568 31758 38620 31764
rect 38580 30734 38608 31758
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 38568 30728 38620 30734
rect 58164 30728 58216 30734
rect 38568 30670 38620 30676
rect 58162 30696 58164 30705
rect 58216 30696 58218 30705
rect 35992 30252 36044 30258
rect 35992 30194 36044 30200
rect 36452 30252 36504 30258
rect 36452 30194 36504 30200
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 35716 30048 35768 30054
rect 35716 29990 35768 29996
rect 35728 29646 35756 29990
rect 36004 29714 36032 30194
rect 35992 29708 36044 29714
rect 35992 29650 36044 29656
rect 35716 29640 35768 29646
rect 35900 29640 35952 29646
rect 35716 29582 35768 29588
rect 35820 29600 35900 29628
rect 35820 29510 35848 29600
rect 35900 29582 35952 29588
rect 35532 29504 35584 29510
rect 35532 29446 35584 29452
rect 35808 29504 35860 29510
rect 35808 29446 35860 29452
rect 36004 29238 36032 29650
rect 37476 29510 37504 30194
rect 38580 29646 38608 30670
rect 58162 30631 58218 30640
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 38568 29640 38620 29646
rect 38568 29582 38620 29588
rect 58164 29640 58216 29646
rect 58164 29582 58216 29588
rect 37464 29504 37516 29510
rect 37464 29446 37516 29452
rect 35992 29232 36044 29238
rect 35992 29174 36044 29180
rect 38580 29170 38608 29582
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 58176 29345 58204 29582
rect 58162 29336 58218 29345
rect 58162 29271 58218 29280
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 35624 29164 35676 29170
rect 35624 29106 35676 29112
rect 38568 29164 38620 29170
rect 38568 29106 38620 29112
rect 35440 29028 35492 29034
rect 35440 28970 35492 28976
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 34716 28342 34836 28370
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 34060 28076 34112 28082
rect 34060 28018 34112 28024
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 34532 27470 34560 28018
rect 34716 27470 34744 28342
rect 34796 27872 34848 27878
rect 34796 27814 34848 27820
rect 34808 27470 34836 27814
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35452 27470 35480 28970
rect 35636 28762 35664 29106
rect 35900 29028 35952 29034
rect 35900 28970 35952 28976
rect 35624 28756 35676 28762
rect 35624 28698 35676 28704
rect 35912 28558 35940 28970
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 37280 28076 37332 28082
rect 37280 28018 37332 28024
rect 37292 27674 37320 28018
rect 37280 27668 37332 27674
rect 37280 27610 37332 27616
rect 38580 27470 38608 29106
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 38660 28076 38712 28082
rect 38660 28018 38712 28024
rect 33968 27464 34020 27470
rect 33782 27432 33838 27441
rect 33968 27406 34020 27412
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34796 27464 34848 27470
rect 34796 27406 34848 27412
rect 35072 27464 35124 27470
rect 35072 27406 35124 27412
rect 35440 27464 35492 27470
rect 35440 27406 35492 27412
rect 38568 27464 38620 27470
rect 38568 27406 38620 27412
rect 33782 27367 33784 27376
rect 33836 27367 33838 27376
rect 33784 27338 33836 27344
rect 33980 27130 34008 27406
rect 35084 27130 35112 27406
rect 33968 27124 34020 27130
rect 33968 27066 34020 27072
rect 35072 27124 35124 27130
rect 35072 27066 35124 27072
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 38580 26450 38608 27406
rect 38568 26444 38620 26450
rect 38568 26386 38620 26392
rect 37280 26308 37332 26314
rect 37280 26250 37332 26256
rect 36636 26240 36688 26246
rect 36636 26182 36688 26188
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36648 25226 36676 26182
rect 37292 26042 37320 26250
rect 38016 26240 38068 26246
rect 38016 26182 38068 26188
rect 37280 26036 37332 26042
rect 37280 25978 37332 25984
rect 37188 25900 37240 25906
rect 37188 25842 37240 25848
rect 37832 25900 37884 25906
rect 37832 25842 37884 25848
rect 37924 25900 37976 25906
rect 37924 25842 37976 25848
rect 36728 25288 36780 25294
rect 36728 25230 36780 25236
rect 36636 25220 36688 25226
rect 36636 25162 36688 25168
rect 33876 24608 33928 24614
rect 33876 24550 33928 24556
rect 33612 23174 33732 23202
rect 33508 22704 33560 22710
rect 33508 22646 33560 22652
rect 33508 22500 33560 22506
rect 33508 22442 33560 22448
rect 33520 21894 33548 22442
rect 33612 22166 33640 23174
rect 33888 23118 33916 24550
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35716 23792 35768 23798
rect 35716 23734 35768 23740
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 33876 23112 33928 23118
rect 33876 23054 33928 23060
rect 33692 23044 33744 23050
rect 33692 22986 33744 22992
rect 33704 22778 33732 22986
rect 34704 22976 34756 22982
rect 34704 22918 34756 22924
rect 33692 22772 33744 22778
rect 33692 22714 33744 22720
rect 33600 22160 33652 22166
rect 33600 22102 33652 22108
rect 34716 22030 34744 22918
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 33508 21888 33560 21894
rect 33508 21830 33560 21836
rect 35624 21888 35676 21894
rect 35624 21830 35676 21836
rect 33520 21690 33548 21830
rect 33508 21684 33560 21690
rect 33508 21626 33560 21632
rect 35348 21480 35400 21486
rect 35348 21422 35400 21428
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34796 21072 34848 21078
rect 34796 21014 34848 21020
rect 34808 20058 34836 21014
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34796 20052 34848 20058
rect 34796 19994 34848 20000
rect 35360 19378 35388 21422
rect 35636 21010 35664 21830
rect 35624 21004 35676 21010
rect 35624 20946 35676 20952
rect 35728 19854 35756 23734
rect 35900 22092 35952 22098
rect 35900 22034 35952 22040
rect 35912 21078 35940 22034
rect 35992 21956 36044 21962
rect 35992 21898 36044 21904
rect 35900 21072 35952 21078
rect 35900 21014 35952 21020
rect 35912 20466 35940 21014
rect 36004 20942 36032 21898
rect 36452 21684 36504 21690
rect 36452 21626 36504 21632
rect 35992 20936 36044 20942
rect 35992 20878 36044 20884
rect 36004 20482 36032 20878
rect 36004 20466 36124 20482
rect 35900 20460 35952 20466
rect 35900 20402 35952 20408
rect 36004 20460 36136 20466
rect 36004 20454 36084 20460
rect 35716 19848 35768 19854
rect 35716 19790 35768 19796
rect 35348 19372 35400 19378
rect 35348 19314 35400 19320
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18834 35388 19314
rect 35912 18834 35940 20402
rect 36004 19378 36032 20454
rect 36084 20402 36136 20408
rect 36464 20330 36492 21626
rect 36544 21480 36596 21486
rect 36544 21422 36596 21428
rect 36452 20324 36504 20330
rect 36452 20266 36504 20272
rect 36360 19984 36412 19990
rect 36360 19926 36412 19932
rect 36268 19916 36320 19922
rect 36268 19858 36320 19864
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 35348 18828 35400 18834
rect 35348 18770 35400 18776
rect 35900 18828 35952 18834
rect 35900 18770 35952 18776
rect 35360 18426 35388 18770
rect 35348 18420 35400 18426
rect 35348 18362 35400 18368
rect 35912 18290 35940 18770
rect 36004 18358 36032 19314
rect 36280 19310 36308 19858
rect 36268 19304 36320 19310
rect 36268 19246 36320 19252
rect 36084 18692 36136 18698
rect 36084 18634 36136 18640
rect 35992 18352 36044 18358
rect 35992 18294 36044 18300
rect 33508 18284 33560 18290
rect 33508 18226 33560 18232
rect 35900 18284 35952 18290
rect 35900 18226 35952 18232
rect 33520 18086 33548 18226
rect 33508 18080 33560 18086
rect 33508 18022 33560 18028
rect 33414 16008 33470 16017
rect 33414 15943 33470 15952
rect 33232 15904 33284 15910
rect 33232 15846 33284 15852
rect 33244 15026 33272 15846
rect 33232 15020 33284 15026
rect 33232 14962 33284 14968
rect 33140 13864 33192 13870
rect 33140 13806 33192 13812
rect 33152 13394 33180 13806
rect 33140 13388 33192 13394
rect 33140 13330 33192 13336
rect 33520 13258 33548 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35348 17876 35400 17882
rect 35348 17818 35400 17824
rect 35360 17678 35388 17818
rect 36096 17678 36124 18634
rect 35348 17672 35400 17678
rect 35348 17614 35400 17620
rect 36084 17672 36136 17678
rect 36084 17614 36136 17620
rect 34980 17604 35032 17610
rect 34980 17546 35032 17552
rect 35256 17604 35308 17610
rect 35256 17546 35308 17552
rect 34992 17134 35020 17546
rect 35268 17338 35296 17546
rect 36096 17542 36124 17614
rect 36280 17610 36308 19246
rect 36372 18766 36400 19926
rect 36360 18760 36412 18766
rect 36360 18702 36412 18708
rect 36452 18284 36504 18290
rect 36452 18226 36504 18232
rect 36360 17672 36412 17678
rect 36360 17614 36412 17620
rect 36176 17604 36228 17610
rect 36176 17546 36228 17552
rect 36268 17604 36320 17610
rect 36268 17546 36320 17552
rect 35900 17536 35952 17542
rect 35900 17478 35952 17484
rect 36084 17536 36136 17542
rect 36084 17478 36136 17484
rect 35256 17332 35308 17338
rect 35256 17274 35308 17280
rect 35912 17202 35940 17478
rect 35900 17196 35952 17202
rect 35900 17138 35952 17144
rect 36096 17134 36124 17478
rect 33784 17128 33836 17134
rect 33784 17070 33836 17076
rect 34612 17128 34664 17134
rect 34612 17070 34664 17076
rect 34980 17128 35032 17134
rect 34980 17070 35032 17076
rect 36084 17128 36136 17134
rect 36084 17070 36136 17076
rect 33796 16726 33824 17070
rect 34060 16788 34112 16794
rect 34060 16730 34112 16736
rect 33784 16720 33836 16726
rect 33784 16662 33836 16668
rect 34072 15706 34100 16730
rect 34624 16114 34652 17070
rect 35532 16992 35584 16998
rect 35532 16934 35584 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34704 16652 34756 16658
rect 34704 16594 34756 16600
rect 34716 16538 34744 16594
rect 35544 16590 35572 16934
rect 35900 16788 35952 16794
rect 35900 16730 35952 16736
rect 34980 16584 35032 16590
rect 34716 16510 34836 16538
rect 34980 16526 35032 16532
rect 35532 16584 35584 16590
rect 35532 16526 35584 16532
rect 34704 16448 34756 16454
rect 34704 16390 34756 16396
rect 34612 16108 34664 16114
rect 34612 16050 34664 16056
rect 34520 16040 34572 16046
rect 34520 15982 34572 15988
rect 34060 15700 34112 15706
rect 34060 15642 34112 15648
rect 34072 15502 34100 15642
rect 34060 15496 34112 15502
rect 34060 15438 34112 15444
rect 34072 15162 34100 15438
rect 34060 15156 34112 15162
rect 34060 15098 34112 15104
rect 34072 14958 34100 15098
rect 34532 15026 34560 15982
rect 34612 15428 34664 15434
rect 34612 15370 34664 15376
rect 34520 15020 34572 15026
rect 34520 14962 34572 14968
rect 34060 14952 34112 14958
rect 34060 14894 34112 14900
rect 34532 14414 34560 14962
rect 34624 14618 34652 15370
rect 34716 14958 34744 16390
rect 34808 15502 34836 16510
rect 34992 16250 35020 16526
rect 34980 16244 35032 16250
rect 34980 16186 35032 16192
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34796 15496 34848 15502
rect 34796 15438 34848 15444
rect 34704 14952 34756 14958
rect 34704 14894 34756 14900
rect 34612 14612 34664 14618
rect 34612 14554 34664 14560
rect 34520 14408 34572 14414
rect 34520 14350 34572 14356
rect 33508 13252 33560 13258
rect 33508 13194 33560 13200
rect 34428 13252 34480 13258
rect 34428 13194 34480 13200
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 33060 11694 33088 12922
rect 34440 12442 34468 13194
rect 34428 12436 34480 12442
rect 34428 12378 34480 12384
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 32956 10668 33008 10674
rect 32956 10610 33008 10616
rect 32864 10600 32916 10606
rect 32864 10542 32916 10548
rect 34428 10532 34480 10538
rect 34428 10474 34480 10480
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 32496 10260 32548 10266
rect 32496 10202 32548 10208
rect 32312 10192 32364 10198
rect 32312 10134 32364 10140
rect 31576 9988 31628 9994
rect 31576 9930 31628 9936
rect 32128 9988 32180 9994
rect 32128 9930 32180 9936
rect 31588 9654 31616 9930
rect 31576 9648 31628 9654
rect 31576 9590 31628 9596
rect 32140 9382 32168 9930
rect 33244 9654 33272 10406
rect 33232 9648 33284 9654
rect 33232 9590 33284 9596
rect 32128 9376 32180 9382
rect 32128 9318 32180 9324
rect 32772 9376 32824 9382
rect 32772 9318 32824 9324
rect 32140 8566 32168 9318
rect 32128 8560 32180 8566
rect 32128 8502 32180 8508
rect 32784 7954 32812 9318
rect 34244 8288 34296 8294
rect 34244 8230 34296 8236
rect 32772 7948 32824 7954
rect 32772 7890 32824 7896
rect 32784 6798 32812 7890
rect 34256 7886 34284 8230
rect 34244 7880 34296 7886
rect 34244 7822 34296 7828
rect 33784 7744 33836 7750
rect 33784 7686 33836 7692
rect 32772 6792 32824 6798
rect 32772 6734 32824 6740
rect 31484 6656 31536 6662
rect 31484 6598 31536 6604
rect 31496 6390 31524 6598
rect 31484 6384 31536 6390
rect 31484 6326 31536 6332
rect 32784 5778 32812 6734
rect 33796 6458 33824 7686
rect 34440 7546 34468 10474
rect 34532 10282 34560 14350
rect 34716 14074 34744 14894
rect 34704 14068 34756 14074
rect 34704 14010 34756 14016
rect 34808 13954 34836 15438
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35440 14272 35492 14278
rect 35440 14214 35492 14220
rect 34624 13926 34836 13954
rect 34624 10441 34652 13926
rect 35452 13870 35480 14214
rect 35348 13864 35400 13870
rect 35348 13806 35400 13812
rect 35440 13864 35492 13870
rect 35440 13806 35492 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34704 13320 34756 13326
rect 34704 13262 34756 13268
rect 34716 12306 34744 13262
rect 34796 13252 34848 13258
rect 34796 13194 34848 13200
rect 34704 12300 34756 12306
rect 34704 12242 34756 12248
rect 34716 11286 34744 12242
rect 34808 12170 34836 13194
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35360 12434 35388 13806
rect 35268 12406 35388 12434
rect 35268 12238 35296 12406
rect 35452 12306 35480 13806
rect 35544 12374 35572 16526
rect 35912 16182 35940 16730
rect 35900 16176 35952 16182
rect 35900 16118 35952 16124
rect 35900 15156 35952 15162
rect 35900 15098 35952 15104
rect 35912 14074 35940 15098
rect 35900 14068 35952 14074
rect 35900 14010 35952 14016
rect 35912 13954 35940 14010
rect 36188 14006 36216 17546
rect 36280 17338 36308 17546
rect 36268 17332 36320 17338
rect 36268 17274 36320 17280
rect 36372 16794 36400 17614
rect 36360 16788 36412 16794
rect 36360 16730 36412 16736
rect 36360 16176 36412 16182
rect 36360 16118 36412 16124
rect 36268 14408 36320 14414
rect 36268 14350 36320 14356
rect 36176 14000 36228 14006
rect 35808 13932 35860 13938
rect 35912 13926 36124 13954
rect 36176 13942 36228 13948
rect 35808 13874 35860 13880
rect 35820 12850 35848 13874
rect 35808 12844 35860 12850
rect 35808 12786 35860 12792
rect 35624 12776 35676 12782
rect 35624 12718 35676 12724
rect 35532 12368 35584 12374
rect 35532 12310 35584 12316
rect 35440 12300 35492 12306
rect 35440 12242 35492 12248
rect 35636 12238 35664 12718
rect 35900 12436 35952 12442
rect 35900 12378 35952 12384
rect 35256 12232 35308 12238
rect 35256 12174 35308 12180
rect 35624 12232 35676 12238
rect 35624 12174 35676 12180
rect 34796 12164 34848 12170
rect 34796 12106 34848 12112
rect 34888 12164 34940 12170
rect 34888 12106 34940 12112
rect 34900 11762 34928 12106
rect 34888 11756 34940 11762
rect 34888 11698 34940 11704
rect 35348 11552 35400 11558
rect 35348 11494 35400 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34704 11280 34756 11286
rect 35360 11234 35388 11494
rect 34704 11222 34756 11228
rect 34716 10742 34744 11222
rect 35268 11206 35388 11234
rect 35268 11082 35296 11206
rect 35256 11076 35308 11082
rect 35256 11018 35308 11024
rect 35440 11008 35492 11014
rect 35440 10950 35492 10956
rect 34704 10736 34756 10742
rect 34704 10678 34756 10684
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34610 10432 34666 10441
rect 34610 10367 34666 10376
rect 34532 10254 34744 10282
rect 34808 10266 34836 10610
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34520 10192 34572 10198
rect 34520 10134 34572 10140
rect 34610 10160 34666 10169
rect 34532 8498 34560 10134
rect 34610 10095 34666 10104
rect 34624 9602 34652 10095
rect 34716 9722 34744 10254
rect 34796 10260 34848 10266
rect 34796 10202 34848 10208
rect 34980 10260 35032 10266
rect 34980 10202 35032 10208
rect 34992 10062 35020 10202
rect 35452 10130 35480 10950
rect 35440 10124 35492 10130
rect 35440 10066 35492 10072
rect 34980 10056 35032 10062
rect 35348 10056 35400 10062
rect 34980 9998 35032 10004
rect 35268 10016 35348 10044
rect 35268 9926 35296 10016
rect 35348 9998 35400 10004
rect 35256 9920 35308 9926
rect 35256 9862 35308 9868
rect 35348 9920 35400 9926
rect 35348 9862 35400 9868
rect 34704 9716 34756 9722
rect 34704 9658 34756 9664
rect 34624 9586 34744 9602
rect 34624 9580 34756 9586
rect 34624 9574 34704 9580
rect 34520 8492 34572 8498
rect 34520 8434 34572 8440
rect 34428 7540 34480 7546
rect 34428 7482 34480 7488
rect 34060 7472 34112 7478
rect 34060 7414 34112 7420
rect 34624 7426 34652 9574
rect 34704 9522 34756 9528
rect 34796 9580 34848 9586
rect 34796 9522 34848 9528
rect 34704 8492 34756 8498
rect 34704 8434 34756 8440
rect 34716 8090 34744 8434
rect 34704 8084 34756 8090
rect 34704 8026 34756 8032
rect 34808 8022 34836 9522
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34796 8016 34848 8022
rect 34796 7958 34848 7964
rect 34808 7886 34836 7958
rect 35360 7886 35388 9862
rect 35636 9518 35664 12174
rect 35912 11354 35940 12378
rect 36096 11762 36124 13926
rect 36188 13530 36216 13942
rect 36176 13524 36228 13530
rect 36176 13466 36228 13472
rect 36280 12850 36308 14350
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 36372 12442 36400 16118
rect 36360 12436 36412 12442
rect 36360 12378 36412 12384
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 35900 11348 35952 11354
rect 35900 11290 35952 11296
rect 35912 11150 35940 11290
rect 36360 11280 36412 11286
rect 36360 11222 36412 11228
rect 35900 11144 35952 11150
rect 35900 11086 35952 11092
rect 35900 11008 35952 11014
rect 35900 10950 35952 10956
rect 35912 10470 35940 10950
rect 35900 10464 35952 10470
rect 35900 10406 35952 10412
rect 35912 9654 35940 10406
rect 36268 9920 36320 9926
rect 36268 9862 36320 9868
rect 35900 9648 35952 9654
rect 35900 9590 35952 9596
rect 35992 9648 36044 9654
rect 35992 9590 36044 9596
rect 35440 9512 35492 9518
rect 35440 9454 35492 9460
rect 35624 9512 35676 9518
rect 35624 9454 35676 9460
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 35348 7880 35400 7886
rect 35348 7822 35400 7828
rect 34796 7540 34848 7546
rect 34796 7482 34848 7488
rect 34808 7426 34836 7482
rect 35452 7478 35480 9454
rect 35636 8498 35664 9454
rect 36004 8566 36032 9590
rect 36280 9586 36308 9862
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 36372 9042 36400 11222
rect 36464 9874 36492 18226
rect 36556 16182 36584 21422
rect 36648 20466 36676 25162
rect 36740 24274 36768 25230
rect 36728 24268 36780 24274
rect 36728 24210 36780 24216
rect 36740 23730 36768 24210
rect 36728 23724 36780 23730
rect 36728 23666 36780 23672
rect 36636 20460 36688 20466
rect 36636 20402 36688 20408
rect 36636 20324 36688 20330
rect 36636 20266 36688 20272
rect 36544 16176 36596 16182
rect 36544 16118 36596 16124
rect 36648 15910 36676 20266
rect 36740 17202 36768 23666
rect 37200 21894 37228 25842
rect 37556 25764 37608 25770
rect 37556 25706 37608 25712
rect 37464 25696 37516 25702
rect 37464 25638 37516 25644
rect 37476 25294 37504 25638
rect 37464 25288 37516 25294
rect 37464 25230 37516 25236
rect 37568 25158 37596 25706
rect 37844 25498 37872 25842
rect 37832 25492 37884 25498
rect 37832 25434 37884 25440
rect 37936 25294 37964 25842
rect 38028 25362 38056 26182
rect 38568 25900 38620 25906
rect 38568 25842 38620 25848
rect 38580 25498 38608 25842
rect 38568 25492 38620 25498
rect 38568 25434 38620 25440
rect 38016 25356 38068 25362
rect 38016 25298 38068 25304
rect 37740 25288 37792 25294
rect 37740 25230 37792 25236
rect 37924 25288 37976 25294
rect 37924 25230 37976 25236
rect 37556 25152 37608 25158
rect 37556 25094 37608 25100
rect 37372 24812 37424 24818
rect 37372 24754 37424 24760
rect 37384 23118 37412 24754
rect 37464 24744 37516 24750
rect 37464 24686 37516 24692
rect 37476 24070 37504 24686
rect 37568 24682 37596 25094
rect 37556 24676 37608 24682
rect 37556 24618 37608 24624
rect 37464 24064 37516 24070
rect 37464 24006 37516 24012
rect 37372 23112 37424 23118
rect 37372 23054 37424 23060
rect 37188 21888 37240 21894
rect 37188 21830 37240 21836
rect 37200 21554 37228 21830
rect 37188 21548 37240 21554
rect 37188 21490 37240 21496
rect 36912 21344 36964 21350
rect 36912 21286 36964 21292
rect 36924 20874 36952 21286
rect 36912 20868 36964 20874
rect 36912 20810 36964 20816
rect 36924 20534 36952 20810
rect 36912 20528 36964 20534
rect 36912 20470 36964 20476
rect 37188 18692 37240 18698
rect 37188 18634 37240 18640
rect 36820 18624 36872 18630
rect 36820 18566 36872 18572
rect 37004 18624 37056 18630
rect 37004 18566 37056 18572
rect 36832 17814 36860 18566
rect 36820 17808 36872 17814
rect 36820 17750 36872 17756
rect 36912 17536 36964 17542
rect 36912 17478 36964 17484
rect 36728 17196 36780 17202
rect 36728 17138 36780 17144
rect 36820 17128 36872 17134
rect 36820 17070 36872 17076
rect 36832 16114 36860 17070
rect 36924 16250 36952 17478
rect 36912 16244 36964 16250
rect 36912 16186 36964 16192
rect 36820 16108 36872 16114
rect 36820 16050 36872 16056
rect 36636 15904 36688 15910
rect 36636 15846 36688 15852
rect 36832 15502 36860 16050
rect 36912 15904 36964 15910
rect 36912 15846 36964 15852
rect 36820 15496 36872 15502
rect 36820 15438 36872 15444
rect 36832 14482 36860 15438
rect 36820 14476 36872 14482
rect 36820 14418 36872 14424
rect 36924 13734 36952 15846
rect 36912 13728 36964 13734
rect 36912 13670 36964 13676
rect 36544 13388 36596 13394
rect 36544 13330 36596 13336
rect 36556 12434 36584 13330
rect 36820 12844 36872 12850
rect 36820 12786 36872 12792
rect 36556 12406 36676 12434
rect 36544 9920 36596 9926
rect 36464 9868 36544 9874
rect 36464 9862 36596 9868
rect 36464 9846 36584 9862
rect 36648 9722 36676 12406
rect 36832 10062 36860 12786
rect 37016 10606 37044 18566
rect 37200 18358 37228 18634
rect 37188 18352 37240 18358
rect 37188 18294 37240 18300
rect 37096 18148 37148 18154
rect 37096 18090 37148 18096
rect 37108 16454 37136 18090
rect 37280 17672 37332 17678
rect 37200 17620 37280 17626
rect 37200 17614 37332 17620
rect 37200 17598 37320 17614
rect 37200 17338 37228 17598
rect 37188 17332 37240 17338
rect 37188 17274 37240 17280
rect 37096 16448 37148 16454
rect 37096 16390 37148 16396
rect 37108 15366 37136 16390
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 37200 15502 37228 16050
rect 37188 15496 37240 15502
rect 37188 15438 37240 15444
rect 37096 15360 37148 15366
rect 37096 15302 37148 15308
rect 37108 14958 37136 15302
rect 37200 15162 37228 15438
rect 37280 15428 37332 15434
rect 37280 15370 37332 15376
rect 37292 15162 37320 15370
rect 37188 15156 37240 15162
rect 37188 15098 37240 15104
rect 37280 15156 37332 15162
rect 37280 15098 37332 15104
rect 37096 14952 37148 14958
rect 37096 14894 37148 14900
rect 37108 14414 37136 14894
rect 37096 14408 37148 14414
rect 37096 14350 37148 14356
rect 37096 14272 37148 14278
rect 37096 14214 37148 14220
rect 37108 13394 37136 14214
rect 37384 14074 37412 23054
rect 37568 23050 37596 24618
rect 37648 23520 37700 23526
rect 37648 23462 37700 23468
rect 37660 23118 37688 23462
rect 37648 23112 37700 23118
rect 37648 23054 37700 23060
rect 37556 23044 37608 23050
rect 37556 22986 37608 22992
rect 37568 18154 37596 22986
rect 37752 22098 37780 25230
rect 37936 24818 37964 25230
rect 37924 24812 37976 24818
rect 37924 24754 37976 24760
rect 38672 24410 38700 28018
rect 58162 27976 58218 27985
rect 58162 27911 58164 27920
rect 58216 27911 58218 27920
rect 58164 27882 58216 27888
rect 40224 27872 40276 27878
rect 40224 27814 40276 27820
rect 40236 27470 40264 27814
rect 40224 27464 40276 27470
rect 40224 27406 40276 27412
rect 38936 26376 38988 26382
rect 38936 26318 38988 26324
rect 38752 25968 38804 25974
rect 38752 25910 38804 25916
rect 38764 24682 38792 25910
rect 38948 25702 38976 26318
rect 39028 26308 39080 26314
rect 39028 26250 39080 26256
rect 38936 25696 38988 25702
rect 38936 25638 38988 25644
rect 38844 24880 38896 24886
rect 38844 24822 38896 24828
rect 38752 24676 38804 24682
rect 38752 24618 38804 24624
rect 38660 24404 38712 24410
rect 38660 24346 38712 24352
rect 38672 24206 38700 24346
rect 38660 24200 38712 24206
rect 38660 24142 38712 24148
rect 37924 24064 37976 24070
rect 37924 24006 37976 24012
rect 37936 23662 37964 24006
rect 38200 23724 38252 23730
rect 38200 23666 38252 23672
rect 37924 23656 37976 23662
rect 37924 23598 37976 23604
rect 37936 23186 37964 23598
rect 38212 23322 38240 23666
rect 38200 23316 38252 23322
rect 38200 23258 38252 23264
rect 37924 23180 37976 23186
rect 37924 23122 37976 23128
rect 37936 22642 37964 23122
rect 37924 22636 37976 22642
rect 37924 22578 37976 22584
rect 38660 22432 38712 22438
rect 38712 22392 38792 22420
rect 38660 22374 38712 22380
rect 37740 22092 37792 22098
rect 37740 22034 37792 22040
rect 38764 21962 38792 22392
rect 38856 22030 38884 24822
rect 38844 22024 38896 22030
rect 38844 21966 38896 21972
rect 38752 21956 38804 21962
rect 38752 21898 38804 21904
rect 38660 21888 38712 21894
rect 38660 21830 38712 21836
rect 38672 21622 38700 21830
rect 38660 21616 38712 21622
rect 38660 21558 38712 21564
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 37752 21146 37780 21490
rect 37740 21140 37792 21146
rect 37740 21082 37792 21088
rect 38948 20942 38976 25638
rect 39040 24818 39068 26250
rect 40236 25906 40264 27406
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 58164 26784 58216 26790
rect 58164 26726 58216 26732
rect 58176 26625 58204 26726
rect 58162 26616 58218 26625
rect 58162 26551 58218 26560
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 40224 25900 40276 25906
rect 40224 25842 40276 25848
rect 39856 25696 39908 25702
rect 39856 25638 39908 25644
rect 39868 24886 39896 25638
rect 58164 25288 58216 25294
rect 58162 25256 58164 25265
rect 58216 25256 58218 25265
rect 58162 25191 58218 25200
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 39856 24880 39908 24886
rect 39856 24822 39908 24828
rect 39028 24812 39080 24818
rect 39028 24754 39080 24760
rect 39040 24274 39068 24754
rect 40132 24608 40184 24614
rect 40132 24550 40184 24556
rect 39028 24268 39080 24274
rect 39028 24210 39080 24216
rect 39672 23112 39724 23118
rect 39672 23054 39724 23060
rect 39120 22160 39172 22166
rect 39120 22102 39172 22108
rect 39132 21690 39160 22102
rect 39120 21684 39172 21690
rect 39120 21626 39172 21632
rect 38936 20936 38988 20942
rect 38936 20878 38988 20884
rect 39684 20058 39712 23054
rect 39856 22636 39908 22642
rect 39856 22578 39908 22584
rect 39868 22234 39896 22578
rect 40144 22506 40172 24550
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 58176 23905 58204 24142
rect 58162 23896 58218 23905
rect 58162 23831 58218 23840
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 58162 22536 58218 22545
rect 40132 22500 40184 22506
rect 58162 22471 58164 22480
rect 40132 22442 40184 22448
rect 58216 22471 58218 22480
rect 58164 22442 58216 22448
rect 39856 22228 39908 22234
rect 39856 22170 39908 22176
rect 40144 22030 40172 22442
rect 40224 22432 40276 22438
rect 40224 22374 40276 22380
rect 39856 22024 39908 22030
rect 39856 21966 39908 21972
rect 40132 22024 40184 22030
rect 40132 21966 40184 21972
rect 39868 21842 39896 21966
rect 39868 21814 40080 21842
rect 39764 21616 39816 21622
rect 39764 21558 39816 21564
rect 39776 20874 39804 21558
rect 40052 21554 40080 21814
rect 40040 21548 40092 21554
rect 40040 21490 40092 21496
rect 40040 21344 40092 21350
rect 40040 21286 40092 21292
rect 40132 21344 40184 21350
rect 40132 21286 40184 21292
rect 39764 20868 39816 20874
rect 39764 20810 39816 20816
rect 39672 20052 39724 20058
rect 39672 19994 39724 20000
rect 38660 19712 38712 19718
rect 38660 19654 38712 19660
rect 38672 19514 38700 19654
rect 38660 19508 38712 19514
rect 38660 19450 38712 19456
rect 38672 18766 38700 19450
rect 37648 18760 37700 18766
rect 37648 18702 37700 18708
rect 38660 18760 38712 18766
rect 38660 18702 38712 18708
rect 37556 18148 37608 18154
rect 37556 18090 37608 18096
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37476 15434 37504 17614
rect 37568 15910 37596 18090
rect 37556 15904 37608 15910
rect 37556 15846 37608 15852
rect 37464 15428 37516 15434
rect 37464 15370 37516 15376
rect 37556 15360 37608 15366
rect 37556 15302 37608 15308
rect 37568 15026 37596 15302
rect 37556 15020 37608 15026
rect 37556 14962 37608 14968
rect 37372 14068 37424 14074
rect 37372 14010 37424 14016
rect 37660 13410 37688 18702
rect 39776 18698 39804 20810
rect 39856 19712 39908 19718
rect 39856 19654 39908 19660
rect 39868 19446 39896 19654
rect 39856 19440 39908 19446
rect 39856 19382 39908 19388
rect 40052 19378 40080 21286
rect 40144 21010 40172 21286
rect 40132 21004 40184 21010
rect 40132 20946 40184 20952
rect 40236 20942 40264 22374
rect 40316 22024 40368 22030
rect 40316 21966 40368 21972
rect 40500 22024 40552 22030
rect 40552 21972 40632 21978
rect 40500 21966 40632 21972
rect 40328 21842 40356 21966
rect 40512 21950 40632 21966
rect 40328 21814 40540 21842
rect 40408 21548 40460 21554
rect 40408 21490 40460 21496
rect 40224 20936 40276 20942
rect 40224 20878 40276 20884
rect 40420 19378 40448 21490
rect 40512 21146 40540 21814
rect 40604 21554 40632 21950
rect 40684 21956 40736 21962
rect 40684 21898 40736 21904
rect 40960 21956 41012 21962
rect 40960 21898 41012 21904
rect 41144 21956 41196 21962
rect 41144 21898 41196 21904
rect 40696 21690 40724 21898
rect 40684 21684 40736 21690
rect 40684 21626 40736 21632
rect 40592 21548 40644 21554
rect 40592 21490 40644 21496
rect 40500 21140 40552 21146
rect 40500 21082 40552 21088
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40040 19372 40092 19378
rect 40040 19314 40092 19320
rect 40408 19372 40460 19378
rect 40408 19314 40460 19320
rect 39764 18692 39816 18698
rect 39764 18634 39816 18640
rect 38016 18420 38068 18426
rect 38016 18362 38068 18368
rect 37924 17740 37976 17746
rect 37924 17682 37976 17688
rect 37832 17536 37884 17542
rect 37832 17478 37884 17484
rect 37740 16992 37792 16998
rect 37740 16934 37792 16940
rect 37752 16250 37780 16934
rect 37740 16244 37792 16250
rect 37740 16186 37792 16192
rect 37844 15502 37872 17478
rect 37936 16726 37964 17682
rect 37924 16720 37976 16726
rect 37924 16662 37976 16668
rect 37832 15496 37884 15502
rect 37832 15438 37884 15444
rect 37844 14090 37872 15438
rect 37844 14074 37964 14090
rect 37740 14068 37792 14074
rect 37844 14068 37976 14074
rect 37844 14062 37924 14068
rect 37740 14010 37792 14016
rect 37924 14010 37976 14016
rect 37096 13388 37148 13394
rect 37096 13330 37148 13336
rect 37568 13382 37688 13410
rect 37096 13184 37148 13190
rect 37096 13126 37148 13132
rect 37108 12918 37136 13126
rect 37096 12912 37148 12918
rect 37096 12854 37148 12860
rect 37568 12850 37596 13382
rect 37752 13326 37780 14010
rect 37648 13320 37700 13326
rect 37648 13262 37700 13268
rect 37740 13320 37792 13326
rect 37740 13262 37792 13268
rect 37660 12986 37688 13262
rect 37648 12980 37700 12986
rect 37648 12922 37700 12928
rect 37556 12844 37608 12850
rect 37556 12786 37608 12792
rect 37188 12436 37240 12442
rect 37188 12378 37240 12384
rect 37200 11150 37228 12378
rect 37740 11688 37792 11694
rect 37740 11630 37792 11636
rect 37280 11552 37332 11558
rect 37280 11494 37332 11500
rect 37188 11144 37240 11150
rect 37188 11086 37240 11092
rect 37004 10600 37056 10606
rect 37004 10542 37056 10548
rect 36820 10056 36872 10062
rect 36820 9998 36872 10004
rect 36636 9716 36688 9722
rect 36636 9658 36688 9664
rect 37200 9586 37228 11086
rect 37292 10674 37320 11494
rect 37648 11076 37700 11082
rect 37648 11018 37700 11024
rect 37660 10810 37688 11018
rect 37648 10804 37700 10810
rect 37648 10746 37700 10752
rect 37280 10668 37332 10674
rect 37280 10610 37332 10616
rect 37292 10062 37320 10610
rect 37752 10198 37780 11630
rect 37740 10192 37792 10198
rect 37740 10134 37792 10140
rect 37280 10056 37332 10062
rect 37280 9998 37332 10004
rect 37280 9920 37332 9926
rect 37280 9862 37332 9868
rect 37464 9920 37516 9926
rect 37464 9862 37516 9868
rect 37292 9722 37320 9862
rect 37280 9716 37332 9722
rect 37280 9658 37332 9664
rect 37188 9580 37240 9586
rect 37188 9522 37240 9528
rect 36636 9376 36688 9382
rect 36636 9318 36688 9324
rect 36360 9036 36412 9042
rect 36360 8978 36412 8984
rect 36648 8974 36676 9318
rect 36636 8968 36688 8974
rect 36636 8910 36688 8916
rect 35992 8560 36044 8566
rect 35992 8502 36044 8508
rect 35624 8492 35676 8498
rect 35624 8434 35676 8440
rect 35532 7880 35584 7886
rect 35532 7822 35584 7828
rect 34072 6866 34100 7414
rect 34624 7410 34836 7426
rect 35440 7472 35492 7478
rect 35440 7414 35492 7420
rect 34624 7404 34848 7410
rect 34624 7398 34796 7404
rect 34796 7346 34848 7352
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34060 6860 34112 6866
rect 34060 6802 34112 6808
rect 33784 6452 33836 6458
rect 33784 6394 33836 6400
rect 34796 6316 34848 6322
rect 34796 6258 34848 6264
rect 34336 6112 34388 6118
rect 34336 6054 34388 6060
rect 32772 5772 32824 5778
rect 32772 5714 32824 5720
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 30656 4616 30708 4622
rect 30656 4558 30708 4564
rect 30932 4616 30984 4622
rect 30932 4558 30984 4564
rect 31576 4616 31628 4622
rect 31576 4558 31628 4564
rect 31588 4282 31616 4558
rect 31576 4276 31628 4282
rect 31576 4218 31628 4224
rect 30564 4208 30616 4214
rect 30564 4150 30616 4156
rect 32784 4146 32812 5714
rect 34348 4146 34376 6054
rect 34808 5914 34836 6258
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5908 34848 5914
rect 34796 5850 34848 5856
rect 35360 5710 35388 7346
rect 35348 5704 35400 5710
rect 35348 5646 35400 5652
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 30196 4140 30248 4146
rect 30196 4082 30248 4088
rect 32772 4140 32824 4146
rect 32772 4082 32824 4088
rect 34336 4140 34388 4146
rect 34336 4082 34388 4088
rect 35360 4010 35388 5646
rect 35544 5642 35572 7822
rect 35636 6322 35664 8434
rect 35808 7540 35860 7546
rect 36004 7528 36032 8502
rect 37200 7886 37228 9522
rect 37292 9518 37320 9658
rect 37280 9512 37332 9518
rect 37280 9454 37332 9460
rect 37476 9450 37504 9862
rect 37752 9589 37780 10134
rect 38028 10130 38056 18362
rect 39776 18358 39804 18634
rect 39764 18352 39816 18358
rect 39764 18294 39816 18300
rect 39028 18148 39080 18154
rect 39028 18090 39080 18096
rect 38752 18080 38804 18086
rect 38752 18022 38804 18028
rect 38764 17882 38792 18022
rect 38752 17876 38804 17882
rect 38752 17818 38804 17824
rect 38844 17672 38896 17678
rect 38844 17614 38896 17620
rect 38568 17604 38620 17610
rect 38568 17546 38620 17552
rect 38580 17202 38608 17546
rect 38568 17196 38620 17202
rect 38568 17138 38620 17144
rect 38200 17128 38252 17134
rect 38200 17070 38252 17076
rect 38212 14414 38240 17070
rect 38660 16516 38712 16522
rect 38660 16458 38712 16464
rect 38672 16046 38700 16458
rect 38856 16250 38884 17614
rect 39040 17338 39068 18090
rect 39212 17536 39264 17542
rect 39212 17478 39264 17484
rect 39028 17332 39080 17338
rect 39028 17274 39080 17280
rect 38844 16244 38896 16250
rect 38844 16186 38896 16192
rect 39028 16244 39080 16250
rect 39028 16186 39080 16192
rect 38660 16040 38712 16046
rect 38660 15982 38712 15988
rect 38384 15360 38436 15366
rect 38384 15302 38436 15308
rect 38200 14408 38252 14414
rect 38200 14350 38252 14356
rect 38212 13326 38240 14350
rect 38292 14340 38344 14346
rect 38292 14282 38344 14288
rect 38304 13870 38332 14282
rect 38292 13864 38344 13870
rect 38292 13806 38344 13812
rect 38200 13320 38252 13326
rect 38200 13262 38252 13268
rect 38304 13258 38332 13806
rect 38396 13326 38424 15302
rect 38568 15020 38620 15026
rect 38568 14962 38620 14968
rect 38580 13326 38608 14962
rect 39040 14890 39068 16186
rect 39224 16114 39252 17478
rect 39776 16998 39804 18294
rect 40052 18290 40080 19314
rect 39856 18284 39908 18290
rect 39856 18226 39908 18232
rect 40040 18284 40092 18290
rect 40040 18226 40092 18232
rect 39868 17882 39896 18226
rect 39856 17876 39908 17882
rect 39856 17818 39908 17824
rect 40052 16998 40080 18226
rect 40420 18170 40448 19314
rect 40512 18970 40540 19450
rect 40696 19242 40724 21626
rect 40972 21622 41000 21898
rect 40960 21616 41012 21622
rect 40960 21558 41012 21564
rect 41156 21350 41184 21898
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 41144 21344 41196 21350
rect 41144 21286 41196 21292
rect 58164 21344 58216 21350
rect 58164 21286 58216 21292
rect 58176 21185 58204 21286
rect 58162 21176 58218 21185
rect 58162 21111 58218 21120
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 40868 20052 40920 20058
rect 40868 19994 40920 20000
rect 40880 19378 40908 19994
rect 58164 19848 58216 19854
rect 58162 19816 58164 19825
rect 58216 19816 58218 19825
rect 58162 19751 58218 19760
rect 41052 19712 41104 19718
rect 41052 19654 41104 19660
rect 41064 19514 41092 19654
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 41052 19508 41104 19514
rect 41052 19450 41104 19456
rect 40868 19372 40920 19378
rect 40868 19314 40920 19320
rect 40684 19236 40736 19242
rect 40684 19178 40736 19184
rect 40500 18964 40552 18970
rect 40500 18906 40552 18912
rect 40420 18142 40540 18170
rect 40512 17678 40540 18142
rect 40592 18080 40644 18086
rect 40592 18022 40644 18028
rect 40500 17672 40552 17678
rect 40500 17614 40552 17620
rect 40512 17134 40540 17614
rect 40604 17610 40632 18022
rect 40592 17604 40644 17610
rect 40592 17546 40644 17552
rect 40696 17542 40724 19178
rect 58164 18760 58216 18766
rect 58164 18702 58216 18708
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 58176 18465 58204 18702
rect 58162 18456 58218 18465
rect 58162 18391 58218 18400
rect 40684 17536 40736 17542
rect 40684 17478 40736 17484
rect 40500 17128 40552 17134
rect 40500 17070 40552 17076
rect 39764 16992 39816 16998
rect 39764 16934 39816 16940
rect 40040 16992 40092 16998
rect 40040 16934 40092 16940
rect 40052 16658 40080 16934
rect 40040 16652 40092 16658
rect 40040 16594 40092 16600
rect 39212 16108 39264 16114
rect 39212 16050 39264 16056
rect 40052 15026 40080 16594
rect 40040 15020 40092 15026
rect 40040 14962 40092 14968
rect 39028 14884 39080 14890
rect 39028 14826 39080 14832
rect 38844 13932 38896 13938
rect 38844 13874 38896 13880
rect 38856 13530 38884 13874
rect 38844 13524 38896 13530
rect 38844 13466 38896 13472
rect 39040 13462 39068 14826
rect 40052 13938 40080 14962
rect 40224 14476 40276 14482
rect 40224 14418 40276 14424
rect 40236 14006 40264 14418
rect 40696 14414 40724 17478
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 58162 17096 58218 17105
rect 58162 17031 58164 17040
rect 58216 17031 58218 17040
rect 58164 17002 58216 17008
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 58164 15904 58216 15910
rect 58164 15846 58216 15852
rect 58176 15745 58204 15846
rect 58162 15736 58218 15745
rect 58162 15671 58218 15680
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 40684 14408 40736 14414
rect 58164 14408 58216 14414
rect 40684 14350 40736 14356
rect 58162 14376 58164 14385
rect 58216 14376 58218 14385
rect 58162 14311 58218 14320
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 40224 14000 40276 14006
rect 40224 13942 40276 13948
rect 40040 13932 40092 13938
rect 40040 13874 40092 13880
rect 39028 13456 39080 13462
rect 39028 13398 39080 13404
rect 38384 13320 38436 13326
rect 38384 13262 38436 13268
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 38292 13252 38344 13258
rect 38292 13194 38344 13200
rect 38304 11762 38332 13194
rect 38580 12102 38608 13262
rect 39120 13184 39172 13190
rect 39120 13126 39172 13132
rect 38568 12096 38620 12102
rect 38568 12038 38620 12044
rect 38292 11756 38344 11762
rect 38292 11698 38344 11704
rect 38936 11688 38988 11694
rect 38936 11630 38988 11636
rect 38568 11280 38620 11286
rect 38568 11222 38620 11228
rect 38580 10742 38608 11222
rect 38948 11150 38976 11630
rect 39132 11558 39160 13126
rect 40052 12850 40080 13874
rect 40236 13326 40264 13942
rect 40224 13320 40276 13326
rect 40224 13262 40276 13268
rect 58164 13320 58216 13326
rect 58164 13262 58216 13268
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 58176 13025 58204 13262
rect 58162 13016 58218 13025
rect 58162 12951 58218 12960
rect 40040 12844 40092 12850
rect 40040 12786 40092 12792
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 58162 11656 58218 11665
rect 58162 11591 58164 11600
rect 58216 11591 58218 11600
rect 58164 11562 58216 11568
rect 39120 11552 39172 11558
rect 39120 11494 39172 11500
rect 39132 11150 39160 11494
rect 38936 11144 38988 11150
rect 38936 11086 38988 11092
rect 39120 11144 39172 11150
rect 39120 11086 39172 11092
rect 39304 11008 39356 11014
rect 39304 10950 39356 10956
rect 38568 10736 38620 10742
rect 38568 10678 38620 10684
rect 38016 10124 38068 10130
rect 38016 10066 38068 10072
rect 37727 9583 37780 9589
rect 37779 9531 37780 9583
rect 37727 9525 37780 9531
rect 37464 9444 37516 9450
rect 37464 9386 37516 9392
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 37188 7880 37240 7886
rect 37188 7822 37240 7828
rect 37200 7562 37228 7822
rect 35808 7482 35860 7488
rect 35912 7500 36032 7528
rect 37108 7534 37228 7562
rect 37384 7546 37412 7958
rect 37752 7954 37780 9525
rect 38028 9178 38056 10066
rect 38384 9988 38436 9994
rect 38384 9930 38436 9936
rect 38016 9172 38068 9178
rect 38016 9114 38068 9120
rect 37740 7948 37792 7954
rect 37740 7890 37792 7896
rect 37372 7540 37424 7546
rect 35820 7410 35848 7482
rect 35808 7404 35860 7410
rect 35808 7346 35860 7352
rect 35912 6458 35940 7500
rect 36726 7440 36782 7449
rect 35992 7404 36044 7410
rect 35992 7346 36044 7352
rect 36084 7404 36136 7410
rect 37108 7410 37136 7534
rect 37372 7482 37424 7488
rect 37188 7472 37240 7478
rect 37188 7414 37240 7420
rect 36726 7375 36728 7384
rect 36084 7346 36136 7352
rect 36780 7375 36782 7384
rect 37096 7404 37148 7410
rect 36728 7346 36780 7352
rect 37096 7346 37148 7352
rect 35900 6452 35952 6458
rect 35900 6394 35952 6400
rect 35624 6316 35676 6322
rect 35624 6258 35676 6264
rect 35900 6316 35952 6322
rect 35900 6258 35952 6264
rect 35912 5914 35940 6258
rect 35900 5908 35952 5914
rect 35900 5850 35952 5856
rect 36004 5710 36032 7346
rect 36096 7002 36124 7346
rect 36084 6996 36136 7002
rect 36084 6938 36136 6944
rect 36096 6322 36124 6938
rect 37200 6662 37228 7414
rect 37464 7404 37516 7410
rect 37464 7346 37516 7352
rect 37280 6724 37332 6730
rect 37280 6666 37332 6672
rect 37188 6656 37240 6662
rect 37188 6598 37240 6604
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 35992 5704 36044 5710
rect 35992 5646 36044 5652
rect 35532 5636 35584 5642
rect 35532 5578 35584 5584
rect 36004 4826 36032 5646
rect 36096 5370 36124 6258
rect 37004 6112 37056 6118
rect 37004 6054 37056 6060
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 35992 4820 36044 4826
rect 35992 4762 36044 4768
rect 37016 4622 37044 6054
rect 37200 5710 37228 6598
rect 37292 6322 37320 6666
rect 37280 6316 37332 6322
rect 37280 6258 37332 6264
rect 37188 5704 37240 5710
rect 37188 5646 37240 5652
rect 37292 4690 37320 6258
rect 37476 5914 37504 7346
rect 37752 7274 37780 7890
rect 37832 7744 37884 7750
rect 37832 7686 37884 7692
rect 37740 7268 37792 7274
rect 37740 7210 37792 7216
rect 37844 6390 37872 7686
rect 37922 7440 37978 7449
rect 38396 7410 38424 9930
rect 38580 9586 38608 10678
rect 39316 10674 39344 10950
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 39304 10668 39356 10674
rect 39304 10610 39356 10616
rect 58164 10464 58216 10470
rect 58164 10406 58216 10412
rect 58176 10305 58204 10406
rect 58162 10296 58218 10305
rect 58162 10231 58218 10240
rect 39948 9920 40000 9926
rect 39948 9862 40000 9868
rect 39960 9722 39988 9862
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 39948 9716 40000 9722
rect 39948 9658 40000 9664
rect 38568 9580 38620 9586
rect 38568 9522 38620 9528
rect 58164 8968 58216 8974
rect 58162 8936 58164 8945
rect 58216 8936 58218 8945
rect 58162 8871 58218 8880
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 58164 7880 58216 7886
rect 58164 7822 58216 7828
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 58176 7585 58204 7822
rect 58162 7576 58218 7585
rect 58162 7511 58218 7520
rect 37922 7375 37924 7384
rect 37976 7375 37978 7384
rect 38384 7404 38436 7410
rect 37924 7346 37976 7352
rect 38384 7346 38436 7352
rect 38016 7200 38068 7206
rect 38016 7142 38068 7148
rect 38028 6798 38056 7142
rect 38016 6792 38068 6798
rect 38016 6734 38068 6740
rect 37832 6384 37884 6390
rect 37832 6326 37884 6332
rect 37464 5908 37516 5914
rect 37464 5850 37516 5856
rect 38396 5642 38424 7346
rect 39120 7336 39172 7342
rect 39120 7278 39172 7284
rect 39132 6458 39160 7278
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 39120 6452 39172 6458
rect 39120 6394 39172 6400
rect 58162 6216 58218 6225
rect 58162 6151 58164 6160
rect 58216 6151 58218 6160
rect 58164 6122 58216 6128
rect 38384 5636 38436 5642
rect 38384 5578 38436 5584
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 53748 5160 53800 5166
rect 53748 5102 53800 5108
rect 53656 5024 53708 5030
rect 53656 4966 53708 4972
rect 52184 4752 52236 4758
rect 52184 4694 52236 4700
rect 37280 4684 37332 4690
rect 37280 4626 37332 4632
rect 37004 4616 37056 4622
rect 37004 4558 37056 4564
rect 52092 4616 52144 4622
rect 52092 4558 52144 4564
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 51816 4072 51868 4078
rect 51816 4014 51868 4020
rect 35348 4004 35400 4010
rect 35348 3946 35400 3952
rect 29460 3936 29512 3942
rect 29460 3878 29512 3884
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 51356 3936 51408 3942
rect 51356 3878 51408 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 46296 3664 46348 3670
rect 46296 3606 46348 3612
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 44364 3528 44416 3534
rect 44364 3470 44416 3476
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 32772 2984 32824 2990
rect 28998 2952 29054 2961
rect 32772 2926 32824 2932
rect 28998 2887 29054 2896
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 28920 800 28948 2382
rect 29196 800 29224 2790
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 29472 800 29500 2382
rect 29748 800 29776 2790
rect 30024 800 30052 2790
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30300 800 30328 2382
rect 30576 800 30604 2790
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 30852 800 30880 2382
rect 31128 800 31156 2382
rect 31404 800 31432 2382
rect 31680 800 31708 2790
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 31956 800 31984 2450
rect 32232 800 32260 2790
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32508 800 32536 2382
rect 32784 800 32812 2926
rect 33876 2916 33928 2922
rect 33876 2858 33928 2864
rect 33324 2848 33376 2854
rect 33324 2790 33376 2796
rect 33048 2508 33100 2514
rect 33048 2450 33100 2456
rect 33060 800 33088 2450
rect 33336 800 33364 2790
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33612 800 33640 2382
rect 33888 800 33916 2858
rect 34428 2848 34480 2854
rect 34428 2790 34480 2796
rect 34152 2576 34204 2582
rect 34152 2518 34204 2524
rect 34164 800 34192 2518
rect 34440 800 34468 2790
rect 34716 800 34744 3470
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 1850 35388 3470
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 34992 1822 35388 1850
rect 34992 800 35020 1822
rect 35452 1442 35480 2790
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 35268 1414 35480 1442
rect 35268 800 35296 1414
rect 35544 800 35572 2450
rect 35820 800 35848 3470
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36096 800 36124 2382
rect 36372 800 36400 2790
rect 36648 800 36676 3470
rect 37188 2916 37240 2922
rect 37188 2858 37240 2864
rect 36912 2372 36964 2378
rect 36912 2314 36964 2320
rect 36924 800 36952 2314
rect 37200 800 37228 2858
rect 37476 800 37504 3470
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 37740 2848 37792 2854
rect 37740 2790 37792 2796
rect 37752 800 37780 2790
rect 38016 2576 38068 2582
rect 38016 2518 38068 2524
rect 38028 800 38056 2518
rect 38304 800 38332 2926
rect 38580 800 38608 3470
rect 39120 2916 39172 2922
rect 39120 2858 39172 2864
rect 38844 2508 38896 2514
rect 38844 2450 38896 2456
rect 38856 800 38884 2450
rect 39132 800 39160 2858
rect 39672 2848 39724 2854
rect 39672 2790 39724 2796
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39408 800 39436 2382
rect 39684 800 39712 2790
rect 39960 800 39988 3470
rect 40224 2916 40276 2922
rect 40224 2858 40276 2864
rect 40236 800 40264 2858
rect 40512 800 40540 3470
rect 40776 2508 40828 2514
rect 40776 2450 40828 2456
rect 40788 800 40816 2450
rect 41064 800 41092 3470
rect 42156 2984 42208 2990
rect 42156 2926 42208 2932
rect 41604 2848 41656 2854
rect 41604 2790 41656 2796
rect 41328 2440 41380 2446
rect 41328 2382 41380 2388
rect 41340 800 41368 2382
rect 41616 800 41644 2790
rect 41880 2576 41932 2582
rect 41880 2518 41932 2524
rect 41892 800 41920 2518
rect 42168 800 42196 2926
rect 42444 800 42472 3470
rect 42720 800 42748 3470
rect 42984 2916 43036 2922
rect 42984 2858 43036 2864
rect 44088 2916 44140 2922
rect 44088 2858 44140 2864
rect 42996 800 43024 2858
rect 43536 2848 43588 2854
rect 43536 2790 43588 2796
rect 43260 2508 43312 2514
rect 43260 2450 43312 2456
rect 43272 800 43300 2450
rect 43548 800 43576 2790
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 44100 800 44128 2858
rect 44376 800 44404 3470
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44640 2372 44692 2378
rect 44640 2314 44692 2320
rect 44652 800 44680 2314
rect 44928 800 44956 2790
rect 45204 800 45232 3470
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 45480 800 45508 2790
rect 45744 2576 45796 2582
rect 45744 2518 45796 2524
rect 45756 800 45784 2518
rect 46032 800 46060 3470
rect 46308 800 46336 3606
rect 50804 3596 50856 3602
rect 50804 3538 50856 3544
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 47400 2916 47452 2922
rect 47400 2858 47452 2864
rect 46848 2848 46900 2854
rect 46848 2790 46900 2796
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 46584 800 46612 2450
rect 46860 800 46888 2790
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 47136 800 47164 2382
rect 47412 800 47440 2858
rect 47688 800 47716 3470
rect 47952 2848 48004 2854
rect 47952 2790 48004 2796
rect 47964 800 47992 2790
rect 48240 800 48268 3470
rect 48780 2916 48832 2922
rect 48780 2858 48832 2864
rect 49884 2916 49936 2922
rect 49884 2858 49936 2864
rect 48504 2508 48556 2514
rect 48504 2450 48556 2456
rect 48516 800 48544 2450
rect 48792 800 48820 2858
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 49068 800 49096 2382
rect 49344 800 49372 2790
rect 49608 2576 49660 2582
rect 49608 2518 49660 2524
rect 49620 800 49648 2518
rect 49896 800 49924 2858
rect 50172 800 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1850 50660 3470
rect 50712 2848 50764 2854
rect 50712 2790 50764 2796
rect 50448 1822 50660 1850
rect 50448 800 50476 1822
rect 50724 1442 50752 2790
rect 50632 1414 50752 1442
rect 50632 800 50660 1414
rect 50816 1306 50844 3538
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50896 2440 50948 2446
rect 50896 2382 50948 2388
rect 50724 1278 50844 1306
rect 50724 800 50752 1278
rect 50908 1170 50936 2382
rect 50816 1142 50936 1170
rect 50816 800 50844 1142
rect 51000 1034 51028 2858
rect 50908 1006 51028 1034
rect 50908 800 50936 1006
rect 50988 944 51040 950
rect 50988 886 51040 892
rect 51000 800 51028 886
rect 51092 800 51120 3878
rect 51172 3528 51224 3534
rect 51172 3470 51224 3476
rect 51184 800 51212 3470
rect 51264 2304 51316 2310
rect 51264 2246 51316 2252
rect 51276 800 51304 2246
rect 51368 800 51396 3878
rect 51448 3664 51500 3670
rect 51448 3606 51500 3612
rect 51460 800 51488 3606
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 51540 2848 51592 2854
rect 51540 2790 51592 2796
rect 51552 800 51580 2790
rect 51644 800 51672 3538
rect 51724 3052 51776 3058
rect 51724 2994 51776 3000
rect 51736 800 51764 2994
rect 51828 800 51856 4014
rect 51908 3120 51960 3126
rect 51908 3062 51960 3068
rect 51920 800 51948 3062
rect 52000 2644 52052 2650
rect 52000 2586 52052 2592
rect 52012 800 52040 2586
rect 52104 800 52132 4558
rect 52196 800 52224 4694
rect 53196 4684 53248 4690
rect 53196 4626 53248 4632
rect 52644 4616 52696 4622
rect 52644 4558 52696 4564
rect 52460 3936 52512 3942
rect 52460 3878 52512 3884
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 52288 800 52316 3470
rect 52368 2100 52420 2106
rect 52368 2042 52420 2048
rect 52380 800 52408 2042
rect 52472 800 52500 3878
rect 52552 2440 52604 2446
rect 52552 2382 52604 2388
rect 52564 1154 52592 2382
rect 52552 1148 52604 1154
rect 52552 1090 52604 1096
rect 52552 944 52604 950
rect 52552 886 52604 892
rect 52564 800 52592 886
rect 52656 800 52684 4558
rect 53012 4140 53064 4146
rect 53012 4082 53064 4088
rect 52828 4004 52880 4010
rect 52828 3946 52880 3952
rect 52736 3732 52788 3738
rect 52736 3674 52788 3680
rect 52748 1426 52776 3674
rect 52736 1420 52788 1426
rect 52736 1362 52788 1368
rect 52840 1170 52868 3946
rect 53024 2774 53052 4082
rect 53104 2984 53156 2990
rect 53104 2926 53156 2932
rect 52748 1142 52868 1170
rect 52932 2746 53052 2774
rect 52748 800 52776 1142
rect 52932 1034 52960 2746
rect 53012 1420 53064 1426
rect 53012 1362 53064 1368
rect 52840 1006 52960 1034
rect 52840 800 52868 1006
rect 52920 944 52972 950
rect 52920 886 52972 892
rect 52932 800 52960 886
rect 53024 800 53052 1362
rect 53116 800 53144 2926
rect 53208 800 53236 4626
rect 53288 3460 53340 3466
rect 53288 3402 53340 3408
rect 53300 800 53328 3402
rect 53378 2952 53434 2961
rect 53378 2887 53434 2896
rect 53392 800 53420 2887
rect 53470 2816 53526 2825
rect 53470 2751 53526 2760
rect 53484 800 53512 2751
rect 53564 2032 53616 2038
rect 53564 1974 53616 1980
rect 53576 800 53604 1974
rect 53668 800 53696 4966
rect 53760 800 53788 5102
rect 54116 5092 54168 5098
rect 54116 5034 54168 5040
rect 53932 4752 53984 4758
rect 53932 4694 53984 4700
rect 53840 3596 53892 3602
rect 53840 3538 53892 3544
rect 53852 800 53880 3538
rect 53944 800 53972 4694
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 54036 800 54064 4014
rect 54128 800 54156 5034
rect 58164 5024 58216 5030
rect 58164 4966 58216 4972
rect 58176 4865 58204 4966
rect 58162 4856 58218 4865
rect 58162 4791 58218 4800
rect 54300 4684 54352 4690
rect 54300 4626 54352 4632
rect 54208 2916 54260 2922
rect 54208 2858 54260 2864
rect 54220 800 54248 2858
rect 54312 800 54340 4626
rect 55312 3936 55364 3942
rect 55312 3878 55364 3884
rect 58440 3936 58492 3942
rect 58440 3878 58492 3884
rect 54760 3052 54812 3058
rect 54760 2994 54812 3000
rect 54772 882 54800 2994
rect 55324 2825 55352 3878
rect 57520 3528 57572 3534
rect 58164 3528 58216 3534
rect 57520 3470 57572 3476
rect 58162 3496 58164 3505
rect 58216 3496 58218 3505
rect 56600 2984 56652 2990
rect 56598 2952 56600 2961
rect 56652 2952 56654 2961
rect 56598 2887 56654 2896
rect 55310 2816 55366 2825
rect 55310 2751 55366 2760
rect 55956 2440 56008 2446
rect 55956 2382 56008 2388
rect 56600 2440 56652 2446
rect 56600 2382 56652 2388
rect 55968 2106 55996 2382
rect 55956 2100 56008 2106
rect 55956 2042 56008 2048
rect 56612 1426 56640 2382
rect 57532 2145 57560 3470
rect 58162 3431 58218 3440
rect 57888 2508 57940 2514
rect 57888 2450 57940 2456
rect 57518 2136 57574 2145
rect 57518 2071 57574 2080
rect 57900 2038 57928 2450
rect 57888 2032 57940 2038
rect 57888 1974 57940 1980
rect 56600 1420 56652 1426
rect 56600 1362 56652 1368
rect 54760 876 54812 882
rect 54760 818 54812 824
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 58452 785 58480 3878
rect 58438 776 58494 785
rect 58438 711 58494 720
<< via2 >>
rect 58438 59200 58494 59256
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 57518 57840 57574 57896
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 57886 56480 57942 56536
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 58162 55140 58218 55176
rect 58162 55120 58164 55140
rect 58164 55120 58216 55140
rect 58216 55120 58218 55140
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 57886 53760 57942 53816
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 57886 52436 57888 52456
rect 57888 52436 57940 52456
rect 57940 52436 57942 52456
rect 57886 52400 57942 52436
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 58162 51040 58218 51096
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 58162 49716 58164 49736
rect 58164 49716 58216 49736
rect 58216 49716 58218 49736
rect 58162 49680 58218 49716
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 58162 48320 58218 48376
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 58162 46996 58164 47016
rect 58164 46996 58216 47016
rect 58216 46996 58218 47016
rect 58162 46960 58218 46996
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 58162 45600 58218 45656
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 58162 44260 58218 44296
rect 58162 44240 58164 44260
rect 58164 44240 58216 44260
rect 58216 44240 58218 44260
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 58162 42880 58218 42936
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4618 33360 4674 33416
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4986 33224 5042 33280
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1674 2896 1730 2952
rect 2410 5752 2466 5808
rect 2778 3168 2834 3224
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 5446 26288 5502 26344
rect 7194 26288 7250 26344
rect 5262 21936 5318 21992
rect 5722 19116 5724 19136
rect 5724 19116 5776 19136
rect 5776 19116 5778 19136
rect 5722 19080 5778 19116
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3974 8356 4030 8392
rect 3974 8336 3976 8356
rect 3976 8336 4028 8356
rect 4028 8336 4030 8356
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 3882 5480 3938 5536
rect 3790 4564 3792 4584
rect 3792 4564 3844 4584
rect 3844 4564 3846 4584
rect 3790 4528 3846 4564
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 5262 9324 5264 9344
rect 5264 9324 5316 9344
rect 5316 9324 5318 9344
rect 5262 9288 5318 9324
rect 5538 11076 5594 11112
rect 5538 11056 5540 11076
rect 5540 11056 5592 11076
rect 5592 11056 5594 11076
rect 5354 3884 5356 3904
rect 5356 3884 5408 3904
rect 5408 3884 5410 3904
rect 5354 3848 5410 3884
rect 5538 3984 5594 4040
rect 4986 3052 5042 3088
rect 4986 3032 4988 3052
rect 4988 3032 5040 3052
rect 5040 3032 5042 3052
rect 5354 2896 5410 2952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6458 13812 6460 13832
rect 6460 13812 6512 13832
rect 6512 13812 6514 13832
rect 6458 13776 6514 13812
rect 7654 16108 7710 16144
rect 7654 16088 7656 16108
rect 7656 16088 7708 16108
rect 7708 16088 7710 16108
rect 6642 11056 6698 11112
rect 5906 4528 5962 4584
rect 5814 3848 5870 3904
rect 5630 2624 5686 2680
rect 6182 2624 6238 2680
rect 10506 17620 10508 17640
rect 10508 17620 10560 17640
rect 10560 17620 10562 17640
rect 10506 17584 10562 17620
rect 9586 14220 9588 14240
rect 9588 14220 9640 14240
rect 9640 14220 9642 14240
rect 9586 14184 9642 14220
rect 6826 4276 6882 4312
rect 6826 4256 6828 4276
rect 6828 4256 6880 4276
rect 6880 4256 6882 4276
rect 6642 2644 6698 2680
rect 6642 2624 6644 2644
rect 6644 2624 6696 2644
rect 6696 2624 6698 2644
rect 7378 5752 7434 5808
rect 7838 5344 7894 5400
rect 8022 3984 8078 4040
rect 9310 9868 9312 9888
rect 9312 9868 9364 9888
rect 9364 9868 9366 9888
rect 9310 9832 9366 9868
rect 8758 5480 8814 5536
rect 8390 2896 8446 2952
rect 9310 4004 9366 4040
rect 9310 3984 9312 4004
rect 9312 3984 9364 4004
rect 9364 3984 9366 4004
rect 8850 3168 8906 3224
rect 9494 5752 9550 5808
rect 9494 5480 9550 5536
rect 9494 3052 9550 3088
rect 9494 3032 9496 3052
rect 9496 3032 9548 3052
rect 9548 3032 9550 3052
rect 11334 24132 11390 24168
rect 11334 24112 11336 24132
rect 11336 24112 11388 24132
rect 11388 24112 11390 24132
rect 11058 21936 11114 21992
rect 11702 23044 11758 23080
rect 11702 23024 11704 23044
rect 11704 23024 11756 23044
rect 11756 23024 11758 23044
rect 9862 2352 9918 2408
rect 10414 3168 10470 3224
rect 10966 3732 11022 3768
rect 10966 3712 10968 3732
rect 10968 3712 11020 3732
rect 11020 3712 11022 3732
rect 10966 3168 11022 3224
rect 11610 7520 11666 7576
rect 11242 3984 11298 4040
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 12346 24148 12348 24168
rect 12348 24148 12400 24168
rect 12400 24148 12402 24168
rect 12346 24112 12402 24148
rect 12898 24812 12954 24848
rect 12898 24792 12900 24812
rect 12900 24792 12952 24812
rect 12952 24792 12954 24812
rect 12162 21292 12164 21312
rect 12164 21292 12216 21312
rect 12216 21292 12218 21312
rect 12162 21256 12218 21292
rect 12806 20576 12862 20632
rect 12070 5616 12126 5672
rect 11518 2524 11520 2544
rect 11520 2524 11572 2544
rect 11572 2524 11574 2544
rect 11518 2488 11574 2524
rect 12714 10512 12770 10568
rect 13634 16632 13690 16688
rect 15198 18672 15254 18728
rect 13542 12824 13598 12880
rect 14646 12844 14702 12880
rect 14646 12824 14648 12844
rect 14648 12824 14700 12844
rect 14700 12824 14702 12844
rect 12530 8372 12532 8392
rect 12532 8372 12584 8392
rect 12584 8372 12586 8392
rect 12530 8336 12586 8372
rect 12530 8064 12586 8120
rect 12346 2352 12402 2408
rect 13266 8084 13322 8120
rect 13266 8064 13268 8084
rect 13268 8064 13320 8084
rect 13320 8064 13322 8084
rect 16854 18536 16910 18592
rect 17590 23024 17646 23080
rect 16946 16652 17002 16688
rect 16946 16632 16948 16652
rect 16948 16632 17000 16652
rect 17000 16632 17002 16652
rect 14922 5788 14924 5808
rect 14924 5788 14976 5808
rect 14976 5788 14978 5808
rect 14922 5752 14978 5788
rect 15198 6452 15254 6488
rect 15198 6432 15200 6452
rect 15200 6432 15252 6452
rect 15252 6432 15254 6452
rect 15566 6452 15622 6488
rect 15566 6432 15568 6452
rect 15568 6432 15620 6452
rect 15620 6432 15622 6452
rect 17590 18692 17646 18728
rect 17590 18672 17592 18692
rect 17592 18672 17644 18692
rect 17644 18672 17646 18692
rect 18326 24928 18382 24984
rect 14002 4256 14058 4312
rect 18234 18572 18236 18592
rect 18236 18572 18288 18592
rect 18288 18572 18290 18592
rect 18234 18536 18290 18572
rect 18050 17584 18106 17640
rect 18234 16632 18290 16688
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 18602 21528 18658 21584
rect 18602 20576 18658 20632
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19246 22208 19302 22264
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19890 18692 19946 18728
rect 19890 18672 19892 18692
rect 19892 18672 19944 18692
rect 19944 18672 19946 18692
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19706 18300 19708 18320
rect 19708 18300 19760 18320
rect 19760 18300 19762 18320
rect 19706 18264 19762 18300
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20258 18400 20314 18456
rect 20534 21800 20590 21856
rect 20442 18672 20498 18728
rect 20166 16632 20222 16688
rect 21086 25880 21142 25936
rect 23662 35980 23664 36000
rect 23664 35980 23716 36000
rect 23716 35980 23718 36000
rect 23662 35944 23718 35980
rect 22190 25900 22246 25936
rect 22190 25880 22192 25900
rect 22192 25880 22244 25900
rect 22244 25880 22246 25900
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20902 11600 20958 11656
rect 21730 14340 21786 14376
rect 21730 14320 21732 14340
rect 21732 14320 21784 14340
rect 21784 14320 21786 14340
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 58162 41556 58164 41576
rect 58164 41556 58216 41576
rect 58216 41556 58218 41576
rect 58162 41520 58218 41556
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 23754 24812 23810 24848
rect 23754 24792 23756 24812
rect 23756 24792 23808 24812
rect 23808 24792 23810 24812
rect 25226 32272 25282 32328
rect 24122 25880 24178 25936
rect 23386 21936 23442 21992
rect 25318 21936 25374 21992
rect 23202 16652 23258 16688
rect 23202 16632 23204 16652
rect 23204 16632 23256 16652
rect 23256 16632 23258 16652
rect 23202 16088 23258 16144
rect 19246 8336 19302 8392
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19522 7792 19578 7848
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19430 7384 19486 7440
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19062 5752 19118 5808
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19982 5228 20038 5264
rect 19982 5208 19984 5228
rect 19984 5208 20036 5228
rect 20036 5208 20038 5228
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20718 8372 20720 8392
rect 20720 8372 20772 8392
rect 20772 8372 20774 8392
rect 20718 8336 20774 8372
rect 25870 21936 25926 21992
rect 25042 15988 25044 16008
rect 25044 15988 25096 16008
rect 25096 15988 25098 16008
rect 25042 15952 25098 15988
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 26698 14320 26754 14376
rect 27986 16632 28042 16688
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 58162 40160 58218 40216
rect 29090 24656 29146 24712
rect 30654 28872 30710 28928
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 31758 31728 31814 31784
rect 32126 21800 32182 21856
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 32770 27376 32826 27432
rect 31942 21528 31998 21584
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 58162 38820 58218 38856
rect 58162 38800 58164 38820
rect 58164 38800 58216 38820
rect 58216 38800 58218 38820
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 58162 37440 58218 37496
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 58162 36116 58164 36136
rect 58164 36116 58216 36136
rect 58216 36116 58218 36136
rect 58162 36080 58218 36116
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 58162 34720 58218 34776
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 58162 33380 58218 33416
rect 58162 33360 58164 33380
rect 58164 33360 58216 33380
rect 58216 33360 58218 33380
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 58162 32000 58218 32056
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 58162 30676 58164 30696
rect 58164 30676 58216 30696
rect 58216 30676 58218 30696
rect 58162 30640 58218 30676
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 58162 29280 58218 29336
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 33782 27396 33838 27432
rect 33782 27376 33784 27396
rect 33784 27376 33836 27396
rect 33836 27376 33838 27396
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 33414 15952 33470 16008
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34610 10376 34666 10432
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34610 10104 34666 10160
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 58162 27940 58218 27976
rect 58162 27920 58164 27940
rect 58164 27920 58216 27940
rect 58216 27920 58218 27940
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 58162 26560 58218 26616
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 58162 25236 58164 25256
rect 58164 25236 58216 25256
rect 58216 25236 58218 25256
rect 58162 25200 58218 25236
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 58162 23840 58218 23896
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 58162 22500 58218 22536
rect 58162 22480 58164 22500
rect 58164 22480 58216 22500
rect 58216 22480 58218 22500
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 58162 21120 58218 21176
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 58162 19796 58164 19816
rect 58164 19796 58216 19816
rect 58216 19796 58218 19816
rect 58162 19760 58218 19796
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 58162 18400 58218 18456
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 58162 17060 58218 17096
rect 58162 17040 58164 17060
rect 58164 17040 58216 17060
rect 58216 17040 58218 17060
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 58162 15680 58218 15736
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 58162 14356 58164 14376
rect 58164 14356 58216 14376
rect 58216 14356 58218 14376
rect 58162 14320 58218 14356
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 58162 12960 58218 13016
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 58162 11620 58218 11656
rect 58162 11600 58164 11620
rect 58164 11600 58216 11620
rect 58216 11600 58218 11620
rect 36726 7404 36782 7440
rect 36726 7384 36728 7404
rect 36728 7384 36780 7404
rect 36780 7384 36782 7404
rect 37922 7404 37978 7440
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 58162 10240 58218 10296
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 58162 8916 58164 8936
rect 58164 8916 58216 8936
rect 58216 8916 58218 8936
rect 58162 8880 58218 8916
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 58162 7520 58218 7576
rect 37922 7384 37924 7404
rect 37924 7384 37976 7404
rect 37976 7384 37978 7404
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 58162 6180 58218 6216
rect 58162 6160 58164 6180
rect 58164 6160 58216 6180
rect 58216 6160 58218 6180
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 28998 2896 29054 2952
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 53378 2896 53434 2952
rect 53470 2760 53526 2816
rect 58162 4800 58218 4856
rect 58162 3476 58164 3496
rect 58164 3476 58216 3496
rect 58216 3476 58218 3496
rect 56598 2932 56600 2952
rect 56600 2932 56652 2952
rect 56652 2932 56654 2952
rect 56598 2896 56654 2932
rect 55310 2760 55366 2816
rect 58162 3440 58218 3476
rect 57518 2080 57574 2136
rect 58438 720 58494 776
<< metal3 >>
rect 58433 59258 58499 59261
rect 59200 59258 60000 59288
rect 58433 59256 60000 59258
rect 58433 59200 58438 59256
rect 58494 59200 60000 59256
rect 58433 59198 60000 59200
rect 58433 59195 58499 59198
rect 59200 59168 60000 59198
rect 57513 57898 57579 57901
rect 59200 57898 60000 57928
rect 57513 57896 60000 57898
rect 57513 57840 57518 57896
rect 57574 57840 60000 57896
rect 57513 57838 60000 57840
rect 57513 57835 57579 57838
rect 59200 57808 60000 57838
rect 19570 57696 19886 57697
rect 0 57536 800 57656
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 57881 56538 57947 56541
rect 59200 56538 60000 56568
rect 57881 56536 60000 56538
rect 57881 56480 57886 56536
rect 57942 56480 60000 56536
rect 57881 56478 60000 56480
rect 57881 56475 57947 56478
rect 59200 56448 60000 56478
rect 0 56040 800 56160
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 58157 55178 58223 55181
rect 59200 55178 60000 55208
rect 58157 55176 60000 55178
rect 58157 55120 58162 55176
rect 58218 55120 60000 55176
rect 58157 55118 60000 55120
rect 58157 55115 58223 55118
rect 59200 55088 60000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 0 54544 800 54664
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 57881 53818 57947 53821
rect 59200 53818 60000 53848
rect 57881 53816 60000 53818
rect 57881 53760 57886 53816
rect 57942 53760 60000 53816
rect 57881 53758 60000 53760
rect 57881 53755 57947 53758
rect 59200 53728 60000 53758
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 0 53048 800 53168
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 57881 52458 57947 52461
rect 59200 52458 60000 52488
rect 57881 52456 60000 52458
rect 57881 52400 57886 52456
rect 57942 52400 60000 52456
rect 57881 52398 60000 52400
rect 57881 52395 57947 52398
rect 59200 52368 60000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51552 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 58157 51098 58223 51101
rect 59200 51098 60000 51128
rect 58157 51096 60000 51098
rect 58157 51040 58162 51096
rect 58218 51040 60000 51096
rect 58157 51038 60000 51040
rect 58157 51035 58223 51038
rect 59200 51008 60000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 0 50056 800 50176
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 58157 49738 58223 49741
rect 59200 49738 60000 49768
rect 58157 49736 60000 49738
rect 58157 49680 58162 49736
rect 58218 49680 60000 49736
rect 58157 49678 60000 49680
rect 58157 49675 58223 49678
rect 59200 49648 60000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48560 800 48680
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58157 48378 58223 48381
rect 59200 48378 60000 48408
rect 58157 48376 60000 48378
rect 58157 48320 58162 48376
rect 58218 48320 60000 48376
rect 58157 48318 60000 48320
rect 58157 48315 58223 48318
rect 59200 48288 60000 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 0 47064 800 47184
rect 58157 47018 58223 47021
rect 59200 47018 60000 47048
rect 58157 47016 60000 47018
rect 58157 46960 58162 47016
rect 58218 46960 60000 47016
rect 58157 46958 60000 46960
rect 58157 46955 58223 46958
rect 59200 46928 60000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 0 45568 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 58157 45658 58223 45661
rect 59200 45658 60000 45688
rect 58157 45656 60000 45658
rect 58157 45600 58162 45656
rect 58218 45600 60000 45656
rect 58157 45598 60000 45600
rect 58157 45595 58223 45598
rect 59200 45568 60000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 58157 44298 58223 44301
rect 59200 44298 60000 44328
rect 58157 44296 60000 44298
rect 58157 44240 58162 44296
rect 58218 44240 60000 44296
rect 58157 44238 60000 44240
rect 58157 44235 58223 44238
rect 59200 44208 60000 44238
rect 0 44072 800 44192
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 58157 42938 58223 42941
rect 59200 42938 60000 42968
rect 58157 42936 60000 42938
rect 58157 42880 58162 42936
rect 58218 42880 60000 42936
rect 58157 42878 60000 42880
rect 58157 42875 58223 42878
rect 59200 42848 60000 42878
rect 0 42576 800 42696
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 58157 41578 58223 41581
rect 59200 41578 60000 41608
rect 58157 41576 60000 41578
rect 58157 41520 58162 41576
rect 58218 41520 60000 41576
rect 58157 41518 60000 41520
rect 58157 41515 58223 41518
rect 59200 41488 60000 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41080 800 41200
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 58157 40218 58223 40221
rect 59200 40218 60000 40248
rect 58157 40216 60000 40218
rect 58157 40160 58162 40216
rect 58218 40160 60000 40216
rect 58157 40158 60000 40160
rect 58157 40155 58223 40158
rect 59200 40128 60000 40158
rect 4210 39744 4526 39745
rect 0 39584 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 58157 38858 58223 38861
rect 59200 38858 60000 38888
rect 58157 38856 60000 38858
rect 58157 38800 58162 38856
rect 58218 38800 60000 38856
rect 58157 38798 60000 38800
rect 58157 38795 58223 38798
rect 59200 38768 60000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 0 38088 800 38208
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 58157 37498 58223 37501
rect 59200 37498 60000 37528
rect 58157 37496 60000 37498
rect 58157 37440 58162 37496
rect 58218 37440 60000 37496
rect 58157 37438 60000 37440
rect 58157 37435 58223 37438
rect 59200 37408 60000 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36592 800 36712
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 58157 36138 58223 36141
rect 59200 36138 60000 36168
rect 58157 36136 60000 36138
rect 58157 36080 58162 36136
rect 58218 36080 60000 36136
rect 58157 36078 60000 36080
rect 58157 36075 58223 36078
rect 59200 36048 60000 36078
rect 23657 36002 23723 36005
rect 23790 36002 23796 36004
rect 23657 36000 23796 36002
rect 23657 35944 23662 36000
rect 23718 35944 23796 36000
rect 23657 35942 23796 35944
rect 23657 35939 23723 35942
rect 23790 35940 23796 35942
rect 23860 35940 23866 36004
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 35096 800 35216
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 58157 34778 58223 34781
rect 59200 34778 60000 34808
rect 58157 34776 60000 34778
rect 58157 34720 58162 34776
rect 58218 34720 60000 34776
rect 58157 34718 60000 34720
rect 58157 34715 58223 34718
rect 59200 34688 60000 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 0 33600 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 4613 33418 4679 33421
rect 58157 33418 58223 33421
rect 59200 33418 60000 33448
rect 4613 33416 4722 33418
rect 4613 33360 4618 33416
rect 4674 33360 4722 33416
rect 4613 33355 4722 33360
rect 58157 33416 60000 33418
rect 58157 33360 58162 33416
rect 58218 33360 60000 33416
rect 58157 33358 60000 33360
rect 58157 33355 58223 33358
rect 4662 33282 4722 33355
rect 59200 33328 60000 33358
rect 4981 33282 5047 33285
rect 4662 33280 5047 33282
rect 4662 33224 4986 33280
rect 5042 33224 5047 33280
rect 4662 33222 5047 33224
rect 4981 33219 5047 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 24526 32268 24532 32332
rect 24596 32330 24602 32332
rect 25221 32330 25287 32333
rect 24596 32328 25287 32330
rect 24596 32272 25226 32328
rect 25282 32272 25287 32328
rect 24596 32270 25287 32272
rect 24596 32268 24602 32270
rect 25221 32267 25287 32270
rect 0 32104 800 32224
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 58157 32058 58223 32061
rect 59200 32058 60000 32088
rect 58157 32056 60000 32058
rect 58157 32000 58162 32056
rect 58218 32000 60000 32056
rect 58157 31998 60000 32000
rect 58157 31995 58223 31998
rect 59200 31968 60000 31998
rect 31753 31788 31819 31789
rect 31702 31786 31708 31788
rect 31626 31726 31708 31786
rect 31772 31786 31819 31788
rect 31772 31784 31864 31786
rect 31814 31728 31864 31784
rect 31702 31724 31708 31726
rect 31772 31726 31864 31728
rect 31772 31724 31819 31726
rect 31753 31723 31819 31724
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 0 30608 800 30728
rect 58157 30698 58223 30701
rect 59200 30698 60000 30728
rect 58157 30696 60000 30698
rect 58157 30640 58162 30696
rect 58218 30640 60000 30696
rect 58157 30638 60000 30640
rect 58157 30635 58223 30638
rect 59200 30608 60000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 58157 29338 58223 29341
rect 59200 29338 60000 29368
rect 58157 29336 60000 29338
rect 58157 29280 58162 29336
rect 58218 29280 60000 29336
rect 58157 29278 60000 29280
rect 58157 29275 58223 29278
rect 59200 29248 60000 29278
rect 0 29112 800 29232
rect 30649 28930 30715 28933
rect 31886 28930 31892 28932
rect 30649 28928 31892 28930
rect 30649 28872 30654 28928
rect 30710 28872 31892 28928
rect 30649 28870 31892 28872
rect 30649 28867 30715 28870
rect 31886 28868 31892 28870
rect 31956 28868 31962 28932
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 58157 27978 58223 27981
rect 59200 27978 60000 28008
rect 58157 27976 60000 27978
rect 58157 27920 58162 27976
rect 58218 27920 60000 27976
rect 58157 27918 60000 27920
rect 58157 27915 58223 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 0 27616 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 32765 27434 32831 27437
rect 33777 27434 33843 27437
rect 32765 27432 33843 27434
rect 32765 27376 32770 27432
rect 32826 27376 33782 27432
rect 33838 27376 33843 27432
rect 32765 27374 33843 27376
rect 32765 27371 32831 27374
rect 33777 27371 33843 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 58157 26618 58223 26621
rect 59200 26618 60000 26648
rect 58157 26616 60000 26618
rect 58157 26560 58162 26616
rect 58218 26560 60000 26616
rect 58157 26558 60000 26560
rect 58157 26555 58223 26558
rect 59200 26528 60000 26558
rect 5441 26346 5507 26349
rect 7189 26346 7255 26349
rect 5441 26344 7255 26346
rect 5441 26288 5446 26344
rect 5502 26288 7194 26344
rect 7250 26288 7255 26344
rect 5441 26286 7255 26288
rect 5441 26283 5507 26286
rect 7189 26283 7255 26286
rect 0 26120 800 26240
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 21081 25938 21147 25941
rect 22185 25938 22251 25941
rect 24117 25938 24183 25941
rect 21081 25936 24183 25938
rect 21081 25880 21086 25936
rect 21142 25880 22190 25936
rect 22246 25880 24122 25936
rect 24178 25880 24183 25936
rect 21081 25878 24183 25880
rect 21081 25875 21147 25878
rect 22185 25875 22251 25878
rect 24117 25875 24183 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 58157 25258 58223 25261
rect 59200 25258 60000 25288
rect 58157 25256 60000 25258
rect 58157 25200 58162 25256
rect 58218 25200 60000 25256
rect 58157 25198 60000 25200
rect 58157 25195 58223 25198
rect 59200 25168 60000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 11646 24924 11652 24988
rect 11716 24986 11722 24988
rect 18321 24986 18387 24989
rect 11716 24984 18387 24986
rect 11716 24928 18326 24984
rect 18382 24928 18387 24984
rect 11716 24926 18387 24928
rect 11716 24924 11722 24926
rect 18321 24923 18387 24926
rect 12893 24850 12959 24853
rect 23749 24852 23815 24853
rect 12893 24848 22110 24850
rect 12893 24792 12898 24848
rect 12954 24792 22110 24848
rect 12893 24790 22110 24792
rect 12893 24787 12959 24790
rect 0 24624 800 24744
rect 22050 24714 22110 24790
rect 23749 24848 23796 24852
rect 23860 24850 23866 24852
rect 23749 24792 23754 24848
rect 23749 24788 23796 24792
rect 23860 24790 23906 24850
rect 23860 24788 23866 24790
rect 23749 24787 23815 24788
rect 29085 24714 29151 24717
rect 22050 24712 29151 24714
rect 22050 24656 29090 24712
rect 29146 24656 29151 24712
rect 22050 24654 29151 24656
rect 29085 24651 29151 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 11329 24170 11395 24173
rect 12341 24170 12407 24173
rect 11329 24168 12407 24170
rect 11329 24112 11334 24168
rect 11390 24112 12346 24168
rect 12402 24112 12407 24168
rect 11329 24110 12407 24112
rect 11329 24107 11395 24110
rect 12341 24107 12407 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 58157 23898 58223 23901
rect 59200 23898 60000 23928
rect 58157 23896 60000 23898
rect 58157 23840 58162 23896
rect 58218 23840 60000 23896
rect 58157 23838 60000 23840
rect 58157 23835 58223 23838
rect 59200 23808 60000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23128 800 23248
rect 11697 23082 11763 23085
rect 17585 23082 17651 23085
rect 11697 23080 17651 23082
rect 11697 23024 11702 23080
rect 11758 23024 17590 23080
rect 17646 23024 17651 23080
rect 11697 23022 17651 23024
rect 11697 23019 11763 23022
rect 17585 23019 17651 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 58157 22538 58223 22541
rect 59200 22538 60000 22568
rect 58157 22536 60000 22538
rect 58157 22480 58162 22536
rect 58218 22480 60000 22536
rect 58157 22478 60000 22480
rect 58157 22475 58223 22478
rect 59200 22448 60000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19241 22268 19307 22269
rect 19190 22266 19196 22268
rect 19150 22206 19196 22266
rect 19260 22264 19307 22268
rect 19302 22208 19307 22264
rect 19190 22204 19196 22206
rect 19260 22204 19307 22208
rect 19241 22203 19307 22204
rect 5257 21994 5323 21997
rect 11053 21994 11119 21997
rect 5257 21992 11119 21994
rect 5257 21936 5262 21992
rect 5318 21936 11058 21992
rect 11114 21936 11119 21992
rect 5257 21934 11119 21936
rect 5257 21931 5323 21934
rect 11053 21931 11119 21934
rect 23381 21994 23447 21997
rect 24526 21994 24532 21996
rect 23381 21992 24532 21994
rect 23381 21936 23386 21992
rect 23442 21936 24532 21992
rect 23381 21934 24532 21936
rect 23381 21931 23447 21934
rect 24526 21932 24532 21934
rect 24596 21932 24602 21996
rect 25313 21994 25379 21997
rect 25865 21994 25931 21997
rect 25313 21992 25931 21994
rect 25313 21936 25318 21992
rect 25374 21936 25870 21992
rect 25926 21936 25931 21992
rect 25313 21934 25931 21936
rect 25313 21931 25379 21934
rect 25865 21931 25931 21934
rect 20529 21858 20595 21861
rect 32121 21858 32187 21861
rect 20529 21856 32187 21858
rect 20529 21800 20534 21856
rect 20590 21800 32126 21856
rect 32182 21800 32187 21856
rect 20529 21798 32187 21800
rect 20529 21795 20595 21798
rect 32121 21795 32187 21798
rect 19570 21792 19886 21793
rect 0 21632 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 18597 21586 18663 21589
rect 31937 21586 32003 21589
rect 18597 21584 32003 21586
rect 18597 21528 18602 21584
rect 18658 21528 31942 21584
rect 31998 21528 32003 21584
rect 18597 21526 32003 21528
rect 18597 21523 18663 21526
rect 31937 21523 32003 21526
rect 12157 21316 12223 21317
rect 12157 21314 12204 21316
rect 12112 21312 12204 21314
rect 12112 21256 12162 21312
rect 12112 21254 12204 21256
rect 12157 21252 12204 21254
rect 12268 21252 12274 21316
rect 12157 21251 12223 21252
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 58157 21178 58223 21181
rect 59200 21178 60000 21208
rect 58157 21176 60000 21178
rect 58157 21120 58162 21176
rect 58218 21120 60000 21176
rect 58157 21118 60000 21120
rect 58157 21115 58223 21118
rect 59200 21088 60000 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 12801 20634 12867 20637
rect 18597 20634 18663 20637
rect 12801 20632 18663 20634
rect 12801 20576 12806 20632
rect 12862 20576 18602 20632
rect 18658 20576 18663 20632
rect 12801 20574 18663 20576
rect 12801 20571 12867 20574
rect 18597 20571 18663 20574
rect 0 20136 800 20256
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 58157 19818 58223 19821
rect 59200 19818 60000 19848
rect 58157 19816 60000 19818
rect 58157 19760 58162 19816
rect 58218 19760 60000 19816
rect 58157 19758 60000 19760
rect 58157 19755 58223 19758
rect 59200 19728 60000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 5717 19140 5783 19141
rect 5717 19138 5764 19140
rect 5672 19136 5764 19138
rect 5672 19080 5722 19136
rect 5672 19078 5764 19080
rect 5717 19076 5764 19078
rect 5828 19076 5834 19140
rect 5717 19075 5783 19076
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 0 18640 800 18760
rect 15193 18730 15259 18733
rect 17585 18730 17651 18733
rect 15193 18728 17651 18730
rect 15193 18672 15198 18728
rect 15254 18672 17590 18728
rect 17646 18672 17651 18728
rect 15193 18670 17651 18672
rect 15193 18667 15259 18670
rect 17585 18667 17651 18670
rect 19885 18730 19951 18733
rect 20437 18730 20503 18733
rect 19885 18728 20503 18730
rect 19885 18672 19890 18728
rect 19946 18672 20442 18728
rect 20498 18672 20503 18728
rect 19885 18670 20503 18672
rect 19885 18667 19951 18670
rect 20437 18667 20503 18670
rect 16849 18594 16915 18597
rect 18229 18594 18295 18597
rect 16849 18592 18295 18594
rect 16849 18536 16854 18592
rect 16910 18536 18234 18592
rect 18290 18536 18295 18592
rect 16849 18534 18295 18536
rect 16849 18531 16915 18534
rect 18229 18531 18295 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 20253 18458 20319 18461
rect 20118 18456 20319 18458
rect 20118 18400 20258 18456
rect 20314 18400 20319 18456
rect 20118 18398 20319 18400
rect 19701 18322 19767 18325
rect 20118 18322 20178 18398
rect 20253 18395 20319 18398
rect 58157 18458 58223 18461
rect 59200 18458 60000 18488
rect 58157 18456 60000 18458
rect 58157 18400 58162 18456
rect 58218 18400 60000 18456
rect 58157 18398 60000 18400
rect 58157 18395 58223 18398
rect 59200 18368 60000 18398
rect 19701 18320 20178 18322
rect 19701 18264 19706 18320
rect 19762 18264 20178 18320
rect 19701 18262 20178 18264
rect 19701 18259 19767 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 10501 17642 10567 17645
rect 18045 17642 18111 17645
rect 10501 17640 18111 17642
rect 10501 17584 10506 17640
rect 10562 17584 18050 17640
rect 18106 17584 18111 17640
rect 10501 17582 18111 17584
rect 10501 17579 10567 17582
rect 18045 17579 18111 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 17144 800 17264
rect 58157 17098 58223 17101
rect 59200 17098 60000 17128
rect 58157 17096 60000 17098
rect 58157 17040 58162 17096
rect 58218 17040 60000 17096
rect 58157 17038 60000 17040
rect 58157 17035 58223 17038
rect 59200 17008 60000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 13629 16690 13695 16693
rect 16941 16690 17007 16693
rect 18229 16690 18295 16693
rect 20161 16690 20227 16693
rect 13629 16688 20227 16690
rect 13629 16632 13634 16688
rect 13690 16632 16946 16688
rect 17002 16632 18234 16688
rect 18290 16632 20166 16688
rect 20222 16632 20227 16688
rect 13629 16630 20227 16632
rect 13629 16627 13695 16630
rect 16941 16627 17007 16630
rect 18229 16627 18295 16630
rect 20161 16627 20227 16630
rect 23197 16690 23263 16693
rect 27981 16690 28047 16693
rect 23197 16688 28047 16690
rect 23197 16632 23202 16688
rect 23258 16632 27986 16688
rect 28042 16632 28047 16688
rect 23197 16630 28047 16632
rect 23197 16627 23263 16630
rect 27981 16627 28047 16630
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 7649 16146 7715 16149
rect 23197 16146 23263 16149
rect 7649 16144 23263 16146
rect 7649 16088 7654 16144
rect 7710 16088 23202 16144
rect 23258 16088 23263 16144
rect 7649 16086 23263 16088
rect 7649 16083 7715 16086
rect 23197 16083 23263 16086
rect 25037 16010 25103 16013
rect 33409 16010 33475 16013
rect 25037 16008 33475 16010
rect 25037 15952 25042 16008
rect 25098 15952 33414 16008
rect 33470 15952 33475 16008
rect 25037 15950 33475 15952
rect 25037 15947 25103 15950
rect 33409 15947 33475 15950
rect 4210 15808 4526 15809
rect 0 15648 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 58157 15738 58223 15741
rect 59200 15738 60000 15768
rect 58157 15736 60000 15738
rect 58157 15680 58162 15736
rect 58218 15680 60000 15736
rect 58157 15678 60000 15680
rect 58157 15675 58223 15678
rect 59200 15648 60000 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 21725 14378 21791 14381
rect 26693 14378 26759 14381
rect 21725 14376 26759 14378
rect 21725 14320 21730 14376
rect 21786 14320 26698 14376
rect 26754 14320 26759 14376
rect 21725 14318 26759 14320
rect 21725 14315 21791 14318
rect 26693 14315 26759 14318
rect 58157 14378 58223 14381
rect 59200 14378 60000 14408
rect 58157 14376 60000 14378
rect 58157 14320 58162 14376
rect 58218 14320 60000 14376
rect 58157 14318 60000 14320
rect 58157 14315 58223 14318
rect 59200 14288 60000 14318
rect 0 14152 800 14272
rect 5942 14180 5948 14244
rect 6012 14242 6018 14244
rect 9581 14242 9647 14245
rect 6012 14240 9647 14242
rect 6012 14184 9586 14240
rect 9642 14184 9647 14240
rect 6012 14182 9647 14184
rect 6012 14180 6018 14182
rect 9581 14179 9647 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 6453 13834 6519 13837
rect 10542 13834 10548 13836
rect 6453 13832 10548 13834
rect 6453 13776 6458 13832
rect 6514 13776 10548 13832
rect 6453 13774 10548 13776
rect 6453 13771 6519 13774
rect 10542 13772 10548 13774
rect 10612 13772 10618 13836
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 58157 13018 58223 13021
rect 59200 13018 60000 13048
rect 58157 13016 60000 13018
rect 58157 12960 58162 13016
rect 58218 12960 60000 13016
rect 58157 12958 60000 12960
rect 58157 12955 58223 12958
rect 59200 12928 60000 12958
rect 13537 12882 13603 12885
rect 14641 12882 14707 12885
rect 13537 12880 14707 12882
rect 13537 12824 13542 12880
rect 13598 12824 14646 12880
rect 14702 12824 14707 12880
rect 13537 12822 14707 12824
rect 13537 12819 13603 12822
rect 14641 12819 14707 12822
rect 0 12656 800 12776
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 7046 11596 7052 11660
rect 7116 11658 7122 11660
rect 20897 11658 20963 11661
rect 7116 11656 20963 11658
rect 7116 11600 20902 11656
rect 20958 11600 20963 11656
rect 7116 11598 20963 11600
rect 7116 11596 7122 11598
rect 20897 11595 20963 11598
rect 58157 11658 58223 11661
rect 59200 11658 60000 11688
rect 58157 11656 60000 11658
rect 58157 11600 58162 11656
rect 58218 11600 60000 11656
rect 58157 11598 60000 11600
rect 58157 11595 58223 11598
rect 59200 11568 60000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 11160 800 11280
rect 5533 11114 5599 11117
rect 6494 11114 6500 11116
rect 5533 11112 6500 11114
rect 5533 11056 5538 11112
rect 5594 11056 6500 11112
rect 5533 11054 6500 11056
rect 5533 11051 5599 11054
rect 6494 11052 6500 11054
rect 6564 11114 6570 11116
rect 6637 11114 6703 11117
rect 6564 11112 6703 11114
rect 6564 11056 6642 11112
rect 6698 11056 6703 11112
rect 6564 11054 6703 11056
rect 6564 11052 6570 11054
rect 6637 11051 6703 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 10726 10508 10732 10572
rect 10796 10570 10802 10572
rect 12709 10570 12775 10573
rect 10796 10568 12775 10570
rect 10796 10512 12714 10568
rect 12770 10512 12775 10568
rect 10796 10510 12775 10512
rect 10796 10508 10802 10510
rect 12709 10507 12775 10510
rect 34605 10434 34671 10437
rect 34605 10432 34714 10434
rect 34605 10376 34610 10432
rect 34666 10376 34714 10432
rect 34605 10371 34714 10376
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34654 10165 34714 10371
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 58157 10298 58223 10301
rect 59200 10298 60000 10328
rect 58157 10296 60000 10298
rect 58157 10240 58162 10296
rect 58218 10240 60000 10296
rect 58157 10238 60000 10240
rect 58157 10235 58223 10238
rect 59200 10208 60000 10238
rect 34605 10160 34714 10165
rect 34605 10104 34610 10160
rect 34666 10104 34714 10160
rect 34605 10102 34714 10104
rect 34605 10099 34671 10102
rect 8150 9828 8156 9892
rect 8220 9890 8226 9892
rect 9305 9890 9371 9893
rect 8220 9888 9371 9890
rect 8220 9832 9310 9888
rect 9366 9832 9371 9888
rect 8220 9830 9371 9832
rect 8220 9828 8226 9830
rect 9305 9827 9371 9830
rect 19570 9824 19886 9825
rect 0 9664 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 5257 9346 5323 9349
rect 5390 9346 5396 9348
rect 5257 9344 5396 9346
rect 5257 9288 5262 9344
rect 5318 9288 5396 9344
rect 5257 9286 5396 9288
rect 5257 9283 5323 9286
rect 5390 9284 5396 9286
rect 5460 9284 5466 9348
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 58157 8938 58223 8941
rect 59200 8938 60000 8968
rect 58157 8936 60000 8938
rect 58157 8880 58162 8936
rect 58218 8880 60000 8936
rect 58157 8878 60000 8880
rect 58157 8875 58223 8878
rect 59200 8848 60000 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 3969 8396 4035 8397
rect 3918 8332 3924 8396
rect 3988 8394 4035 8396
rect 3988 8392 4080 8394
rect 4030 8336 4080 8392
rect 3988 8334 4080 8336
rect 3988 8332 4035 8334
rect 10910 8332 10916 8396
rect 10980 8394 10986 8396
rect 12525 8394 12591 8397
rect 10980 8392 12591 8394
rect 10980 8336 12530 8392
rect 12586 8336 12591 8392
rect 10980 8334 12591 8336
rect 10980 8332 10986 8334
rect 3969 8331 4035 8332
rect 12525 8331 12591 8334
rect 19241 8394 19307 8397
rect 20713 8394 20779 8397
rect 19241 8392 20779 8394
rect 19241 8336 19246 8392
rect 19302 8336 20718 8392
rect 20774 8336 20779 8392
rect 19241 8334 20779 8336
rect 19241 8331 19307 8334
rect 20713 8331 20779 8334
rect 0 8168 800 8288
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 12525 8122 12591 8125
rect 13261 8122 13327 8125
rect 19190 8122 19196 8124
rect 12525 8120 19196 8122
rect 12525 8064 12530 8120
rect 12586 8064 13266 8120
rect 13322 8064 19196 8120
rect 12525 8062 19196 8064
rect 12525 8059 12591 8062
rect 13261 8059 13327 8062
rect 19190 8060 19196 8062
rect 19260 8060 19266 8124
rect 19517 7850 19583 7853
rect 19382 7848 19583 7850
rect 19382 7792 19522 7848
rect 19578 7792 19583 7848
rect 19382 7790 19583 7792
rect 11605 7580 11671 7581
rect 11605 7578 11652 7580
rect 11560 7576 11652 7578
rect 11560 7520 11610 7576
rect 11560 7518 11652 7520
rect 11605 7516 11652 7518
rect 11716 7516 11722 7580
rect 11605 7515 11671 7516
rect 19382 7445 19442 7790
rect 19517 7787 19583 7790
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 58157 7578 58223 7581
rect 59200 7578 60000 7608
rect 58157 7576 60000 7578
rect 58157 7520 58162 7576
rect 58218 7520 60000 7576
rect 58157 7518 60000 7520
rect 58157 7515 58223 7518
rect 59200 7488 60000 7518
rect 19382 7440 19491 7445
rect 19382 7384 19430 7440
rect 19486 7384 19491 7440
rect 19382 7382 19491 7384
rect 19425 7379 19491 7382
rect 36721 7442 36787 7445
rect 37917 7442 37983 7445
rect 36721 7440 37983 7442
rect 36721 7384 36726 7440
rect 36782 7384 37922 7440
rect 37978 7384 37983 7440
rect 36721 7382 37983 7384
rect 36721 7379 36787 7382
rect 37917 7379 37983 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6672 800 6792
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 15193 6490 15259 6493
rect 15561 6490 15627 6493
rect 15193 6488 15627 6490
rect 15193 6432 15198 6488
rect 15254 6432 15566 6488
rect 15622 6432 15627 6488
rect 15193 6430 15627 6432
rect 15193 6427 15259 6430
rect 15561 6427 15627 6430
rect 58157 6218 58223 6221
rect 59200 6218 60000 6248
rect 58157 6216 60000 6218
rect 58157 6160 58162 6216
rect 58218 6160 60000 6216
rect 58157 6158 60000 6160
rect 58157 6155 58223 6158
rect 59200 6128 60000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 2405 5810 2471 5813
rect 7373 5810 7439 5813
rect 9489 5810 9555 5813
rect 2405 5808 9555 5810
rect 2405 5752 2410 5808
rect 2466 5752 7378 5808
rect 7434 5752 9494 5808
rect 9550 5752 9555 5808
rect 2405 5750 9555 5752
rect 2405 5747 2471 5750
rect 7373 5747 7439 5750
rect 9489 5747 9555 5750
rect 14917 5810 14983 5813
rect 19057 5810 19123 5813
rect 14917 5808 19123 5810
rect 14917 5752 14922 5808
rect 14978 5752 19062 5808
rect 19118 5752 19123 5808
rect 14917 5750 19123 5752
rect 14917 5747 14983 5750
rect 19057 5747 19123 5750
rect 9622 5612 9628 5676
rect 9692 5674 9698 5676
rect 12065 5674 12131 5677
rect 9692 5672 12131 5674
rect 9692 5616 12070 5672
rect 12126 5616 12131 5672
rect 9692 5614 12131 5616
rect 9692 5612 9698 5614
rect 12065 5611 12131 5614
rect 3877 5538 3943 5541
rect 8753 5538 8819 5541
rect 9489 5538 9555 5541
rect 3877 5536 9555 5538
rect 3877 5480 3882 5536
rect 3938 5480 8758 5536
rect 8814 5480 9494 5536
rect 9550 5480 9555 5536
rect 3877 5478 9555 5480
rect 3877 5475 3943 5478
rect 8753 5475 8819 5478
rect 9489 5475 9555 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 7833 5404 7899 5405
rect 7782 5340 7788 5404
rect 7852 5402 7899 5404
rect 7852 5400 7944 5402
rect 7894 5344 7944 5400
rect 7852 5342 7944 5344
rect 7852 5340 7899 5342
rect 7833 5339 7899 5340
rect 0 5176 800 5296
rect 5574 5204 5580 5268
rect 5644 5266 5650 5268
rect 19977 5266 20043 5269
rect 5644 5264 20043 5266
rect 5644 5208 19982 5264
rect 20038 5208 20043 5264
rect 5644 5206 20043 5208
rect 5644 5204 5650 5206
rect 19977 5203 20043 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 58157 4858 58223 4861
rect 59200 4858 60000 4888
rect 58157 4856 60000 4858
rect 58157 4800 58162 4856
rect 58218 4800 60000 4856
rect 58157 4798 60000 4800
rect 58157 4795 58223 4798
rect 59200 4768 60000 4798
rect 3785 4586 3851 4589
rect 5901 4586 5967 4589
rect 3785 4584 5967 4586
rect 3785 4528 3790 4584
rect 3846 4528 5906 4584
rect 5962 4528 5967 4584
rect 3785 4526 5967 4528
rect 3785 4523 3851 4526
rect 5901 4523 5967 4526
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 6821 4314 6887 4317
rect 13997 4314 14063 4317
rect 6821 4312 14063 4314
rect 6821 4256 6826 4312
rect 6882 4256 14002 4312
rect 14058 4256 14063 4312
rect 6821 4254 14063 4256
rect 6821 4251 6887 4254
rect 13997 4251 14063 4254
rect 5533 4042 5599 4045
rect 7046 4042 7052 4044
rect 5533 4040 7052 4042
rect 5533 3984 5538 4040
rect 5594 3984 7052 4040
rect 5533 3982 7052 3984
rect 5533 3979 5599 3982
rect 7046 3980 7052 3982
rect 7116 3980 7122 4044
rect 8017 4042 8083 4045
rect 8150 4042 8156 4044
rect 8017 4040 8156 4042
rect 8017 3984 8022 4040
rect 8078 3984 8156 4040
rect 8017 3982 8156 3984
rect 8017 3979 8083 3982
rect 8150 3980 8156 3982
rect 8220 3980 8226 4044
rect 9305 4042 9371 4045
rect 11237 4042 11303 4045
rect 9305 4040 11303 4042
rect 9305 3984 9310 4040
rect 9366 3984 11242 4040
rect 11298 3984 11303 4040
rect 9305 3982 11303 3984
rect 9305 3979 9371 3982
rect 11237 3979 11303 3982
rect 5349 3906 5415 3909
rect 5574 3906 5580 3908
rect 5349 3904 5580 3906
rect 5349 3848 5354 3904
rect 5410 3848 5580 3904
rect 5349 3846 5580 3848
rect 5349 3843 5415 3846
rect 5574 3844 5580 3846
rect 5644 3844 5650 3908
rect 5809 3906 5875 3909
rect 5942 3906 5948 3908
rect 5809 3904 5948 3906
rect 5809 3848 5814 3904
rect 5870 3848 5948 3904
rect 5809 3846 5948 3848
rect 5809 3843 5875 3846
rect 5942 3844 5948 3846
rect 6012 3844 6018 3908
rect 4210 3840 4526 3841
rect 0 3680 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 10961 3772 11027 3773
rect 10910 3708 10916 3772
rect 10980 3770 11027 3772
rect 10980 3768 11072 3770
rect 11022 3712 11072 3768
rect 10980 3710 11072 3712
rect 10980 3708 11027 3710
rect 10961 3707 11027 3708
rect 58157 3498 58223 3501
rect 59200 3498 60000 3528
rect 58157 3496 60000 3498
rect 58157 3440 58162 3496
rect 58218 3440 60000 3496
rect 58157 3438 60000 3440
rect 58157 3435 58223 3438
rect 59200 3408 60000 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 2773 3226 2839 3229
rect 7782 3226 7788 3228
rect 2773 3224 7788 3226
rect 2773 3168 2778 3224
rect 2834 3168 7788 3224
rect 2773 3166 7788 3168
rect 2773 3163 2839 3166
rect 7782 3164 7788 3166
rect 7852 3226 7858 3228
rect 8845 3226 8911 3229
rect 7852 3224 8911 3226
rect 7852 3168 8850 3224
rect 8906 3168 8911 3224
rect 7852 3166 8911 3168
rect 7852 3164 7858 3166
rect 8845 3163 8911 3166
rect 10409 3226 10475 3229
rect 10542 3226 10548 3228
rect 10409 3224 10548 3226
rect 10409 3168 10414 3224
rect 10470 3168 10548 3224
rect 10409 3166 10548 3168
rect 10409 3163 10475 3166
rect 10542 3164 10548 3166
rect 10612 3164 10618 3228
rect 10726 3164 10732 3228
rect 10796 3226 10802 3228
rect 10961 3226 11027 3229
rect 10796 3224 11027 3226
rect 10796 3168 10966 3224
rect 11022 3168 11027 3224
rect 10796 3166 11027 3168
rect 10796 3164 10802 3166
rect 4981 3090 5047 3093
rect 9489 3090 9555 3093
rect 9622 3090 9628 3092
rect 4981 3088 8402 3090
rect 4981 3032 4986 3088
rect 5042 3032 8402 3088
rect 4981 3030 8402 3032
rect 4981 3027 5047 3030
rect 8342 2957 8402 3030
rect 9489 3088 9628 3090
rect 9489 3032 9494 3088
rect 9550 3032 9628 3088
rect 9489 3030 9628 3032
rect 9489 3027 9555 3030
rect 9622 3028 9628 3030
rect 9692 3028 9698 3092
rect 1669 2954 1735 2957
rect 5349 2954 5415 2957
rect 1669 2952 5415 2954
rect 1669 2896 1674 2952
rect 1730 2896 5354 2952
rect 5410 2896 5415 2952
rect 1669 2894 5415 2896
rect 8342 2952 8451 2957
rect 8342 2896 8390 2952
rect 8446 2896 8451 2952
rect 8342 2894 8451 2896
rect 10550 2954 10610 3164
rect 10961 3163 11027 3166
rect 28993 2954 29059 2957
rect 10550 2952 29059 2954
rect 10550 2896 28998 2952
rect 29054 2896 29059 2952
rect 10550 2894 29059 2896
rect 1669 2891 1735 2894
rect 5349 2891 5415 2894
rect 8385 2891 8451 2894
rect 28993 2891 29059 2894
rect 53373 2954 53439 2957
rect 56593 2954 56659 2957
rect 53373 2952 56659 2954
rect 53373 2896 53378 2952
rect 53434 2896 56598 2952
rect 56654 2896 56659 2952
rect 53373 2894 56659 2896
rect 53373 2891 53439 2894
rect 56593 2891 56659 2894
rect 53465 2818 53531 2821
rect 55305 2818 55371 2821
rect 53465 2816 55371 2818
rect 53465 2760 53470 2816
rect 53526 2760 55310 2816
rect 55366 2760 55371 2816
rect 53465 2758 55371 2760
rect 53465 2755 53531 2758
rect 55305 2755 55371 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 5625 2682 5691 2685
rect 6177 2682 6243 2685
rect 5625 2680 6243 2682
rect 5625 2624 5630 2680
rect 5686 2624 6182 2680
rect 6238 2624 6243 2680
rect 5625 2622 6243 2624
rect 5625 2619 5691 2622
rect 6177 2619 6243 2622
rect 6494 2620 6500 2684
rect 6564 2682 6570 2684
rect 6637 2682 6703 2685
rect 6564 2680 6703 2682
rect 6564 2624 6642 2680
rect 6698 2624 6703 2680
rect 6564 2622 6703 2624
rect 6564 2620 6570 2622
rect 6637 2619 6703 2622
rect 5390 2484 5396 2548
rect 5460 2546 5466 2548
rect 11513 2546 11579 2549
rect 5460 2544 11579 2546
rect 5460 2488 11518 2544
rect 11574 2488 11579 2544
rect 5460 2486 11579 2488
rect 5460 2484 5466 2486
rect 11513 2483 11579 2486
rect 3918 2348 3924 2412
rect 3988 2410 3994 2412
rect 9857 2410 9923 2413
rect 12198 2410 12204 2412
rect 3988 2408 12204 2410
rect 3988 2352 9862 2408
rect 9918 2352 12204 2408
rect 3988 2350 12204 2352
rect 3988 2348 3994 2350
rect 9857 2347 9923 2350
rect 12198 2348 12204 2350
rect 12268 2410 12274 2412
rect 12341 2410 12407 2413
rect 12268 2408 12407 2410
rect 12268 2352 12346 2408
rect 12402 2352 12407 2408
rect 12268 2350 12407 2352
rect 12268 2348 12274 2350
rect 12341 2347 12407 2350
rect 0 2184 800 2304
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 57513 2138 57579 2141
rect 59200 2138 60000 2168
rect 57513 2136 60000 2138
rect 57513 2080 57518 2136
rect 57574 2080 60000 2136
rect 57513 2078 60000 2080
rect 57513 2075 57579 2078
rect 59200 2048 60000 2078
rect 58433 778 58499 781
rect 59200 778 60000 808
rect 58433 776 60000 778
rect 58433 720 58438 776
rect 58494 720 60000 776
rect 58433 718 60000 720
rect 58433 715 58499 718
rect 59200 688 60000 718
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 23796 35940 23860 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 24532 32268 24596 32332
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 31708 31784 31772 31788
rect 31708 31728 31758 31784
rect 31758 31728 31772 31784
rect 31708 31724 31772 31728
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 31892 28868 31956 28932
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 11652 24924 11716 24988
rect 23796 24848 23860 24852
rect 23796 24792 23810 24848
rect 23810 24792 23860 24848
rect 23796 24788 23860 24792
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19196 22264 19260 22268
rect 19196 22208 19246 22264
rect 19246 22208 19260 22264
rect 19196 22204 19260 22208
rect 24532 21932 24596 21996
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 12204 21312 12268 21316
rect 12204 21256 12218 21312
rect 12218 21256 12268 21312
rect 12204 21252 12268 21256
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 5764 19136 5828 19140
rect 5764 19080 5778 19136
rect 5778 19080 5828 19136
rect 5764 19076 5828 19080
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 5948 14180 6012 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 10548 13772 10612 13836
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 7052 11596 7116 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 6500 11052 6564 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 10732 10508 10796 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 8156 9828 8220 9892
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 5396 9284 5460 9348
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 3924 8392 3988 8396
rect 3924 8336 3974 8392
rect 3974 8336 3988 8392
rect 3924 8332 3988 8336
rect 10916 8332 10980 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19196 8060 19260 8124
rect 11652 7576 11716 7580
rect 11652 7520 11666 7576
rect 11666 7520 11716 7576
rect 11652 7516 11716 7520
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 9628 5612 9692 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 7788 5400 7852 5404
rect 7788 5344 7838 5400
rect 7838 5344 7852 5400
rect 7788 5340 7852 5344
rect 5580 5204 5644 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 7052 3980 7116 4044
rect 8156 3980 8220 4044
rect 5580 3844 5644 3908
rect 5948 3844 6012 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 10916 3768 10980 3772
rect 10916 3712 10966 3768
rect 10966 3712 10980 3768
rect 10916 3708 10980 3712
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 7788 3164 7852 3228
rect 10548 3164 10612 3228
rect 10732 3164 10796 3228
rect 9628 3028 9692 3092
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 6500 2620 6564 2684
rect 5396 2484 5460 2548
rect 3924 2348 3988 2412
rect 12204 2348 12268 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 23795 36004 23861 36005
rect 23795 35940 23796 36004
rect 23860 35940 23861 36004
rect 23795 35939 23861 35940
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 11651 24988 11717 24989
rect 11651 24924 11652 24988
rect 11716 24924 11717 24988
rect 11651 24923 11717 24924
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 5763 19140 5829 19141
rect 5763 19076 5764 19140
rect 5828 19076 5829 19140
rect 5763 19075 5829 19076
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 5766 12450 5826 19075
rect 5947 14244 6013 14245
rect 5947 14180 5948 14244
rect 6012 14180 6013 14244
rect 5947 14179 6013 14180
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 5582 12390 5826 12450
rect 5395 9348 5461 9349
rect 5395 9284 5396 9348
rect 5460 9284 5461 9348
rect 5395 9283 5461 9284
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 3923 8396 3989 8397
rect 3923 8332 3924 8396
rect 3988 8332 3989 8396
rect 3923 8331 3989 8332
rect 3926 2413 3986 8331
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 3923 2412 3989 2413
rect 3923 2348 3924 2412
rect 3988 2348 3989 2412
rect 3923 2347 3989 2348
rect 4208 2128 4528 2688
rect 5398 2549 5458 9283
rect 5582 5269 5642 12390
rect 5579 5268 5645 5269
rect 5579 5204 5580 5268
rect 5644 5204 5645 5268
rect 5579 5203 5645 5204
rect 5582 3909 5642 5203
rect 5950 3909 6010 14179
rect 10547 13836 10613 13837
rect 10547 13772 10548 13836
rect 10612 13772 10613 13836
rect 10547 13771 10613 13772
rect 7051 11660 7117 11661
rect 7051 11596 7052 11660
rect 7116 11596 7117 11660
rect 7051 11595 7117 11596
rect 6499 11116 6565 11117
rect 6499 11052 6500 11116
rect 6564 11052 6565 11116
rect 6499 11051 6565 11052
rect 5579 3908 5645 3909
rect 5579 3844 5580 3908
rect 5644 3844 5645 3908
rect 5579 3843 5645 3844
rect 5947 3908 6013 3909
rect 5947 3844 5948 3908
rect 6012 3844 6013 3908
rect 5947 3843 6013 3844
rect 6502 2685 6562 11051
rect 7054 4045 7114 11595
rect 8155 9892 8221 9893
rect 8155 9828 8156 9892
rect 8220 9828 8221 9892
rect 8155 9827 8221 9828
rect 7787 5404 7853 5405
rect 7787 5340 7788 5404
rect 7852 5340 7853 5404
rect 7787 5339 7853 5340
rect 7051 4044 7117 4045
rect 7051 3980 7052 4044
rect 7116 3980 7117 4044
rect 7051 3979 7117 3980
rect 7790 3229 7850 5339
rect 8158 4045 8218 9827
rect 9627 5676 9693 5677
rect 9627 5612 9628 5676
rect 9692 5612 9693 5676
rect 9627 5611 9693 5612
rect 8155 4044 8221 4045
rect 8155 3980 8156 4044
rect 8220 3980 8221 4044
rect 8155 3979 8221 3980
rect 7787 3228 7853 3229
rect 7787 3164 7788 3228
rect 7852 3164 7853 3228
rect 7787 3163 7853 3164
rect 9630 3093 9690 5611
rect 10550 3229 10610 13771
rect 10731 10572 10797 10573
rect 10731 10508 10732 10572
rect 10796 10508 10797 10572
rect 10731 10507 10797 10508
rect 10734 3229 10794 10507
rect 10915 8396 10981 8397
rect 10915 8332 10916 8396
rect 10980 8332 10981 8396
rect 10915 8331 10981 8332
rect 10918 3773 10978 8331
rect 11654 7581 11714 24923
rect 19568 23968 19888 24992
rect 23798 24853 23858 35939
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 24531 32332 24597 32333
rect 24531 32268 24532 32332
rect 24596 32268 24597 32332
rect 24531 32267 24597 32268
rect 23795 24852 23861 24853
rect 23795 24788 23796 24852
rect 23860 24788 23861 24852
rect 23795 24787 23861 24788
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19195 22268 19261 22269
rect 19195 22204 19196 22268
rect 19260 22204 19261 22268
rect 19195 22203 19261 22204
rect 12203 21316 12269 21317
rect 12203 21252 12204 21316
rect 12268 21252 12269 21316
rect 12203 21251 12269 21252
rect 11651 7580 11717 7581
rect 11651 7516 11652 7580
rect 11716 7516 11717 7580
rect 11651 7515 11717 7516
rect 10915 3772 10981 3773
rect 10915 3708 10916 3772
rect 10980 3708 10981 3772
rect 10915 3707 10981 3708
rect 10547 3228 10613 3229
rect 10547 3164 10548 3228
rect 10612 3164 10613 3228
rect 10547 3163 10613 3164
rect 10731 3228 10797 3229
rect 10731 3164 10732 3228
rect 10796 3164 10797 3228
rect 10731 3163 10797 3164
rect 9627 3092 9693 3093
rect 9627 3028 9628 3092
rect 9692 3028 9693 3092
rect 9627 3027 9693 3028
rect 6499 2684 6565 2685
rect 6499 2620 6500 2684
rect 6564 2620 6565 2684
rect 6499 2619 6565 2620
rect 5395 2548 5461 2549
rect 5395 2484 5396 2548
rect 5460 2484 5461 2548
rect 5395 2483 5461 2484
rect 12206 2413 12266 21251
rect 19198 8125 19258 22203
rect 19568 21792 19888 22816
rect 24534 21997 24594 32267
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 31707 31788 31773 31789
rect 31707 31724 31708 31788
rect 31772 31770 31773 31788
rect 31772 31724 31954 31770
rect 31707 31723 31954 31724
rect 31710 31710 31954 31723
rect 31894 28933 31954 31710
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 31891 28932 31957 28933
rect 31891 28868 31892 28932
rect 31956 28868 31957 28932
rect 31891 28867 31957 28868
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 24531 21996 24597 21997
rect 24531 21932 24532 21996
rect 24596 21932 24597 21996
rect 24531 21931 24597 21932
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19195 8124 19261 8125
rect 19195 8060 19196 8124
rect 19260 8060 19261 8124
rect 19195 8059 19261 8060
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 12203 2412 12269 2413
rect 12203 2348 12204 2412
rect 12268 2348 12269 2412
rect 12203 2347 12269 2348
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B
timestamp 1649977179
transform 1 0 10304 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A0
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A0
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A0
timestamp 1649977179
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A0
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A0
timestamp 1649977179
transform 1 0 4508 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A0
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A0
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A0
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A0
timestamp 1649977179
transform 1 0 13524 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A0
timestamp 1649977179
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A0
timestamp 1649977179
transform 1 0 5152 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A0
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1649977179
transform -1 0 5336 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1649977179
transform 1 0 16836 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1649977179
transform 1 0 10488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B
timestamp 1649977179
transform -1 0 10120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1649977179
transform -1 0 12788 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1649977179
transform -1 0 12972 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1649977179
transform 1 0 4876 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1649977179
transform -1 0 5060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1649977179
transform -1 0 8372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1649977179
transform 1 0 3036 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1649977179
transform 1 0 5152 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1649977179
transform 1 0 3312 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1649977179
transform 1 0 6808 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1649977179
transform -1 0 5336 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1649977179
transform 1 0 7912 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1649977179
transform 1 0 26036 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1649977179
transform -1 0 12052 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1649977179
transform -1 0 14996 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A1
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1649977179
transform 1 0 23460 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1649977179
transform -1 0 21712 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1649977179
transform -1 0 13340 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1649977179
transform 1 0 21712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1649977179
transform 1 0 13432 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1649977179
transform 1 0 16008 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1649977179
transform 1 0 11868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1649977179
transform 1 0 13984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C1
timestamp 1649977179
transform 1 0 13432 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1649977179
transform 1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1649977179
transform 1 0 14628 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__C1
timestamp 1649977179
transform -1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1649977179
transform 1 0 28796 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1649977179
transform 1 0 30452 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1649977179
transform 1 0 28888 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1649977179
transform 1 0 27048 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__C1
timestamp 1649977179
transform 1 0 26496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1649977179
transform 1 0 26864 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__C1
timestamp 1649977179
transform 1 0 27048 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1649977179
transform 1 0 27140 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__C1
timestamp 1649977179
transform -1 0 28980 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1649977179
transform 1 0 29716 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1649977179
transform 1 0 29072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1
timestamp 1649977179
transform 1 0 35236 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp 1649977179
transform 1 0 35328 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1
timestamp 1649977179
transform 1 0 35236 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1649977179
transform 1 0 28244 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1649977179
transform 1 0 34960 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A1
timestamp 1649977179
transform 1 0 34868 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1649977179
transform -1 0 35144 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1649977179
transform 1 0 32476 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1649977179
transform 1 0 21160 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B
timestamp 1649977179
transform -1 0 21620 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1649977179
transform 1 0 28704 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1649977179
transform 1 0 30360 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1649977179
transform 1 0 29900 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1
timestamp 1649977179
transform 1 0 27140 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1649977179
transform -1 0 27416 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A1
timestamp 1649977179
transform 1 0 28888 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A1
timestamp 1649977179
transform 1 0 29900 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A1
timestamp 1649977179
transform 1 0 31280 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1649977179
transform 1 0 32292 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1649977179
transform 1 0 34776 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A1
timestamp 1649977179
transform 1 0 33396 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A1
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A1
timestamp 1649977179
transform 1 0 33672 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A1
timestamp 1649977179
transform 1 0 33580 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1649977179
transform 1 0 29716 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1649977179
transform -1 0 30636 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C1
timestamp 1649977179
transform 1 0 30636 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1649977179
transform -1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B
timestamp 1649977179
transform -1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1649977179
transform 1 0 14076 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1649977179
transform 1 0 16560 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1649977179
transform 1 0 5704 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__C1
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A1
timestamp 1649977179
transform 1 0 3128 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__C1
timestamp 1649977179
transform -1 0 5244 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C1
timestamp 1649977179
transform 1 0 5428 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1649977179
transform 1 0 4508 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__C1
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1649977179
transform 1 0 21896 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1649977179
transform -1 0 19780 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1649977179
transform 1 0 6900 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__C1
timestamp 1649977179
transform -1 0 8372 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1649977179
transform 1 0 20516 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__C1
timestamp 1649977179
transform 1 0 18584 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__C1
timestamp 1649977179
transform -1 0 20516 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1649977179
transform -1 0 17940 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__C1
timestamp 1649977179
transform -1 0 18676 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1649977179
transform 1 0 20700 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__C1
timestamp 1649977179
transform 1 0 19412 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A1
timestamp 1649977179
transform 1 0 20148 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1649977179
transform 1 0 14904 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1649977179
transform 1 0 17480 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B
timestamp 1649977179
transform 1 0 16928 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1649977179
transform -1 0 15548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1649977179
transform 1 0 9016 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1649977179
transform 1 0 10672 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1649977179
transform 1 0 23276 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1649977179
transform -1 0 12696 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A1
timestamp 1649977179
transform 1 0 12052 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__C1
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1649977179
transform 1 0 14168 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__C1
timestamp 1649977179
transform 1 0 16008 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A1
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__C1
timestamp 1649977179
transform -1 0 23644 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1649977179
transform 1 0 24288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__C1
timestamp 1649977179
transform -1 0 24196 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1649977179
transform 1 0 23736 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A1
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A1
timestamp 1649977179
transform 1 0 24472 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1649977179
transform 1 0 25208 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1649977179
transform 1 0 25024 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A1
timestamp 1649977179
transform 1 0 23736 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1649977179
transform 1 0 19596 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B
timestamp 1649977179
transform 1 0 19872 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1649977179
transform 1 0 25024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1649977179
transform 1 0 23000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1649977179
transform -1 0 24564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1649977179
transform -1 0 24840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1649977179
transform -1 0 16192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A1
timestamp 1649977179
transform 1 0 23368 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A1
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1
timestamp 1649977179
transform -1 0 26496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A1
timestamp 1649977179
transform 1 0 28888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1649977179
transform -1 0 31372 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1649977179
transform -1 0 33948 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A1
timestamp 1649977179
transform 1 0 31924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1649977179
transform 1 0 31924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform 1 0 29440 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1649977179
transform -1 0 29992 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1649977179
transform 1 0 26404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A1
timestamp 1649977179
transform -1 0 32568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1649977179
transform 1 0 26772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A1
timestamp 1649977179
transform -1 0 29072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1649977179
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1649977179
transform 1 0 19596 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A1
timestamp 1649977179
transform 1 0 22632 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1649977179
transform 1 0 20700 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B
timestamp 1649977179
transform 1 0 19688 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1649977179
transform -1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A1
timestamp 1649977179
transform -1 0 15456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A1
timestamp 1649977179
transform -1 0 15088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A1
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__C1
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A1
timestamp 1649977179
transform 1 0 18216 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__C1
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1
timestamp 1649977179
transform 1 0 31280 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__C1
timestamp 1649977179
transform 1 0 28796 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A1
timestamp 1649977179
transform 1 0 31188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__C1
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1
timestamp 1649977179
transform 1 0 30728 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__C1
timestamp 1649977179
transform -1 0 29716 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A1
timestamp 1649977179
transform -1 0 27232 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__C1
timestamp 1649977179
transform 1 0 26312 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1649977179
transform -1 0 27324 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__C1
timestamp 1649977179
transform 1 0 27324 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1649977179
transform 1 0 19872 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__C1
timestamp 1649977179
transform 1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1649977179
transform 1 0 20976 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__C1
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1649977179
transform -1 0 23920 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B
timestamp 1649977179
transform 1 0 22724 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1649977179
transform 1 0 34040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1649977179
transform 1 0 34040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1649977179
transform -1 0 35972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__C1
timestamp 1649977179
transform 1 0 34040 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A1
timestamp 1649977179
transform 1 0 36616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A1
timestamp 1649977179
transform 1 0 36616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A1
timestamp 1649977179
transform 1 0 37260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 1649977179
transform -1 0 39100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A1
timestamp 1649977179
transform 1 0 37076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A1
timestamp 1649977179
transform -1 0 40664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1
timestamp 1649977179
transform 1 0 38088 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1
timestamp 1649977179
transform 1 0 40204 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A1
timestamp 1649977179
transform -1 0 41124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A1
timestamp 1649977179
transform 1 0 37996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A1
timestamp 1649977179
transform 1 0 34040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1649977179
transform 1 0 21344 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B
timestamp 1649977179
transform 1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1649977179
transform -1 0 36340 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A
timestamp 1649977179
transform 1 0 34040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1
timestamp 1649977179
transform -1 0 33856 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A1
timestamp 1649977179
transform -1 0 33948 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A1
timestamp 1649977179
transform -1 0 35696 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1
timestamp 1649977179
transform 1 0 35512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1
timestamp 1649977179
transform 1 0 36524 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1649977179
transform 1 0 36616 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A1
timestamp 1649977179
transform 1 0 37352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__A1
timestamp 1649977179
transform 1 0 37352 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A1
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1649977179
transform 1 0 38088 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1649977179
transform 1 0 36616 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1649977179
transform 1 0 32752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1649977179
transform 1 0 21896 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1649977179
transform 1 0 27048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A
timestamp 1649977179
transform 1 0 26128 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A1
timestamp 1649977179
transform 1 0 25576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A1
timestamp 1649977179
transform -1 0 26864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A1
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1649977179
transform 1 0 27876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1649977179
transform -1 0 27508 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A1
timestamp 1649977179
transform 1 0 32476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1649977179
transform 1 0 13340 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1649977179
transform -1 0 25300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A1
timestamp 1649977179
transform 1 0 31464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A1
timestamp 1649977179
transform 1 0 32384 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A1
timestamp 1649977179
transform 1 0 33396 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A1
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1649977179
transform 1 0 25484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1649977179
transform -1 0 3312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1649977179
transform 1 0 16652 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1649977179
transform 1 0 19412 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1649977179
transform 1 0 7636 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A
timestamp 1649977179
transform -1 0 17020 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1649977179
transform 1 0 6532 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A
timestamp 1649977179
transform 1 0 5704 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A1
timestamp 1649977179
transform 1 0 4600 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1649977179
transform 1 0 4508 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A1
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1649977179
transform -1 0 2484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A
timestamp 1649977179
transform 1 0 5704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A1
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1649977179
transform 1 0 6440 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A1
timestamp 1649977179
transform 1 0 5244 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1649977179
transform 1 0 21160 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1649977179
transform 1 0 19320 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A
timestamp 1649977179
transform -1 0 20608 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1649977179
transform 1 0 21896 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 1649977179
transform 1 0 22724 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A1
timestamp 1649977179
transform -1 0 23828 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A1
timestamp 1649977179
transform -1 0 23276 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A
timestamp 1649977179
transform -1 0 20516 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1649977179
transform 1 0 20792 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 1649977179
transform 1 0 23460 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A1
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A
timestamp 1649977179
transform 1 0 12144 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__B
timestamp 1649977179
transform 1 0 19412 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A
timestamp 1649977179
transform 1 0 16192 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A1
timestamp 1649977179
transform 1 0 17204 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A2
timestamp 1649977179
transform 1 0 17664 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 1649977179
transform 1 0 12052 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__B
timestamp 1649977179
transform 1 0 18952 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1649977179
transform 1 0 18032 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A2
timestamp 1649977179
transform 1 0 18584 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1649977179
transform -1 0 19044 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1649977179
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1649977179
transform 1 0 15272 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1649977179
transform 1 0 16376 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A1
timestamp 1649977179
transform -1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 1649977179
transform 1 0 14076 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1649977179
transform -1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A1
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A1
timestamp 1649977179
transform 1 0 24472 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A1
timestamp 1649977179
transform 1 0 24564 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A1
timestamp 1649977179
transform -1 0 27140 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1649977179
transform -1 0 11040 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A1
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__C1
timestamp 1649977179
transform 1 0 23736 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__A1
timestamp 1649977179
transform -1 0 25208 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__C1
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A1
timestamp 1649977179
transform -1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__C1
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__A1
timestamp 1649977179
transform -1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__C1
timestamp 1649977179
transform -1 0 21988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1649977179
transform -1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 1649977179
transform 1 0 10396 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A
timestamp 1649977179
transform 1 0 14352 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A1
timestamp 1649977179
transform 1 0 5336 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__C1
timestamp 1649977179
transform 1 0 7820 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A1
timestamp 1649977179
transform -1 0 2760 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__C1
timestamp 1649977179
transform 1 0 4232 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1649977179
transform 1 0 5244 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__C1
timestamp 1649977179
transform -1 0 4876 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A1
timestamp 1649977179
transform 1 0 6348 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__C1
timestamp 1649977179
transform 1 0 8004 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A1
timestamp 1649977179
transform 1 0 5704 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__C1
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A1
timestamp 1649977179
transform 1 0 13524 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__C1
timestamp 1649977179
transform 1 0 11868 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A1
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A1
timestamp 1649977179
transform 1 0 16744 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A1
timestamp 1649977179
transform 1 0 18216 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A1
timestamp 1649977179
transform -1 0 17480 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A1
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A1
timestamp 1649977179
transform 1 0 12696 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A
timestamp 1649977179
transform 1 0 9752 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A1
timestamp 1649977179
transform -1 0 4324 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A1
timestamp 1649977179
transform 1 0 5060 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A1
timestamp 1649977179
transform -1 0 4140 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A1
timestamp 1649977179
transform -1 0 5244 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A1
timestamp 1649977179
transform 1 0 9936 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A1
timestamp 1649977179
transform -1 0 11316 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A1
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__A1
timestamp 1649977179
transform 1 0 11224 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A1
timestamp 1649977179
transform 1 0 11592 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__A1
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A1
timestamp 1649977179
transform -1 0 9292 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__A
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__A1
timestamp 1649977179
transform 1 0 9476 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A1
timestamp 1649977179
transform 1 0 9568 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A
timestamp 1649977179
transform 1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__A1
timestamp 1649977179
transform 1 0 11316 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A1
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A1
timestamp 1649977179
transform 1 0 13340 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A1
timestamp 1649977179
transform 1 0 21344 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__A1
timestamp 1649977179
transform -1 0 19780 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__A
timestamp 1649977179
transform -1 0 20240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A1
timestamp 1649977179
transform 1 0 21896 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__A1
timestamp 1649977179
transform -1 0 21344 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A1
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A1
timestamp 1649977179
transform -1 0 17756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A1
timestamp 1649977179
transform -1 0 17480 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__A
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__A
timestamp 1649977179
transform -1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__A
timestamp 1649977179
transform -1 0 20240 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__A
timestamp 1649977179
transform -1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A1
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A1
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__A1
timestamp 1649977179
transform 1 0 14628 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__A
timestamp 1649977179
transform -1 0 17940 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A1
timestamp 1649977179
transform -1 0 20884 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A1
timestamp 1649977179
transform -1 0 18492 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__A
timestamp 1649977179
transform -1 0 24932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__A1
timestamp 1649977179
transform 1 0 28888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__A1
timestamp 1649977179
transform 1 0 29624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A1
timestamp 1649977179
transform -1 0 31372 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A1
timestamp 1649977179
transform 1 0 26404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__A1
timestamp 1649977179
transform 1 0 25944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__A1
timestamp 1649977179
transform 1 0 17204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__C1
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A1
timestamp 1649977179
transform -1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__C1
timestamp 1649977179
transform -1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__D
timestamp 1649977179
transform 1 0 25576 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__C1
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__A
timestamp 1649977179
transform -1 0 23920 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__D
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__C1
timestamp 1649977179
transform 1 0 7636 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__A
timestamp 1649977179
transform 1 0 25300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__D
timestamp 1649977179
transform 1 0 25024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__C1
timestamp 1649977179
transform -1 0 7544 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__B2
timestamp 1649977179
transform -1 0 29072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__A
timestamp 1649977179
transform 1 0 31188 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__A
timestamp 1649977179
transform -1 0 30820 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__A2
timestamp 1649977179
transform 1 0 14628 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__B1
timestamp 1649977179
transform -1 0 15088 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__A
timestamp 1649977179
transform -1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__A1
timestamp 1649977179
transform 1 0 6624 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__A2
timestamp 1649977179
transform -1 0 17388 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__B1
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__A
timestamp 1649977179
transform 1 0 10120 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1620__A1
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__A2
timestamp 1649977179
transform -1 0 23920 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__B1
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1631__B
timestamp 1649977179
transform -1 0 15364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__A2
timestamp 1649977179
transform -1 0 22816 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__B1
timestamp 1649977179
transform 1 0 22356 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1646__B1
timestamp 1649977179
transform -1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__A2
timestamp 1649977179
transform 1 0 22632 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__B1
timestamp 1649977179
transform 1 0 22080 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1659__B1
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1671__B1
timestamp 1649977179
transform -1 0 11776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1683__B1
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1688__D
timestamp 1649977179
transform -1 0 25116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__B1
timestamp 1649977179
transform -1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1700__D
timestamp 1649977179
transform -1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1707__B1
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1708__A
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 20884 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_wb_clk_i_A
timestamp 1649977179
transform -1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_wb_clk_i_A
timestamp 1649977179
transform -1 0 12420 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 28336 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1649977179
transform 1 0 11592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1649977179
transform -1 0 16100 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1649977179
transform 1 0 12880 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1649977179
transform 1 0 7636 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1649977179
transform 1 0 7912 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1649977179
transform 1 0 5612 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1649977179
transform 1 0 20056 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1649977179
transform 1 0 15824 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1649977179
transform 1 0 25208 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1649977179
transform -1 0 30544 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1649977179
transform 1 0 34224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1649977179
transform 1 0 36616 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1649977179
transform 1 0 36432 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1649977179
transform 1 0 32568 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1649977179
transform -1 0 28704 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1649977179
transform 1 0 33396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1649977179
transform 1 0 39008 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1649977179
transform 1 0 35880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1649977179
transform 1 0 34040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_wb_clk_i_A
timestamp 1649977179
transform 1 0 31464 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_wb_clk_i_A
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_wb_clk_i_A
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_28_wb_clk_i_A
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_29_wb_clk_i_A
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_30_wb_clk_i_A
timestamp 1649977179
transform 1 0 17940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_31_wb_clk_i_A
timestamp 1649977179
transform 1 0 12144 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_32_wb_clk_i_A
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_33_wb_clk_i_A
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 2024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 8464 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 7912 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 16836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 4876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 4048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 6624 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 13432 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 9476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 10212 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output36_A
timestamp 1649977179
transform -1 0 2024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output37_A
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1649977179
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_171
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_178
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1649977179
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_323
timestamp 1649977179
transform 1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1649977179
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_340
timestamp 1649977179
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1649977179
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1649977179
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1649977179
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1649977179
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_17
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_72
timestamp 1649977179
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1649977179
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_143
timestamp 1649977179
transform 1 0 14260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_150
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_157
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_171
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1649977179
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_303
timestamp 1649977179
transform 1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1649977179
transform 1 0 29624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_324 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_340
timestamp 1649977179
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_354
timestamp 1649977179
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1649977179
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1649977179
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1649977179
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1649977179
transform 1 0 58512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1649977179
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp 1649977179
transform 1 0 11960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1649977179
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_183
timestamp 1649977179
transform 1 0 17940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_204
timestamp 1649977179
transform 1 0 19872 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_213
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_222
timestamp 1649977179
transform 1 0 21528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_226
timestamp 1649977179
transform 1 0 21896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_230
timestamp 1649977179
transform 1 0 22264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_237
timestamp 1649977179
transform 1 0 22908 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_246
timestamp 1649977179
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_258
timestamp 1649977179
transform 1 0 24840 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_267
timestamp 1649977179
transform 1 0 25668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1649977179
transform 1 0 27508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_294
timestamp 1649977179
transform 1 0 28152 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1649977179
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1649977179
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_376
timestamp 1649977179
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1649977179
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_390
timestamp 1649977179
transform 1 0 36984 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_399
timestamp 1649977179
transform 1 0 37812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_407
timestamp 1649977179
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1649977179
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1649977179
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_440
timestamp 1649977179
transform 1 0 41584 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_448
timestamp 1649977179
transform 1 0 42320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1649977179
transform 1 0 42780 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_460
timestamp 1649977179
transform 1 0 43424 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1649977179
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1649977179
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1649977179
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1649977179
transform 1 0 46552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_510
timestamp 1649977179
transform 1 0 48024 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_517
timestamp 1649977179
transform 1 0 48668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_529
timestamp 1649977179
transform 1 0 49772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_537
timestamp 1649977179
transform 1 0 50508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_544
timestamp 1649977179
transform 1 0 51152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_551
timestamp 1649977179
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_558
timestamp 1649977179
transform 1 0 52440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1649977179
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_610
timestamp 1649977179
transform 1 0 57224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_614
timestamp 1649977179
transform 1 0 57592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1649977179
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_9
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_16
timestamp 1649977179
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1649977179
transform 1 0 3956 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_75
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_97
timestamp 1649977179
transform 1 0 10028 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_117
timestamp 1649977179
transform 1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_124
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_138
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_152
timestamp 1649977179
transform 1 0 15088 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_158
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_197
timestamp 1649977179
transform 1 0 19228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1649977179
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_313
timestamp 1649977179
transform 1 0 29900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1649977179
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_368
timestamp 1649977179
transform 1 0 34960 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_380
timestamp 1649977179
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_547
timestamp 1649977179
transform 1 0 51428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_554
timestamp 1649977179
transform 1 0 52072 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_564
timestamp 1649977179
transform 1 0 52992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1649977179
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_578
timestamp 1649977179
transform 1 0 54280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_592
timestamp 1649977179
transform 1 0 55568 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_599
timestamp 1649977179
transform 1 0 56212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_611
timestamp 1649977179
transform 1 0 57316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1649977179
transform 1 0 58236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_10
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_39
timestamp 1649977179
transform 1 0 4692 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_49
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_61
timestamp 1649977179
transform 1 0 6716 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_123
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_130
timestamp 1649977179
transform 1 0 13064 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_145
timestamp 1649977179
transform 1 0 14444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_174
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_186
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_220
timestamp 1649977179
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_232
timestamp 1649977179
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1649977179
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_259
timestamp 1649977179
transform 1 0 24932 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_267
timestamp 1649977179
transform 1 0 25668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_272
timestamp 1649977179
transform 1 0 26128 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_284
timestamp 1649977179
transform 1 0 27232 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_293
timestamp 1649977179
transform 1 0 28060 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1649977179
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_313
timestamp 1649977179
transform 1 0 29900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_322
timestamp 1649977179
transform 1 0 30728 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_331
timestamp 1649977179
transform 1 0 31556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_343
timestamp 1649977179
transform 1 0 32660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1649977179
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_394
timestamp 1649977179
transform 1 0 37352 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_406
timestamp 1649977179
transform 1 0 38456 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_418
timestamp 1649977179
transform 1 0 39560 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_553
timestamp 1649977179
transform 1 0 51980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_558
timestamp 1649977179
transform 1 0 52440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_565
timestamp 1649977179
transform 1 0 53084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_572
timestamp 1649977179
transform 1 0 53728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_579
timestamp 1649977179
transform 1 0 54372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_592
timestamp 1649977179
transform 1 0 55568 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_599
timestamp 1649977179
transform 1 0 56212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_611
timestamp 1649977179
transform 1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1649977179
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_12
timestamp 1649977179
transform 1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_40
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_44
timestamp 1649977179
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_76
timestamp 1649977179
transform 1 0 8096 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_84
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1649977179
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_121
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_134
timestamp 1649977179
transform 1 0 13432 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_144
timestamp 1649977179
transform 1 0 14352 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1649977179
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1649977179
transform 1 0 18032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_188
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_209
timestamp 1649977179
transform 1 0 20332 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1649977179
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp 1649977179
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_269
timestamp 1649977179
transform 1 0 25852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1649977179
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_309
timestamp 1649977179
transform 1 0 29532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_312
timestamp 1649977179
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_324
timestamp 1649977179
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_376
timestamp 1649977179
transform 1 0 35696 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1649977179
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_569
timestamp 1649977179
transform 1 0 53452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_575
timestamp 1649977179
transform 1 0 54004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_582
timestamp 1649977179
transform 1 0 54648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_589
timestamp 1649977179
transform 1 0 55292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_601
timestamp 1649977179
transform 1 0 56396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_613
timestamp 1649977179
transform 1 0 57500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1649977179
transform 1 0 58236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_33
timestamp 1649977179
transform 1 0 4140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_39
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1649977179
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_64
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_91
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_104
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_115
timestamp 1649977179
transform 1 0 11684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_122
timestamp 1649977179
transform 1 0 12328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1649977179
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_154
timestamp 1649977179
transform 1 0 15272 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_174
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_180
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_183
timestamp 1649977179
transform 1 0 17940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_203
timestamp 1649977179
transform 1 0 19780 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_258
timestamp 1649977179
transform 1 0 24840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_270
timestamp 1649977179
transform 1 0 25944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1649977179
transform 1 0 26312 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_317
timestamp 1649977179
transform 1 0 30268 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_337
timestamp 1649977179
transform 1 0 32108 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_349
timestamp 1649977179
transform 1 0 33212 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_361
timestamp 1649977179
transform 1 0 34316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1649977179
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_374
timestamp 1649977179
transform 1 0 35512 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_380
timestamp 1649977179
transform 1 0 36064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_388
timestamp 1649977179
transform 1 0 36800 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_395
timestamp 1649977179
transform 1 0 37444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_407
timestamp 1649977179
transform 1 0 38548 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_37
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1649977179
transform 1 0 7360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_72
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_79
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1649977179
transform 1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_99
timestamp 1649977179
transform 1 0 10212 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_131
timestamp 1649977179
transform 1 0 13156 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_143
timestamp 1649977179
transform 1 0 14260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_174
timestamp 1649977179
transform 1 0 17112 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_186
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_199
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_211
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_230
timestamp 1649977179
transform 1 0 22264 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_238
timestamp 1649977179
transform 1 0 23000 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_257
timestamp 1649977179
transform 1 0 24748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_265
timestamp 1649977179
transform 1 0 25484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_298
timestamp 1649977179
transform 1 0 28520 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_311
timestamp 1649977179
transform 1 0 29716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_323
timestamp 1649977179
transform 1 0 30820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_357
timestamp 1649977179
transform 1 0 33948 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_369
timestamp 1649977179
transform 1 0 35052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_375
timestamp 1649977179
transform 1 0 35604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_384
timestamp 1649977179
transform 1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_397
timestamp 1649977179
transform 1 0 37628 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_414
timestamp 1649977179
transform 1 0 39192 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_426
timestamp 1649977179
transform 1 0 40296 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_438
timestamp 1649977179
transform 1 0 41400 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_446
timestamp 1649977179
transform 1 0 42136 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1649977179
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1649977179
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_19
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1649977179
transform 1 0 4048 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_48
timestamp 1649977179
transform 1 0 5520 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_60
timestamp 1649977179
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_64
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_74
timestamp 1649977179
transform 1 0 7912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1649977179
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_126
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1649977179
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_172
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_180
timestamp 1649977179
transform 1 0 17664 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_185
timestamp 1649977179
transform 1 0 18124 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_229
timestamp 1649977179
transform 1 0 22172 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp 1649977179
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1649977179
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_255
timestamp 1649977179
transform 1 0 24564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_259
timestamp 1649977179
transform 1 0 24932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_280
timestamp 1649977179
transform 1 0 26864 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_288
timestamp 1649977179
transform 1 0 27600 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_294
timestamp 1649977179
transform 1 0 28152 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1649977179
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_315
timestamp 1649977179
transform 1 0 30084 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_332
timestamp 1649977179
transform 1 0 31648 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_344
timestamp 1649977179
transform 1 0 32752 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_356
timestamp 1649977179
transform 1 0 33856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1649977179
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_369
timestamp 1649977179
transform 1 0 35052 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_390
timestamp 1649977179
transform 1 0 36984 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_398
timestamp 1649977179
transform 1 0 37720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp 1649977179
transform 1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1649977179
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1649977179
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1649977179
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1649977179
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_10
timestamp 1649977179
transform 1 0 2024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_30
timestamp 1649977179
transform 1 0 3864 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_38
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_41
timestamp 1649977179
transform 1 0 4876 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_49
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_59
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_88
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_91
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_97
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_116
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_146
timestamp 1649977179
transform 1 0 14536 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_154
timestamp 1649977179
transform 1 0 15272 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_174
timestamp 1649977179
transform 1 0 17112 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_186
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_200
timestamp 1649977179
transform 1 0 19504 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_236
timestamp 1649977179
transform 1 0 22816 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1649977179
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_260
timestamp 1649977179
transform 1 0 25024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_264
timestamp 1649977179
transform 1 0 25392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1649977179
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1649977179
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_283
timestamp 1649977179
transform 1 0 27140 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_291
timestamp 1649977179
transform 1 0 27876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_297
timestamp 1649977179
transform 1 0 28428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_326
timestamp 1649977179
transform 1 0 31096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1649977179
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_369
timestamp 1649977179
transform 1 0 35052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_380
timestamp 1649977179
transform 1 0 36064 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_388
timestamp 1649977179
transform 1 0 36800 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_401
timestamp 1649977179
transform 1 0 37996 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_410
timestamp 1649977179
transform 1 0 38824 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_422
timestamp 1649977179
transform 1 0 39928 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_434
timestamp 1649977179
transform 1 0 41032 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1649977179
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1649977179
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_19
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_31
timestamp 1649977179
transform 1 0 3956 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_45
timestamp 1649977179
transform 1 0 5244 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_55
timestamp 1649977179
transform 1 0 6164 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_71
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_74
timestamp 1649977179
transform 1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_99
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1649977179
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_127
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_164
timestamp 1649977179
transform 1 0 16192 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_172
timestamp 1649977179
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_183
timestamp 1649977179
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_202
timestamp 1649977179
transform 1 0 19688 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_208
timestamp 1649977179
transform 1 0 20240 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_220
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_228
timestamp 1649977179
transform 1 0 22080 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_238
timestamp 1649977179
transform 1 0 23000 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_244
timestamp 1649977179
transform 1 0 23552 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_285
timestamp 1649977179
transform 1 0 27324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1649977179
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_341
timestamp 1649977179
transform 1 0 32476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_360
timestamp 1649977179
transform 1 0 34224 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_370
timestamp 1649977179
transform 1 0 35144 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_382
timestamp 1649977179
transform 1 0 36248 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_388
timestamp 1649977179
transform 1 0 36800 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_400
timestamp 1649977179
transform 1 0 37904 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_412
timestamp 1649977179
transform 1 0 39008 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_617
timestamp 1649977179
transform 1 0 57868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1649977179
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_5
timestamp 1649977179
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_11
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_17
timestamp 1649977179
transform 1 0 2668 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_33
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_37
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_40
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_67
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_75
timestamp 1649977179
transform 1 0 8004 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_80
timestamp 1649977179
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_92
timestamp 1649977179
transform 1 0 9568 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_102
timestamp 1649977179
transform 1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_120
timestamp 1649977179
transform 1 0 12144 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_126
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_134
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_151
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_159
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_177
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_183
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_192
timestamp 1649977179
transform 1 0 18768 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_198
timestamp 1649977179
transform 1 0 19320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_209
timestamp 1649977179
transform 1 0 20332 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_215
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp 1649977179
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_239
timestamp 1649977179
transform 1 0 23092 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_251
timestamp 1649977179
transform 1 0 24196 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_255
timestamp 1649977179
transform 1 0 24564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_258
timestamp 1649977179
transform 1 0 24840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_270
timestamp 1649977179
transform 1 0 25944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1649977179
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_292
timestamp 1649977179
transform 1 0 27968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_304
timestamp 1649977179
transform 1 0 29072 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_315
timestamp 1649977179
transform 1 0 30084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_327
timestamp 1649977179
transform 1 0 31188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_353
timestamp 1649977179
transform 1 0 33580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_356
timestamp 1649977179
transform 1 0 33856 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_368
timestamp 1649977179
transform 1 0 34960 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_380
timestamp 1649977179
transform 1 0 36064 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1649977179
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1649977179
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1649977179
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_22
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_37
timestamp 1649977179
transform 1 0 4508 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_43
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_46
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_54
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_67
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_101
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_113
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_132
timestamp 1649977179
transform 1 0 13248 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_171
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_200
timestamp 1649977179
transform 1 0 19504 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1649977179
transform 1 0 20056 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_224
timestamp 1649977179
transform 1 0 21712 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_236
timestamp 1649977179
transform 1 0 22816 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_244
timestamp 1649977179
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_282
timestamp 1649977179
transform 1 0 27048 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_298
timestamp 1649977179
transform 1 0 28520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_328
timestamp 1649977179
transform 1 0 31280 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_340
timestamp 1649977179
transform 1 0 32384 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_352
timestamp 1649977179
transform 1 0 33488 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_399
timestamp 1649977179
transform 1 0 37812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_411
timestamp 1649977179
transform 1 0 38916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1649977179
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_617
timestamp 1649977179
transform 1 0 57868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1649977179
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_40
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_46
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_77
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_94
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1649977179
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_116
timestamp 1649977179
transform 1 0 11776 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_156
timestamp 1649977179
transform 1 0 15456 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1649977179
transform 1 0 17388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_183
timestamp 1649977179
transform 1 0 17940 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_191
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_199
timestamp 1649977179
transform 1 0 19412 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_206
timestamp 1649977179
transform 1 0 20056 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1649977179
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_233
timestamp 1649977179
transform 1 0 22540 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_250
timestamp 1649977179
transform 1 0 24104 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_259
timestamp 1649977179
transform 1 0 24932 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_268
timestamp 1649977179
transform 1 0 25760 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_284
timestamp 1649977179
transform 1 0 27232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_298
timestamp 1649977179
transform 1 0 28520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_306
timestamp 1649977179
transform 1 0 29256 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_319
timestamp 1649977179
transform 1 0 30452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_331
timestamp 1649977179
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_353
timestamp 1649977179
transform 1 0 33580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_368
timestamp 1649977179
transform 1 0 34960 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_376
timestamp 1649977179
transform 1 0 35696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1649977179
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1649977179
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_423
timestamp 1649977179
transform 1 0 40020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_435
timestamp 1649977179
transform 1 0 41124 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1649977179
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_11
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_17
timestamp 1649977179
transform 1 0 2668 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1649977179
transform 1 0 5428 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_58
timestamp 1649977179
transform 1 0 6440 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_69
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_129
timestamp 1649977179
transform 1 0 12972 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_168
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_176
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1649977179
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_192
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_203
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_230
timestamp 1649977179
transform 1 0 22264 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_236
timestamp 1649977179
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1649977179
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_256
timestamp 1649977179
transform 1 0 24656 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_262
timestamp 1649977179
transform 1 0 25208 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_274
timestamp 1649977179
transform 1 0 26312 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_282
timestamp 1649977179
transform 1 0 27048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_290
timestamp 1649977179
transform 1 0 27784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_319
timestamp 1649977179
transform 1 0 30452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_336
timestamp 1649977179
transform 1 0 32016 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_342
timestamp 1649977179
transform 1 0 32568 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_354
timestamp 1649977179
transform 1 0 33672 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1649977179
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_373
timestamp 1649977179
transform 1 0 35420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_379
timestamp 1649977179
transform 1 0 35972 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_383
timestamp 1649977179
transform 1 0 36340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_395
timestamp 1649977179
transform 1 0 37444 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_404
timestamp 1649977179
transform 1 0 38272 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_416
timestamp 1649977179
transform 1 0 39376 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_37
timestamp 1649977179
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1649977179
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_67
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_75
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_85
timestamp 1649977179
transform 1 0 8924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_97
timestamp 1649977179
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_117
timestamp 1649977179
transform 1 0 11868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1649977179
transform 1 0 18400 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_200
timestamp 1649977179
transform 1 0 19504 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_211
timestamp 1649977179
transform 1 0 20516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_232
timestamp 1649977179
transform 1 0 22448 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1649977179
transform 1 0 23184 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_263
timestamp 1649977179
transform 1 0 25300 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1649977179
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_287
timestamp 1649977179
transform 1 0 27508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1649977179
transform 1 0 28244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1649977179
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_330
timestamp 1649977179
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_345
timestamp 1649977179
transform 1 0 32844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_357
timestamp 1649977179
transform 1 0 33948 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_379
timestamp 1649977179
transform 1 0 35972 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_398
timestamp 1649977179
transform 1 0 37720 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_422
timestamp 1649977179
transform 1 0 39928 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_434
timestamp 1649977179
transform 1 0 41032 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_446
timestamp 1649977179
transform 1 0 42136 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1649977179
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_39
timestamp 1649977179
transform 1 0 4692 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_43
timestamp 1649977179
transform 1 0 5060 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_71
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_110
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_118
timestamp 1649977179
transform 1 0 11960 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_126
timestamp 1649977179
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_186
timestamp 1649977179
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1649977179
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_241
timestamp 1649977179
transform 1 0 23276 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1649977179
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_255
timestamp 1649977179
transform 1 0 24564 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1649977179
transform 1 0 25668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_275
timestamp 1649977179
transform 1 0 26404 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_282
timestamp 1649977179
transform 1 0 27048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_294
timestamp 1649977179
transform 1 0 28152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_298
timestamp 1649977179
transform 1 0 28520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_304
timestamp 1649977179
transform 1 0 29072 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_316
timestamp 1649977179
transform 1 0 30176 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_328
timestamp 1649977179
transform 1 0 31280 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_337
timestamp 1649977179
transform 1 0 32108 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_343
timestamp 1649977179
transform 1 0 32660 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_354
timestamp 1649977179
transform 1 0 33672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1649977179
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_372
timestamp 1649977179
transform 1 0 35328 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_380
timestamp 1649977179
transform 1 0 36064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_404
timestamp 1649977179
transform 1 0 38272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1649977179
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_21
timestamp 1649977179
transform 1 0 3036 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_38
timestamp 1649977179
transform 1 0 4600 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_73
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_94
timestamp 1649977179
transform 1 0 9752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_117
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_129
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_155
timestamp 1649977179
transform 1 0 15364 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_195
timestamp 1649977179
transform 1 0 19044 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1649977179
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_236
timestamp 1649977179
transform 1 0 22816 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_248
timestamp 1649977179
transform 1 0 23920 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_256
timestamp 1649977179
transform 1 0 24656 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1649977179
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_300
timestamp 1649977179
transform 1 0 28704 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_312
timestamp 1649977179
transform 1 0 29808 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_324
timestamp 1649977179
transform 1 0 30912 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1649977179
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_351
timestamp 1649977179
transform 1 0 33396 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_357
timestamp 1649977179
transform 1 0 33948 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_369
timestamp 1649977179
transform 1 0 35052 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_377
timestamp 1649977179
transform 1 0 35788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_383
timestamp 1649977179
transform 1 0 36340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_407
timestamp 1649977179
transform 1 0 38548 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_413
timestamp 1649977179
transform 1 0 39100 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_425
timestamp 1649977179
transform 1 0 40204 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_437
timestamp 1649977179
transform 1 0 41308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_445
timestamp 1649977179
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1649977179
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_54
timestamp 1649977179
transform 1 0 6072 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_103
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_186
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_199
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_219
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_225
timestamp 1649977179
transform 1 0 21804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_228
timestamp 1649977179
transform 1 0 22080 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_236
timestamp 1649977179
transform 1 0 22816 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1649977179
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_268
timestamp 1649977179
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_280
timestamp 1649977179
transform 1 0 26864 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_292
timestamp 1649977179
transform 1 0 27968 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1649977179
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_314
timestamp 1649977179
transform 1 0 29992 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_322
timestamp 1649977179
transform 1 0 30728 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_330
timestamp 1649977179
transform 1 0 31464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_350
timestamp 1649977179
transform 1 0 33304 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_360
timestamp 1649977179
transform 1 0 34224 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_373
timestamp 1649977179
transform 1 0 35420 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_385
timestamp 1649977179
transform 1 0 36524 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_397
timestamp 1649977179
transform 1 0 37628 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_403
timestamp 1649977179
transform 1 0 38180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_415
timestamp 1649977179
transform 1 0 39284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_16
timestamp 1649977179
transform 1 0 2576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1649977179
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_77
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_97
timestamp 1649977179
transform 1 0 10028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_132
timestamp 1649977179
transform 1 0 13248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1649977179
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_200
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_214
timestamp 1649977179
transform 1 0 20792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1649977179
transform 1 0 24748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_275
timestamp 1649977179
transform 1 0 26404 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_283
timestamp 1649977179
transform 1 0 27140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_301
timestamp 1649977179
transform 1 0 28796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_304
timestamp 1649977179
transform 1 0 29072 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_316
timestamp 1649977179
transform 1 0 30176 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_324
timestamp 1649977179
transform 1 0 30912 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_332
timestamp 1649977179
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_345
timestamp 1649977179
transform 1 0 32844 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_351
timestamp 1649977179
transform 1 0 33396 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_363
timestamp 1649977179
transform 1 0 34500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_367
timestamp 1649977179
transform 1 0 34868 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_378
timestamp 1649977179
transform 1 0 35880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_390
timestamp 1649977179
transform 1 0 36984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_398
timestamp 1649977179
transform 1 0 37720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1649977179
transform 1 0 38456 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_423
timestamp 1649977179
transform 1 0 40020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_435
timestamp 1649977179
transform 1 0 41124 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_112
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_124
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1649977179
transform 1 0 13064 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1649977179
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_156
timestamp 1649977179
transform 1 0 15456 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_164
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_200
timestamp 1649977179
transform 1 0 19504 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_206
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_212
timestamp 1649977179
transform 1 0 20608 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_220
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_237
timestamp 1649977179
transform 1 0 22908 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1649977179
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1649977179
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_276
timestamp 1649977179
transform 1 0 26496 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_280
timestamp 1649977179
transform 1 0 26864 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_311
timestamp 1649977179
transform 1 0 29716 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_323
timestamp 1649977179
transform 1 0 30820 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_337
timestamp 1649977179
transform 1 0 32108 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_343
timestamp 1649977179
transform 1 0 32660 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_354
timestamp 1649977179
transform 1 0 33672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1649977179
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_381
timestamp 1649977179
transform 1 0 36156 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_387
timestamp 1649977179
transform 1 0 36708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_411
timestamp 1649977179
transform 1 0 38916 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_425
timestamp 1649977179
transform 1 0 40204 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_437
timestamp 1649977179
transform 1 0 41308 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_449
timestamp 1649977179
transform 1 0 42412 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_461
timestamp 1649977179
transform 1 0 43516 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_473
timestamp 1649977179
transform 1 0 44620 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_617
timestamp 1649977179
transform 1 0 57868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1649977179
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_38
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_42
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_59
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_71
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_89
timestamp 1649977179
transform 1 0 9292 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_135
timestamp 1649977179
transform 1 0 13524 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_147
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_152
timestamp 1649977179
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_180
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_192
timestamp 1649977179
transform 1 0 18768 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_206
timestamp 1649977179
transform 1 0 20056 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_214
timestamp 1649977179
transform 1 0 20792 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1649977179
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_259
timestamp 1649977179
transform 1 0 24932 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_267
timestamp 1649977179
transform 1 0 25668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_285
timestamp 1649977179
transform 1 0 27324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1649977179
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_326
timestamp 1649977179
transform 1 0 31096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1649977179
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_345
timestamp 1649977179
transform 1 0 32844 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_350
timestamp 1649977179
transform 1 0 33304 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_362
timestamp 1649977179
transform 1 0 34408 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_401
timestamp 1649977179
transform 1 0 37996 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_425
timestamp 1649977179
transform 1 0 40204 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_437
timestamp 1649977179
transform 1 0 41308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_445
timestamp 1649977179
transform 1 0 42044 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_34
timestamp 1649977179
transform 1 0 4232 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_51
timestamp 1649977179
transform 1 0 5796 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_64
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_70
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1649977179
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1649977179
transform 1 0 11040 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_116
timestamp 1649977179
transform 1 0 11776 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_128
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_205
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_216
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_222
timestamp 1649977179
transform 1 0 21528 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1649977179
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_259
timestamp 1649977179
transform 1 0 24932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_274
timestamp 1649977179
transform 1 0 26312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_284
timestamp 1649977179
transform 1 0 27232 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_287
timestamp 1649977179
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1649977179
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_314
timestamp 1649977179
transform 1 0 29992 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_326
timestamp 1649977179
transform 1 0 31096 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_338
timestamp 1649977179
transform 1 0 32200 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_350
timestamp 1649977179
transform 1 0 33304 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_360
timestamp 1649977179
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_370
timestamp 1649977179
transform 1 0 35144 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_386
timestamp 1649977179
transform 1 0 36616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_394
timestamp 1649977179
transform 1 0 37352 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_410
timestamp 1649977179
transform 1 0 38824 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_418
timestamp 1649977179
transform 1 0 39560 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_431
timestamp 1649977179
transform 1 0 40756 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_443
timestamp 1649977179
transform 1 0 41860 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_455
timestamp 1649977179
transform 1 0 42964 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_467
timestamp 1649977179
transform 1 0 44068 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1649977179
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_617
timestamp 1649977179
transform 1 0 57868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1649977179
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1649977179
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_41
timestamp 1649977179
transform 1 0 4876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1649977179
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_85
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1649977179
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_124
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_136
timestamp 1649977179
transform 1 0 13616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_144
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1649977179
transform 1 0 17112 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1649977179
transform 1 0 17848 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_199
timestamp 1649977179
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1649977179
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_248
timestamp 1649977179
transform 1 0 23920 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_258
timestamp 1649977179
transform 1 0 24840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_271
timestamp 1649977179
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_313
timestamp 1649977179
transform 1 0 29900 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_325
timestamp 1649977179
transform 1 0 31004 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1649977179
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_353
timestamp 1649977179
transform 1 0 33580 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_357
timestamp 1649977179
transform 1 0 33948 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_360
timestamp 1649977179
transform 1 0 34224 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_369
timestamp 1649977179
transform 1 0 35052 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_381
timestamp 1649977179
transform 1 0 36156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1649977179
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1649977179
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_407
timestamp 1649977179
transform 1 0 38548 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_424
timestamp 1649977179
transform 1 0 40112 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_436
timestamp 1649977179
transform 1 0 41216 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_16
timestamp 1649977179
transform 1 0 2576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_20
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1649977179
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_34
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1649977179
transform 1 0 4784 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_52
timestamp 1649977179
transform 1 0 5888 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1649977179
transform 1 0 7452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1649977179
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 1649977179
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_104
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_116
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_122
timestamp 1649977179
transform 1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_130
timestamp 1649977179
transform 1 0 13064 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_204
timestamp 1649977179
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_213
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_225
timestamp 1649977179
transform 1 0 21804 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_230
timestamp 1649977179
transform 1 0 22264 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_238
timestamp 1649977179
transform 1 0 23000 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_246
timestamp 1649977179
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_255
timestamp 1649977179
transform 1 0 24564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_259
timestamp 1649977179
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_262
timestamp 1649977179
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_268
timestamp 1649977179
transform 1 0 25760 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1649977179
transform 1 0 26312 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_278
timestamp 1649977179
transform 1 0 26680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_284
timestamp 1649977179
transform 1 0 27232 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_292
timestamp 1649977179
transform 1 0 27968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_298
timestamp 1649977179
transform 1 0 28520 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1649977179
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_314
timestamp 1649977179
transform 1 0 29992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_326
timestamp 1649977179
transform 1 0 31096 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_346
timestamp 1649977179
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1649977179
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_370
timestamp 1649977179
transform 1 0 35144 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_383
timestamp 1649977179
transform 1 0 36340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_387
timestamp 1649977179
transform 1 0 36708 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1649977179
transform 1 0 37260 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_402
timestamp 1649977179
transform 1 0 38088 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_414
timestamp 1649977179
transform 1 0 39192 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1649977179
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1649977179
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1649977179
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1649977179
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_11
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_21
timestamp 1649977179
transform 1 0 3036 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_42
timestamp 1649977179
transform 1 0 4968 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1649977179
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_65
timestamp 1649977179
transform 1 0 7084 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_73
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_97
timestamp 1649977179
transform 1 0 10028 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_122
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_136
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_152
timestamp 1649977179
transform 1 0 15088 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_180
timestamp 1649977179
transform 1 0 17664 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_189
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_206
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_209
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_227
timestamp 1649977179
transform 1 0 21988 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_245
timestamp 1649977179
transform 1 0 23644 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_248
timestamp 1649977179
transform 1 0 23920 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_256
timestamp 1649977179
transform 1 0 24656 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_291
timestamp 1649977179
transform 1 0 27876 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_303
timestamp 1649977179
transform 1 0 28980 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_315
timestamp 1649977179
transform 1 0 30084 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1649977179
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_345
timestamp 1649977179
transform 1 0 32844 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_353
timestamp 1649977179
transform 1 0 33580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_365
timestamp 1649977179
transform 1 0 34684 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_369
timestamp 1649977179
transform 1 0 35052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_375
timestamp 1649977179
transform 1 0 35604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_387
timestamp 1649977179
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_396
timestamp 1649977179
transform 1 0 37536 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_404
timestamp 1649977179
transform 1 0 38272 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_416
timestamp 1649977179
transform 1 0 39376 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_428
timestamp 1649977179
transform 1 0 40480 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_440
timestamp 1649977179
transform 1 0 41584 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1649977179
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_33
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_43
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_58
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_70
timestamp 1649977179
transform 1 0 7544 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1649977179
transform 1 0 9660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_104
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_118
timestamp 1649977179
transform 1 0 11960 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1649977179
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1649977179
transform 1 0 14812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_156
timestamp 1649977179
transform 1 0 15456 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_164
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_168
timestamp 1649977179
transform 1 0 16560 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_174
timestamp 1649977179
transform 1 0 17112 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_180
timestamp 1649977179
transform 1 0 17664 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_187
timestamp 1649977179
transform 1 0 18308 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_205
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_212
timestamp 1649977179
transform 1 0 20608 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_222
timestamp 1649977179
transform 1 0 21528 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1649977179
transform 1 0 22080 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_235
timestamp 1649977179
transform 1 0 22724 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_242
timestamp 1649977179
transform 1 0 23368 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1649977179
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_259
timestamp 1649977179
transform 1 0 24932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_271
timestamp 1649977179
transform 1 0 26036 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_274
timestamp 1649977179
transform 1 0 26312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1649977179
transform 1 0 27140 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_291
timestamp 1649977179
transform 1 0 27876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_303
timestamp 1649977179
transform 1 0 28980 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_311
timestamp 1649977179
transform 1 0 29716 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_319
timestamp 1649977179
transform 1 0 30452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_331
timestamp 1649977179
transform 1 0 31556 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_337
timestamp 1649977179
transform 1 0 32108 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_343
timestamp 1649977179
transform 1 0 32660 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_346
timestamp 1649977179
transform 1 0 32936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_374
timestamp 1649977179
transform 1 0 35512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_394
timestamp 1649977179
transform 1 0 37352 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1649977179
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1649977179
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1649977179
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1649977179
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1649977179
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_24
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_32
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_40
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_62
timestamp 1649977179
transform 1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_75
timestamp 1649977179
transform 1 0 8004 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_87
timestamp 1649977179
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_91
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1649977179
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_116
timestamp 1649977179
transform 1 0 11776 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_124
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_136
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_142
timestamp 1649977179
transform 1 0 14168 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_154
timestamp 1649977179
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_186
timestamp 1649977179
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_198
timestamp 1649977179
transform 1 0 19320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_201
timestamp 1649977179
transform 1 0 19596 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1649977179
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_228
timestamp 1649977179
transform 1 0 22080 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1649977179
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_239
timestamp 1649977179
transform 1 0 23092 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_250
timestamp 1649977179
transform 1 0 24104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1649977179
transform 1 0 25024 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_264
timestamp 1649977179
transform 1 0 25392 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_267
timestamp 1649977179
transform 1 0 25668 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_283
timestamp 1649977179
transform 1 0 27140 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_295
timestamp 1649977179
transform 1 0 28244 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_307
timestamp 1649977179
transform 1 0 29348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1649977179
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1649977179
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_365
timestamp 1649977179
transform 1 0 34684 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_379
timestamp 1649977179
transform 1 0 35972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_403
timestamp 1649977179
transform 1 0 38180 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_411
timestamp 1649977179
transform 1 0 38916 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_414
timestamp 1649977179
transform 1 0 39192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_438
timestamp 1649977179
transform 1 0 41400 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_446
timestamp 1649977179
transform 1 0 42136 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1649977179
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_39
timestamp 1649977179
transform 1 0 4692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_51
timestamp 1649977179
transform 1 0 5796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_57
timestamp 1649977179
transform 1 0 6348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_60
timestamp 1649977179
transform 1 0 6624 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1649977179
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_91
timestamp 1649977179
transform 1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_95
timestamp 1649977179
transform 1 0 9844 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1649977179
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_104
timestamp 1649977179
transform 1 0 10672 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_111
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_115
timestamp 1649977179
transform 1 0 11684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1649977179
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1649977179
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_207
timestamp 1649977179
transform 1 0 20148 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_263
timestamp 1649977179
transform 1 0 25300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_275
timestamp 1649977179
transform 1 0 26404 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_287
timestamp 1649977179
transform 1 0 27508 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_299
timestamp 1649977179
transform 1 0 28612 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_312
timestamp 1649977179
transform 1 0 29808 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_316
timestamp 1649977179
transform 1 0 30176 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_323
timestamp 1649977179
transform 1 0 30820 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_335
timestamp 1649977179
transform 1 0 31924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_347
timestamp 1649977179
transform 1 0 33028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_359
timestamp 1649977179
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_374
timestamp 1649977179
transform 1 0 35512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_385
timestamp 1649977179
transform 1 0 36524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_396
timestamp 1649977179
transform 1 0 37536 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_404
timestamp 1649977179
transform 1 0 38272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_412
timestamp 1649977179
transform 1 0 39008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_429
timestamp 1649977179
transform 1 0 40572 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_435
timestamp 1649977179
transform 1 0 41124 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_447
timestamp 1649977179
transform 1 0 42228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_459
timestamp 1649977179
transform 1 0 43332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_471
timestamp 1649977179
transform 1 0 44436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1649977179
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_10
timestamp 1649977179
transform 1 0 2024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_30
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_36
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1649977179
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1649977179
transform 1 0 7636 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_89
timestamp 1649977179
transform 1 0 9292 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_116
timestamp 1649977179
transform 1 0 11776 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_128
timestamp 1649977179
transform 1 0 12880 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_140
timestamp 1649977179
transform 1 0 13984 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_152
timestamp 1649977179
transform 1 0 15088 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_158
timestamp 1649977179
transform 1 0 15640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_174
timestamp 1649977179
transform 1 0 17112 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_183
timestamp 1649977179
transform 1 0 17940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1649977179
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_213
timestamp 1649977179
transform 1 0 20700 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_228
timestamp 1649977179
transform 1 0 22080 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_242
timestamp 1649977179
transform 1 0 23368 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_253
timestamp 1649977179
transform 1 0 24380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_259
timestamp 1649977179
transform 1 0 24932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1649977179
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_297
timestamp 1649977179
transform 1 0 28428 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_311
timestamp 1649977179
transform 1 0 29716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_325
timestamp 1649977179
transform 1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1649977179
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_343
timestamp 1649977179
transform 1 0 32660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_353
timestamp 1649977179
transform 1 0 33580 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_377
timestamp 1649977179
transform 1 0 35788 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1649977179
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_397
timestamp 1649977179
transform 1 0 37628 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_425
timestamp 1649977179
transform 1 0 40204 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_434
timestamp 1649977179
transform 1 0 41032 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_446
timestamp 1649977179
transform 1 0 42136 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1649977179
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_38
timestamp 1649977179
transform 1 0 4600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_46
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_73
timestamp 1649977179
transform 1 0 7820 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1649977179
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_100
timestamp 1649977179
transform 1 0 10304 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_108
timestamp 1649977179
transform 1 0 11040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_113
timestamp 1649977179
transform 1 0 11500 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_119
timestamp 1649977179
transform 1 0 12052 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1649977179
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_170
timestamp 1649977179
transform 1 0 16744 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_190
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_199
timestamp 1649977179
transform 1 0 19412 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_211
timestamp 1649977179
transform 1 0 20516 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_219
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_223
timestamp 1649977179
transform 1 0 21620 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_235
timestamp 1649977179
transform 1 0 22724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_243
timestamp 1649977179
transform 1 0 23460 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1649977179
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_260
timestamp 1649977179
transform 1 0 25024 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_268
timestamp 1649977179
transform 1 0 25760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_275
timestamp 1649977179
transform 1 0 26404 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_284
timestamp 1649977179
transform 1 0 27232 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_296
timestamp 1649977179
transform 1 0 28336 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_316
timestamp 1649977179
transform 1 0 30176 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_322
timestamp 1649977179
transform 1 0 30728 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_339
timestamp 1649977179
transform 1 0 32292 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_351
timestamp 1649977179
transform 1 0 33396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_373
timestamp 1649977179
transform 1 0 35420 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_384
timestamp 1649977179
transform 1 0 36432 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_395
timestamp 1649977179
transform 1 0 37444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_407
timestamp 1649977179
transform 1 0 38548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_426
timestamp 1649977179
transform 1 0 40296 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_438
timestamp 1649977179
transform 1 0 41400 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_450
timestamp 1649977179
transform 1 0 42504 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_462
timestamp 1649977179
transform 1 0 43608 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_474
timestamp 1649977179
transform 1 0 44712 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_617
timestamp 1649977179
transform 1 0 57868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1649977179
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1649977179
transform 1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_25
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_35
timestamp 1649977179
transform 1 0 4324 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_43
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_46
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_60
timestamp 1649977179
transform 1 0 6624 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_72
timestamp 1649977179
transform 1 0 7728 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_84
timestamp 1649977179
transform 1 0 8832 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_92
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_98
timestamp 1649977179
transform 1 0 10120 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_102
timestamp 1649977179
transform 1 0 10488 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_121
timestamp 1649977179
transform 1 0 12236 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_132
timestamp 1649977179
transform 1 0 13248 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1649977179
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_148
timestamp 1649977179
transform 1 0 14720 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1649977179
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_182
timestamp 1649977179
transform 1 0 17848 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_189
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_195
timestamp 1649977179
transform 1 0 19044 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_207
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1649977179
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_284
timestamp 1649977179
transform 1 0 27232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_296
timestamp 1649977179
transform 1 0 28336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_304
timestamp 1649977179
transform 1 0 29072 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_312
timestamp 1649977179
transform 1 0 29808 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_320
timestamp 1649977179
transform 1 0 30544 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_339
timestamp 1649977179
transform 1 0 32292 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_343
timestamp 1649977179
transform 1 0 32660 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_360
timestamp 1649977179
transform 1 0 34224 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_382
timestamp 1649977179
transform 1 0 36248 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1649977179
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_423
timestamp 1649977179
transform 1 0 40020 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_435
timestamp 1649977179
transform 1 0 41124 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1649977179
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_16
timestamp 1649977179
transform 1 0 2576 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_45
timestamp 1649977179
transform 1 0 5244 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_50
timestamp 1649977179
transform 1 0 5704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1649977179
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_64
timestamp 1649977179
transform 1 0 6992 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1649977179
transform 1 0 8096 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_102
timestamp 1649977179
transform 1 0 10488 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_110
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1649977179
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_119
timestamp 1649977179
transform 1 0 12052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1649977179
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_143
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_149
timestamp 1649977179
transform 1 0 14812 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1649977179
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1649977179
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_227
timestamp 1649977179
transform 1 0 21988 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_231
timestamp 1649977179
transform 1 0 22356 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_237
timestamp 1649977179
transform 1 0 22908 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_249
timestamp 1649977179
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_273
timestamp 1649977179
transform 1 0 26220 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_294
timestamp 1649977179
transform 1 0 28152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1649977179
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_327
timestamp 1649977179
transform 1 0 31188 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_339
timestamp 1649977179
transform 1 0 32292 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_347
timestamp 1649977179
transform 1 0 33028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1649977179
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_376
timestamp 1649977179
transform 1 0 35696 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_388
timestamp 1649977179
transform 1 0 36800 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_400
timestamp 1649977179
transform 1 0 37904 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_412
timestamp 1649977179
transform 1 0 39008 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_427
timestamp 1649977179
transform 1 0 40388 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_439
timestamp 1649977179
transform 1 0 41492 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_451
timestamp 1649977179
transform 1 0 42596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_463
timestamp 1649977179
transform 1 0 43700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_617
timestamp 1649977179
transform 1 0 57868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1649977179
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_67
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_73
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_77
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1649977179
transform 1 0 9752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1649977179
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_118
timestamp 1649977179
transform 1 0 11960 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_130
timestamp 1649977179
transform 1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_143
timestamp 1649977179
transform 1 0 14260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1649977179
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1649977179
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_242
timestamp 1649977179
transform 1 0 23368 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_251
timestamp 1649977179
transform 1 0 24196 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_263
timestamp 1649977179
transform 1 0 25300 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_275
timestamp 1649977179
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_311
timestamp 1649977179
transform 1 0 29716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_325
timestamp 1649977179
transform 1 0 31004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_333
timestamp 1649977179
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_343
timestamp 1649977179
transform 1 0 32660 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_355
timestamp 1649977179
transform 1 0 33764 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_367
timestamp 1649977179
transform 1 0 34868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_375
timestamp 1649977179
transform 1 0 35604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_383
timestamp 1649977179
transform 1 0 36340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1649977179
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_49
timestamp 1649977179
transform 1 0 5612 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_70
timestamp 1649977179
transform 1 0 7544 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_76
timestamp 1649977179
transform 1 0 8096 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1649977179
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_94
timestamp 1649977179
transform 1 0 9752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_106
timestamp 1649977179
transform 1 0 10856 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_114
timestamp 1649977179
transform 1 0 11592 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_122
timestamp 1649977179
transform 1 0 12328 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp 1649977179
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1649977179
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_151
timestamp 1649977179
transform 1 0 14996 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_160
timestamp 1649977179
transform 1 0 15824 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_172
timestamp 1649977179
transform 1 0 16928 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_180
timestamp 1649977179
transform 1 0 17664 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1649977179
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_213
timestamp 1649977179
transform 1 0 20700 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_227
timestamp 1649977179
transform 1 0 21988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1649977179
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_256
timestamp 1649977179
transform 1 0 24656 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_262
timestamp 1649977179
transform 1 0 25208 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_282
timestamp 1649977179
transform 1 0 27048 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_297
timestamp 1649977179
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_305
timestamp 1649977179
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_318
timestamp 1649977179
transform 1 0 30360 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_329
timestamp 1649977179
transform 1 0 31372 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_341
timestamp 1649977179
transform 1 0 32476 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_353
timestamp 1649977179
transform 1 0 33580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1649977179
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_373
timestamp 1649977179
transform 1 0 35420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_382
timestamp 1649977179
transform 1 0 36248 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_386
timestamp 1649977179
transform 1 0 36616 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_392
timestamp 1649977179
transform 1 0 37168 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_404
timestamp 1649977179
transform 1 0 38272 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_416
timestamp 1649977179
transform 1 0 39376 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_426
timestamp 1649977179
transform 1 0 40296 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_438
timestamp 1649977179
transform 1 0 41400 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_450
timestamp 1649977179
transform 1 0 42504 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_462
timestamp 1649977179
transform 1 0 43608 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1649977179
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_11
timestamp 1649977179
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_30
timestamp 1649977179
transform 1 0 3864 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_50
timestamp 1649977179
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_67
timestamp 1649977179
transform 1 0 7268 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_73
timestamp 1649977179
transform 1 0 7820 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_90
timestamp 1649977179
transform 1 0 9384 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1649977179
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1649977179
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1649977179
transform 1 0 11684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_121
timestamp 1649977179
transform 1 0 12236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_129
timestamp 1649977179
transform 1 0 12972 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_135
timestamp 1649977179
transform 1 0 13524 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_147
timestamp 1649977179
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_156
timestamp 1649977179
transform 1 0 15456 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1649977179
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_171
timestamp 1649977179
transform 1 0 16836 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_175
timestamp 1649977179
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1649977179
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_190
timestamp 1649977179
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_199
timestamp 1649977179
transform 1 0 19412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_213
timestamp 1649977179
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1649977179
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_243
timestamp 1649977179
transform 1 0 23460 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_254
timestamp 1649977179
transform 1 0 24472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_266
timestamp 1649977179
transform 1 0 25576 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1649977179
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_287
timestamp 1649977179
transform 1 0 27508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_298
timestamp 1649977179
transform 1 0 28520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_306
timestamp 1649977179
transform 1 0 29256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_313
timestamp 1649977179
transform 1 0 29900 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_328
timestamp 1649977179
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_343
timestamp 1649977179
transform 1 0 32660 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_355
timestamp 1649977179
transform 1 0 33764 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_367
timestamp 1649977179
transform 1 0 34868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_371
timestamp 1649977179
transform 1 0 35236 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1649977179
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_401
timestamp 1649977179
transform 1 0 37996 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_425
timestamp 1649977179
transform 1 0 40204 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_437
timestamp 1649977179
transform 1 0 41308 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_445
timestamp 1649977179
transform 1 0 42044 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_621
timestamp 1649977179
transform 1 0 58236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_34
timestamp 1649977179
transform 1 0 4232 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_40
timestamp 1649977179
transform 1 0 4784 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_44
timestamp 1649977179
transform 1 0 5152 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_47
timestamp 1649977179
transform 1 0 5428 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_70
timestamp 1649977179
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1649977179
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_95
timestamp 1649977179
transform 1 0 9844 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_107
timestamp 1649977179
transform 1 0 10948 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_119
timestamp 1649977179
transform 1 0 12052 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_131
timestamp 1649977179
transform 1 0 13156 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1649977179
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_183
timestamp 1649977179
transform 1 0 17940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_202
timestamp 1649977179
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_208
timestamp 1649977179
transform 1 0 20240 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_214
timestamp 1649977179
transform 1 0 20792 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_217
timestamp 1649977179
transform 1 0 21068 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_223
timestamp 1649977179
transform 1 0 21620 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_226
timestamp 1649977179
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_236
timestamp 1649977179
transform 1 0 22816 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_242
timestamp 1649977179
transform 1 0 23368 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_255
timestamp 1649977179
transform 1 0 24564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_275
timestamp 1649977179
transform 1 0 26404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_281
timestamp 1649977179
transform 1 0 26956 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1649977179
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1649977179
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_315
timestamp 1649977179
transform 1 0 30084 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_323
timestamp 1649977179
transform 1 0 30820 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_329
timestamp 1649977179
transform 1 0 31372 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_341
timestamp 1649977179
transform 1 0 32476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_347
timestamp 1649977179
transform 1 0 33028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_353
timestamp 1649977179
transform 1 0 33580 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_361
timestamp 1649977179
transform 1 0 34316 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_373
timestamp 1649977179
transform 1 0 35420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_382
timestamp 1649977179
transform 1 0 36248 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_390
timestamp 1649977179
transform 1 0 36984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_393
timestamp 1649977179
transform 1 0 37260 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_404
timestamp 1649977179
transform 1 0 38272 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1649977179
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_429
timestamp 1649977179
transform 1 0 40572 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_438
timestamp 1649977179
transform 1 0 41400 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_450
timestamp 1649977179
transform 1 0 42504 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_462
timestamp 1649977179
transform 1 0 43608 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_474
timestamp 1649977179
transform 1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_11
timestamp 1649977179
transform 1 0 2116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_65
timestamp 1649977179
transform 1 0 7084 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_71
timestamp 1649977179
transform 1 0 7636 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_83
timestamp 1649977179
transform 1 0 8740 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_89
timestamp 1649977179
transform 1 0 9292 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_97
timestamp 1649977179
transform 1 0 10028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1649977179
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1649977179
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_202
timestamp 1649977179
transform 1 0 19688 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1649977179
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_241
timestamp 1649977179
transform 1 0 23276 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_255
timestamp 1649977179
transform 1 0 24564 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_264
timestamp 1649977179
transform 1 0 25392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_285
timestamp 1649977179
transform 1 0 27324 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_297
timestamp 1649977179
transform 1 0 28428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_310
timestamp 1649977179
transform 1 0 29624 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_318
timestamp 1649977179
transform 1 0 30360 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_330
timestamp 1649977179
transform 1 0 31464 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_342
timestamp 1649977179
transform 1 0 32568 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_346
timestamp 1649977179
transform 1 0 32936 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_355
timestamp 1649977179
transform 1 0 33764 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_367
timestamp 1649977179
transform 1 0 34868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_379
timestamp 1649977179
transform 1 0 35972 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_424
timestamp 1649977179
transform 1 0 40112 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_430
timestamp 1649977179
transform 1 0 40664 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_442
timestamp 1649977179
transform 1 0 41768 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_621
timestamp 1649977179
transform 1 0 58236 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1649977179
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_31
timestamp 1649977179
transform 1 0 3956 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_45
timestamp 1649977179
transform 1 0 5244 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_74
timestamp 1649977179
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1649977179
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_118
timestamp 1649977179
transform 1 0 11960 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_126
timestamp 1649977179
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1649977179
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_149
timestamp 1649977179
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_152
timestamp 1649977179
transform 1 0 15088 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_164
timestamp 1649977179
transform 1 0 16192 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_178
timestamp 1649977179
transform 1 0 17480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_213
timestamp 1649977179
transform 1 0 20700 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_237
timestamp 1649977179
transform 1 0 22908 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_249
timestamp 1649977179
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_256
timestamp 1649977179
transform 1 0 24656 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_268
timestamp 1649977179
transform 1 0 25760 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_280
timestamp 1649977179
transform 1 0 26864 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_284
timestamp 1649977179
transform 1 0 27232 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_329
timestamp 1649977179
transform 1 0 31372 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_332
timestamp 1649977179
transform 1 0 31648 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_344
timestamp 1649977179
transform 1 0 32752 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_353
timestamp 1649977179
transform 1 0 33580 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1649977179
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_381
timestamp 1649977179
transform 1 0 36156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_391
timestamp 1649977179
transform 1 0 37076 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_403
timestamp 1649977179
transform 1 0 38180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_415
timestamp 1649977179
transform 1 0 39284 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1649977179
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1649977179
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1649977179
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1649977179
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_11
timestamp 1649977179
transform 1 0 2116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_18
timestamp 1649977179
transform 1 0 2760 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1649977179
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_67
timestamp 1649977179
transform 1 0 7268 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_73
timestamp 1649977179
transform 1 0 7820 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_85
timestamp 1649977179
transform 1 0 8924 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_101
timestamp 1649977179
transform 1 0 10396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1649977179
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1649977179
transform 1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_135
timestamp 1649977179
transform 1 0 13524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_148
timestamp 1649977179
transform 1 0 14720 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_152
timestamp 1649977179
transform 1 0 15088 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1649977179
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_171
timestamp 1649977179
transform 1 0 16836 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_177
timestamp 1649977179
transform 1 0 17388 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_188
timestamp 1649977179
transform 1 0 18400 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_200
timestamp 1649977179
transform 1 0 19504 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_206
timestamp 1649977179
transform 1 0 20056 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1649977179
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_230
timestamp 1649977179
transform 1 0 22264 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_242
timestamp 1649977179
transform 1 0 23368 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_254
timestamp 1649977179
transform 1 0 24472 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_260
timestamp 1649977179
transform 1 0 25024 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_263
timestamp 1649977179
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_271
timestamp 1649977179
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_292
timestamp 1649977179
transform 1 0 27968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_304
timestamp 1649977179
transform 1 0 29072 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_315
timestamp 1649977179
transform 1 0 30084 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_327
timestamp 1649977179
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_381
timestamp 1649977179
transform 1 0 36156 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1649977179
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_399
timestamp 1649977179
transform 1 0 37812 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_416
timestamp 1649977179
transform 1 0 39376 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_428
timestamp 1649977179
transform 1 0 40480 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_440
timestamp 1649977179
transform 1 0 41584 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_49
timestamp 1649977179
transform 1 0 5612 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_52
timestamp 1649977179
transform 1 0 5888 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_59
timestamp 1649977179
transform 1 0 6532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_63
timestamp 1649977179
transform 1 0 6900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_80
timestamp 1649977179
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_40_98
timestamp 1649977179
transform 1 0 10120 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_106
timestamp 1649977179
transform 1 0 10856 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_112
timestamp 1649977179
transform 1 0 11408 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_124
timestamp 1649977179
transform 1 0 12512 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_130
timestamp 1649977179
transform 1 0 13064 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1649977179
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_143
timestamp 1649977179
transform 1 0 14260 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1649977179
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1649977179
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_164
timestamp 1649977179
transform 1 0 16192 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_170
timestamp 1649977179
transform 1 0 16744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1649977179
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_182
timestamp 1649977179
transform 1 0 17848 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1649977179
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_203
timestamp 1649977179
transform 1 0 19780 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_215
timestamp 1649977179
transform 1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_219
timestamp 1649977179
transform 1 0 21252 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_222
timestamp 1649977179
transform 1 0 21528 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_230
timestamp 1649977179
transform 1 0 22264 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_241
timestamp 1649977179
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_249
timestamp 1649977179
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_273
timestamp 1649977179
transform 1 0 26220 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_277
timestamp 1649977179
transform 1 0 26588 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_285
timestamp 1649977179
transform 1 0 27324 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_294
timestamp 1649977179
transform 1 0 28152 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_306
timestamp 1649977179
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_311
timestamp 1649977179
transform 1 0 29716 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_323
timestamp 1649977179
transform 1 0 30820 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_329
timestamp 1649977179
transform 1 0 31372 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_337
timestamp 1649977179
transform 1 0 32108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1649977179
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_354
timestamp 1649977179
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1649977179
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_383
timestamp 1649977179
transform 1 0 36340 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_386
timestamp 1649977179
transform 1 0 36616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_410
timestamp 1649977179
transform 1 0 38824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1649977179
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1649977179
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1649977179
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1649977179
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_617
timestamp 1649977179
transform 1 0 57868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1649977179
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_32
timestamp 1649977179
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1649977179
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_61
timestamp 1649977179
transform 1 0 6716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_73
timestamp 1649977179
transform 1 0 7820 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_79
timestamp 1649977179
transform 1 0 8372 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_96
timestamp 1649977179
transform 1 0 9936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1649977179
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_115
timestamp 1649977179
transform 1 0 11684 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_121
timestamp 1649977179
transform 1 0 12236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_133
timestamp 1649977179
transform 1 0 13340 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_141
timestamp 1649977179
transform 1 0 14076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_144
timestamp 1649977179
transform 1 0 14352 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_156
timestamp 1649977179
transform 1 0 15456 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1649977179
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_173
timestamp 1649977179
transform 1 0 17020 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_185
timestamp 1649977179
transform 1 0 18124 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_201
timestamp 1649977179
transform 1 0 19596 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_210
timestamp 1649977179
transform 1 0 20424 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1649977179
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_247
timestamp 1649977179
transform 1 0 23828 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_257
timestamp 1649977179
transform 1 0 24748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_268
timestamp 1649977179
transform 1 0 25760 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1649977179
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_284
timestamp 1649977179
transform 1 0 27232 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_296
timestamp 1649977179
transform 1 0 28336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_300
timestamp 1649977179
transform 1 0 28704 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_303
timestamp 1649977179
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_312
timestamp 1649977179
transform 1 0 29808 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1649977179
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_355
timestamp 1649977179
transform 1 0 33764 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_372
timestamp 1649977179
transform 1 0 35328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_384
timestamp 1649977179
transform 1 0 36432 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_396
timestamp 1649977179
transform 1 0 37536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_408
timestamp 1649977179
transform 1 0 38640 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1649977179
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1649977179
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1649977179
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1649977179
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_67
timestamp 1649977179
transform 1 0 7268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_73
timestamp 1649977179
transform 1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1649977179
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_88
timestamp 1649977179
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_100
timestamp 1649977179
transform 1 0 10304 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_106
timestamp 1649977179
transform 1 0 10856 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_118
timestamp 1649977179
transform 1 0 11960 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1649977179
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_145
timestamp 1649977179
transform 1 0 14444 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_171
timestamp 1649977179
transform 1 0 16836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_183
timestamp 1649977179
transform 1 0 17940 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1649977179
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_213
timestamp 1649977179
transform 1 0 20700 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_225
timestamp 1649977179
transform 1 0 21804 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_285
timestamp 1649977179
transform 1 0 27324 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_297
timestamp 1649977179
transform 1 0 28428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1649977179
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_320
timestamp 1649977179
transform 1 0 30544 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_340
timestamp 1649977179
transform 1 0 32384 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_352
timestamp 1649977179
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_383
timestamp 1649977179
transform 1 0 36340 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_393
timestamp 1649977179
transform 1 0 37260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_396
timestamp 1649977179
transform 1 0 37536 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_408
timestamp 1649977179
transform 1 0 38640 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_617
timestamp 1649977179
transform 1 0 57868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1649977179
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_32
timestamp 1649977179
transform 1 0 4048 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_38
timestamp 1649977179
transform 1 0 4600 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_41
timestamp 1649977179
transform 1 0 4876 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1649977179
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_73
timestamp 1649977179
transform 1 0 7820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_85
timestamp 1649977179
transform 1 0 8924 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_96
timestamp 1649977179
transform 1 0 9936 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_104
timestamp 1649977179
transform 1 0 10672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_108
timestamp 1649977179
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_117
timestamp 1649977179
transform 1 0 11868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_128
timestamp 1649977179
transform 1 0 12880 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1649977179
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_151
timestamp 1649977179
transform 1 0 14996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1649977179
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_175
timestamp 1649977179
transform 1 0 17204 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_183
timestamp 1649977179
transform 1 0 17940 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_201
timestamp 1649977179
transform 1 0 19596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_213
timestamp 1649977179
transform 1 0 20700 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1649977179
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_233
timestamp 1649977179
transform 1 0 22540 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_239
timestamp 1649977179
transform 1 0 23092 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_248
timestamp 1649977179
transform 1 0 23920 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_257
timestamp 1649977179
transform 1 0 24748 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_265
timestamp 1649977179
transform 1 0 25484 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_271
timestamp 1649977179
transform 1 0 26036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_285
timestamp 1649977179
transform 1 0 27324 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_302
timestamp 1649977179
transform 1 0 28888 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_318
timestamp 1649977179
transform 1 0 30360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_324
timestamp 1649977179
transform 1 0 30912 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_330
timestamp 1649977179
transform 1 0 31464 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1649977179
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_401
timestamp 1649977179
transform 1 0 37996 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_407
timestamp 1649977179
transform 1 0 38548 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_424
timestamp 1649977179
transform 1 0 40112 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_444
timestamp 1649977179
transform 1 0 41952 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1649977179
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_37
timestamp 1649977179
transform 1 0 4508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_45
timestamp 1649977179
transform 1 0 5244 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_48
timestamp 1649977179
transform 1 0 5520 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_57
timestamp 1649977179
transform 1 0 6348 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_69
timestamp 1649977179
transform 1 0 7452 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1649977179
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_103
timestamp 1649977179
transform 1 0 10580 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_108
timestamp 1649977179
transform 1 0 11040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_118
timestamp 1649977179
transform 1 0 11960 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_126
timestamp 1649977179
transform 1 0 12696 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_130
timestamp 1649977179
transform 1 0 13064 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1649977179
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_151
timestamp 1649977179
transform 1 0 14996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_167
timestamp 1649977179
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1649977179
transform 1 0 17204 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_179
timestamp 1649977179
transform 1 0 17572 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_190
timestamp 1649977179
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_205
timestamp 1649977179
transform 1 0 19964 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_211
timestamp 1649977179
transform 1 0 20516 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_219
timestamp 1649977179
transform 1 0 21252 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_241
timestamp 1649977179
transform 1 0 23276 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1649977179
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1649977179
transform 1 0 24840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_264
timestamp 1649977179
transform 1 0 25392 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_268
timestamp 1649977179
transform 1 0 25760 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_274
timestamp 1649977179
transform 1 0 26312 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_286
timestamp 1649977179
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_298
timestamp 1649977179
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1649977179
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_311
timestamp 1649977179
transform 1 0 29716 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_317
timestamp 1649977179
transform 1 0 30268 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_338
timestamp 1649977179
transform 1 0 32200 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_344
timestamp 1649977179
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1649977179
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_383
timestamp 1649977179
transform 1 0 36340 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_400
timestamp 1649977179
transform 1 0 37904 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_409
timestamp 1649977179
transform 1 0 38732 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_417
timestamp 1649977179
transform 1 0 39468 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1649977179
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1649977179
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1649977179
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1649977179
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1649977179
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_18
timestamp 1649977179
transform 1 0 2760 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_30
timestamp 1649977179
transform 1 0 3864 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_36
timestamp 1649977179
transform 1 0 4416 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1649977179
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_97
timestamp 1649977179
transform 1 0 10028 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1649977179
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_126
timestamp 1649977179
transform 1 0 12696 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1649977179
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_154
timestamp 1649977179
transform 1 0 15272 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_157
timestamp 1649977179
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1649977179
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1649977179
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_183
timestamp 1649977179
transform 1 0 17940 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_191
timestamp 1649977179
transform 1 0 18676 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_199
timestamp 1649977179
transform 1 0 19412 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_213
timestamp 1649977179
transform 1 0 20700 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_221
timestamp 1649977179
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_243
timestamp 1649977179
transform 1 0 23460 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_259
timestamp 1649977179
transform 1 0 24932 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1649977179
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_283
timestamp 1649977179
transform 1 0 27140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_297
timestamp 1649977179
transform 1 0 28428 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_303
timestamp 1649977179
transform 1 0 28980 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_323
timestamp 1649977179
transform 1 0 30820 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_343
timestamp 1649977179
transform 1 0 32660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_347
timestamp 1649977179
transform 1 0 33028 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_364
timestamp 1649977179
transform 1 0 34592 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_370
timestamp 1649977179
transform 1 0 35144 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_382
timestamp 1649977179
transform 1 0 36248 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1649977179
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1649977179
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1649977179
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1649977179
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1649977179
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1649977179
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_34
timestamp 1649977179
transform 1 0 4232 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_38
timestamp 1649977179
transform 1 0 4600 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_47
timestamp 1649977179
transform 1 0 5428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_55
timestamp 1649977179
transform 1 0 6164 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_59
timestamp 1649977179
transform 1 0 6532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_71
timestamp 1649977179
transform 1 0 7636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_93
timestamp 1649977179
transform 1 0 9660 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_103
timestamp 1649977179
transform 1 0 10580 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_131
timestamp 1649977179
transform 1 0 13156 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_147
timestamp 1649977179
transform 1 0 14628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_158
timestamp 1649977179
transform 1 0 15640 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_166
timestamp 1649977179
transform 1 0 16376 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_174
timestamp 1649977179
transform 1 0 17112 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1649977179
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1649977179
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_199
timestamp 1649977179
transform 1 0 19412 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_211
timestamp 1649977179
transform 1 0 20516 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_217
timestamp 1649977179
transform 1 0 21068 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_226
timestamp 1649977179
transform 1 0 21896 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_248
timestamp 1649977179
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_255
timestamp 1649977179
transform 1 0 24564 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_275
timestamp 1649977179
transform 1 0 26404 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_295
timestamp 1649977179
transform 1 0 28244 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_303
timestamp 1649977179
transform 1 0 28980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_325
timestamp 1649977179
transform 1 0 31004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_339
timestamp 1649977179
transform 1 0 32292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_351
timestamp 1649977179
transform 1 0 33396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1649977179
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_373
timestamp 1649977179
transform 1 0 35420 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_385
timestamp 1649977179
transform 1 0 36524 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_409
timestamp 1649977179
transform 1 0 38732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1649977179
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_11
timestamp 1649977179
transform 1 0 2116 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_29
timestamp 1649977179
transform 1 0 3772 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_35
timestamp 1649977179
transform 1 0 4324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_47
timestamp 1649977179
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_61
timestamp 1649977179
transform 1 0 6716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_78
timestamp 1649977179
transform 1 0 8280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_90
timestamp 1649977179
transform 1 0 9384 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_96
timestamp 1649977179
transform 1 0 9936 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1649977179
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_121
timestamp 1649977179
transform 1 0 12236 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_130
timestamp 1649977179
transform 1 0 13064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_143
timestamp 1649977179
transform 1 0 14260 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_157
timestamp 1649977179
transform 1 0 15548 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1649977179
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_173
timestamp 1649977179
transform 1 0 17020 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_179
timestamp 1649977179
transform 1 0 17572 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_182
timestamp 1649977179
transform 1 0 17848 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1649977179
transform 1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_198
timestamp 1649977179
transform 1 0 19320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_201
timestamp 1649977179
transform 1 0 19596 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_209
timestamp 1649977179
transform 1 0 20332 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1649977179
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_228
timestamp 1649977179
transform 1 0 22080 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_240
timestamp 1649977179
transform 1 0 23184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_243
timestamp 1649977179
transform 1 0 23460 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_251
timestamp 1649977179
transform 1 0 24196 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_263
timestamp 1649977179
transform 1 0 25300 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1649977179
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_299
timestamp 1649977179
transform 1 0 28612 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_302
timestamp 1649977179
transform 1 0 28888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_316
timestamp 1649977179
transform 1 0 30176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1649977179
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_347
timestamp 1649977179
transform 1 0 33028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_358
timestamp 1649977179
transform 1 0 34040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_362
timestamp 1649977179
transform 1 0 34408 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_368
timestamp 1649977179
transform 1 0 34960 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_380
timestamp 1649977179
transform 1 0 36064 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_407
timestamp 1649977179
transform 1 0 38548 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_431
timestamp 1649977179
transform 1 0 40756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_443
timestamp 1649977179
transform 1 0 41860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_621
timestamp 1649977179
transform 1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_23
timestamp 1649977179
transform 1 0 3220 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_37
timestamp 1649977179
transform 1 0 4508 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_46
timestamp 1649977179
transform 1 0 5336 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_58
timestamp 1649977179
transform 1 0 6440 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_64
timestamp 1649977179
transform 1 0 6992 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_70
timestamp 1649977179
transform 1 0 7544 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1649977179
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_90
timestamp 1649977179
transform 1 0 9384 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_99
timestamp 1649977179
transform 1 0 10212 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_111
timestamp 1649977179
transform 1 0 11316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_122
timestamp 1649977179
transform 1 0 12328 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_128
timestamp 1649977179
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_146
timestamp 1649977179
transform 1 0 14536 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_152
timestamp 1649977179
transform 1 0 15088 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_169
timestamp 1649977179
transform 1 0 16652 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_181
timestamp 1649977179
transform 1 0 17756 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_190
timestamp 1649977179
transform 1 0 18584 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_205
timestamp 1649977179
transform 1 0 19964 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_211
timestamp 1649977179
transform 1 0 20516 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_219
timestamp 1649977179
transform 1 0 21252 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_224
timestamp 1649977179
transform 1 0 21712 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_234
timestamp 1649977179
transform 1 0 22632 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_242
timestamp 1649977179
transform 1 0 23368 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1649977179
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_261
timestamp 1649977179
transform 1 0 25116 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_267
timestamp 1649977179
transform 1 0 25668 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_279
timestamp 1649977179
transform 1 0 26772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_291
timestamp 1649977179
transform 1 0 27876 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_299
timestamp 1649977179
transform 1 0 28612 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_316
timestamp 1649977179
transform 1 0 30176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_320
timestamp 1649977179
transform 1 0 30544 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_323
timestamp 1649977179
transform 1 0 30820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_347
timestamp 1649977179
transform 1 0 33028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1649977179
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_371
timestamp 1649977179
transform 1 0 35236 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_92
timestamp 1649977179
transform 1 0 9568 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1649977179
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_124
timestamp 1649977179
transform 1 0 12512 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_136
timestamp 1649977179
transform 1 0 13616 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1649977179
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_152
timestamp 1649977179
transform 1 0 15088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1649977179
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_177
timestamp 1649977179
transform 1 0 17388 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_197
timestamp 1649977179
transform 1 0 19228 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_206
timestamp 1649977179
transform 1 0 20056 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_262
timestamp 1649977179
transform 1 0 25208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1649977179
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1649977179
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_311
timestamp 1649977179
transform 1 0 29716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_315
timestamp 1649977179
transform 1 0 30084 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_321
timestamp 1649977179
transform 1 0 30636 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_333
timestamp 1649977179
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_360
timestamp 1649977179
transform 1 0 34224 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_366
timestamp 1649977179
transform 1 0 34776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_369
timestamp 1649977179
transform 1 0 35052 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_381
timestamp 1649977179
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1649977179
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_409
timestamp 1649977179
transform 1 0 38732 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_421
timestamp 1649977179
transform 1 0 39836 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_433
timestamp 1649977179
transform 1 0 40940 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_445
timestamp 1649977179
transform 1 0 42044 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1649977179
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_39
timestamp 1649977179
transform 1 0 4692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_51
timestamp 1649977179
transform 1 0 5796 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_64
timestamp 1649977179
transform 1 0 6992 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_71
timestamp 1649977179
transform 1 0 7636 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_104
timestamp 1649977179
transform 1 0 10672 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_118
timestamp 1649977179
transform 1 0 11960 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_122
timestamp 1649977179
transform 1 0 12328 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_130
timestamp 1649977179
transform 1 0 13064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_136
timestamp 1649977179
transform 1 0 13616 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_164
timestamp 1649977179
transform 1 0 16192 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_170
timestamp 1649977179
transform 1 0 16744 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_182
timestamp 1649977179
transform 1 0 17848 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1649977179
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_205
timestamp 1649977179
transform 1 0 19964 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_213
timestamp 1649977179
transform 1 0 20700 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_225
timestamp 1649977179
transform 1 0 21804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_228
timestamp 1649977179
transform 1 0 22080 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_234
timestamp 1649977179
transform 1 0 22632 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_239
timestamp 1649977179
transform 1 0 23092 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1649977179
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_285
timestamp 1649977179
transform 1 0 27324 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_297
timestamp 1649977179
transform 1 0 28428 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1649977179
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_311
timestamp 1649977179
transform 1 0 29716 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_317
timestamp 1649977179
transform 1 0 30268 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_320
timestamp 1649977179
transform 1 0 30544 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_328
timestamp 1649977179
transform 1 0 31280 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_347
timestamp 1649977179
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1649977179
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_370
timestamp 1649977179
transform 1 0 35144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_382
timestamp 1649977179
transform 1 0 36248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_390
timestamp 1649977179
transform 1 0 36984 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_409
timestamp 1649977179
transform 1 0 38732 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_417
timestamp 1649977179
transform 1 0 39468 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_617
timestamp 1649977179
transform 1 0 57868 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_621
timestamp 1649977179
transform 1 0 58236 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_25
timestamp 1649977179
transform 1 0 3404 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_31
timestamp 1649977179
transform 1 0 3956 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_45
timestamp 1649977179
transform 1 0 5244 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_49
timestamp 1649977179
transform 1 0 5612 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_52
timestamp 1649977179
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_65
timestamp 1649977179
transform 1 0 7084 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_71
timestamp 1649977179
transform 1 0 7636 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_83
timestamp 1649977179
transform 1 0 8740 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_89
timestamp 1649977179
transform 1 0 9292 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_101
timestamp 1649977179
transform 1 0 10396 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_107
timestamp 1649977179
transform 1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_117
timestamp 1649977179
transform 1 0 11868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_123
timestamp 1649977179
transform 1 0 12420 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_130
timestamp 1649977179
transform 1 0 13064 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_134
timestamp 1649977179
transform 1 0 13432 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_143
timestamp 1649977179
transform 1 0 14260 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_157
timestamp 1649977179
transform 1 0 15548 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1649977179
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_175
timestamp 1649977179
transform 1 0 17204 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_187
timestamp 1649977179
transform 1 0 18308 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_196
timestamp 1649977179
transform 1 0 19136 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_235
timestamp 1649977179
transform 1 0 22724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_247
timestamp 1649977179
transform 1 0 23828 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_255
timestamp 1649977179
transform 1 0 24564 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_266
timestamp 1649977179
transform 1 0 25576 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1649977179
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_303
timestamp 1649977179
transform 1 0 28980 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_316
timestamp 1649977179
transform 1 0 30176 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_323
timestamp 1649977179
transform 1 0 30820 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1649977179
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_347
timestamp 1649977179
transform 1 0 33028 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_355
timestamp 1649977179
transform 1 0 33764 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_367
timestamp 1649977179
transform 1 0 34868 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_381
timestamp 1649977179
transform 1 0 36156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_389
timestamp 1649977179
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_398
timestamp 1649977179
transform 1 0 37720 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_410
timestamp 1649977179
transform 1 0 38824 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_422
timestamp 1649977179
transform 1 0 39928 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_434
timestamp 1649977179
transform 1 0 41032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1649977179
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_24
timestamp 1649977179
transform 1 0 3312 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_34
timestamp 1649977179
transform 1 0 4232 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_46
timestamp 1649977179
transform 1 0 5336 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_54
timestamp 1649977179
transform 1 0 6072 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_71
timestamp 1649977179
transform 1 0 7636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_96
timestamp 1649977179
transform 1 0 9936 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_100
timestamp 1649977179
transform 1 0 10304 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_127
timestamp 1649977179
transform 1 0 12788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_136
timestamp 1649977179
transform 1 0 13616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_157
timestamp 1649977179
transform 1 0 15548 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_161
timestamp 1649977179
transform 1 0 15916 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_182
timestamp 1649977179
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1649977179
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_213
timestamp 1649977179
transform 1 0 20700 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_224
timestamp 1649977179
transform 1 0 21712 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_238
timestamp 1649977179
transform 1 0 23000 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_244
timestamp 1649977179
transform 1 0 23552 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1649977179
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_262
timestamp 1649977179
transform 1 0 25208 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_282
timestamp 1649977179
transform 1 0 27048 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_294
timestamp 1649977179
transform 1 0 28152 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1649977179
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_317
timestamp 1649977179
transform 1 0 30268 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_347
timestamp 1649977179
transform 1 0 33028 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1649977179
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_368
timestamp 1649977179
transform 1 0 34960 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_392
timestamp 1649977179
transform 1 0 37168 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_404
timestamp 1649977179
transform 1 0 38272 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1649977179
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_617
timestamp 1649977179
transform 1 0 57868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_621
timestamp 1649977179
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1649977179
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1649977179
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1649977179
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_73
timestamp 1649977179
transform 1 0 7820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_85
timestamp 1649977179
transform 1 0 8924 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_101
timestamp 1649977179
transform 1 0 10396 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1649977179
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_123
timestamp 1649977179
transform 1 0 12420 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_129
timestamp 1649977179
transform 1 0 12972 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_133
timestamp 1649977179
transform 1 0 13340 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1649977179
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_142
timestamp 1649977179
transform 1 0 14168 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_154
timestamp 1649977179
transform 1 0 15272 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1649977179
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_177
timestamp 1649977179
transform 1 0 17388 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_183
timestamp 1649977179
transform 1 0 17940 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_195
timestamp 1649977179
transform 1 0 19044 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_200
timestamp 1649977179
transform 1 0 19504 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_214
timestamp 1649977179
transform 1 0 20792 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1649977179
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_229
timestamp 1649977179
transform 1 0 22172 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_239
timestamp 1649977179
transform 1 0 23092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_245
timestamp 1649977179
transform 1 0 23644 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1649977179
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_262
timestamp 1649977179
transform 1 0 25208 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_270
timestamp 1649977179
transform 1 0 25944 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_304
timestamp 1649977179
transform 1 0 29072 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_310
timestamp 1649977179
transform 1 0 29624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_313
timestamp 1649977179
transform 1 0 29900 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_323
timestamp 1649977179
transform 1 0 30820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_346
timestamp 1649977179
transform 1 0 32936 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_358
timestamp 1649977179
transform 1 0 34040 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_370
timestamp 1649977179
transform 1 0 35144 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1649977179
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1649977179
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_7
timestamp 1649977179
transform 1 0 1748 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1649977179
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_49
timestamp 1649977179
transform 1 0 5612 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_70
timestamp 1649977179
transform 1 0 7544 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_76
timestamp 1649977179
transform 1 0 8096 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_101
timestamp 1649977179
transform 1 0 10396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_113
timestamp 1649977179
transform 1 0 11500 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_132
timestamp 1649977179
transform 1 0 13248 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_143
timestamp 1649977179
transform 1 0 14260 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_155
timestamp 1649977179
transform 1 0 15364 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_179
timestamp 1649977179
transform 1 0 17572 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1649977179
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_206
timestamp 1649977179
transform 1 0 20056 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_212
timestamp 1649977179
transform 1 0 20608 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_224
timestamp 1649977179
transform 1 0 21712 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_232
timestamp 1649977179
transform 1 0 22448 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_237
timestamp 1649977179
transform 1 0 22908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1649977179
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_269
timestamp 1649977179
transform 1 0 25852 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_291
timestamp 1649977179
transform 1 0 27876 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1649977179
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_317
timestamp 1649977179
transform 1 0 30268 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_325
timestamp 1649977179
transform 1 0 31004 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_334
timestamp 1649977179
transform 1 0 31832 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_373
timestamp 1649977179
transform 1 0 35420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_380
timestamp 1649977179
transform 1 0 36064 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_388
timestamp 1649977179
transform 1 0 36800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_406
timestamp 1649977179
transform 1 0 38456 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1649977179
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_31
timestamp 1649977179
transform 1 0 3956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_47
timestamp 1649977179
transform 1 0 5428 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1649977179
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_65
timestamp 1649977179
transform 1 0 7084 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_71
timestamp 1649977179
transform 1 0 7636 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_87
timestamp 1649977179
transform 1 0 9108 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_99
timestamp 1649977179
transform 1 0 10212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_130
timestamp 1649977179
transform 1 0 13064 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_138
timestamp 1649977179
transform 1 0 13800 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_147
timestamp 1649977179
transform 1 0 14628 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_156
timestamp 1649977179
transform 1 0 15456 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_177
timestamp 1649977179
transform 1 0 17388 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_189
timestamp 1649977179
transform 1 0 18492 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_201
timestamp 1649977179
transform 1 0 19596 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_213
timestamp 1649977179
transform 1 0 20700 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1649977179
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_233
timestamp 1649977179
transform 1 0 22540 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_241
timestamp 1649977179
transform 1 0 23276 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_258
timestamp 1649977179
transform 1 0 24840 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_264
timestamp 1649977179
transform 1 0 25392 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1649977179
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_325
timestamp 1649977179
transform 1 0 31004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1649977179
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_347
timestamp 1649977179
transform 1 0 33028 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_359
timestamp 1649977179
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_382
timestamp 1649977179
transform 1 0 36248 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1649977179
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_621
timestamp 1649977179
transform 1 0 58236 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_37
timestamp 1649977179
transform 1 0 4508 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_43
timestamp 1649977179
transform 1 0 5060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_55
timestamp 1649977179
transform 1 0 6164 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_62
timestamp 1649977179
transform 1 0 6808 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_69
timestamp 1649977179
transform 1 0 7452 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_75
timestamp 1649977179
transform 1 0 8004 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1649977179
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1649977179
transform 1 0 9476 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_102
timestamp 1649977179
transform 1 0 10488 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_114
timestamp 1649977179
transform 1 0 11592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_122
timestamp 1649977179
transform 1 0 12328 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_131
timestamp 1649977179
transform 1 0 13156 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_157
timestamp 1649977179
transform 1 0 15548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_169
timestamp 1649977179
transform 1 0 16652 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_182
timestamp 1649977179
transform 1 0 17848 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1649977179
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_205
timestamp 1649977179
transform 1 0 19964 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_224
timestamp 1649977179
transform 1 0 21712 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_232
timestamp 1649977179
transform 1 0 22448 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_235
timestamp 1649977179
transform 1 0 22724 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_243
timestamp 1649977179
transform 1 0 23460 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1649977179
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_263
timestamp 1649977179
transform 1 0 25300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_275
timestamp 1649977179
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_287
timestamp 1649977179
transform 1 0 27508 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_295
timestamp 1649977179
transform 1 0 28244 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1649977179
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_311
timestamp 1649977179
transform 1 0 29716 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_323
timestamp 1649977179
transform 1 0 30820 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_327
timestamp 1649977179
transform 1 0 31188 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_339
timestamp 1649977179
transform 1 0 32292 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_348
timestamp 1649977179
transform 1 0 33120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1649977179
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_374
timestamp 1649977179
transform 1 0 35512 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_386
timestamp 1649977179
transform 1 0 36616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_390
timestamp 1649977179
transform 1 0 36984 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_407
timestamp 1649977179
transform 1 0 38548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_36
timestamp 1649977179
transform 1 0 4416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1649977179
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1649977179
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_57_79
timestamp 1649977179
transform 1 0 8372 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_90
timestamp 1649977179
transform 1 0 9384 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_98
timestamp 1649977179
transform 1 0 10120 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_106
timestamp 1649977179
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_143
timestamp 1649977179
transform 1 0 14260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_151
timestamp 1649977179
transform 1 0 14996 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_158
timestamp 1649977179
transform 1 0 15640 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1649977179
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_177
timestamp 1649977179
transform 1 0 17388 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_189
timestamp 1649977179
transform 1 0 18492 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_203
timestamp 1649977179
transform 1 0 19780 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_209
timestamp 1649977179
transform 1 0 20332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1649977179
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_227
timestamp 1649977179
transform 1 0 21988 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_235
timestamp 1649977179
transform 1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_239
timestamp 1649977179
transform 1 0 23092 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_245
timestamp 1649977179
transform 1 0 23644 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_257
timestamp 1649977179
transform 1 0 24748 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_263
timestamp 1649977179
transform 1 0 25300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1649977179
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_301
timestamp 1649977179
transform 1 0 28796 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_306
timestamp 1649977179
transform 1 0 29256 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_318
timestamp 1649977179
transform 1 0 30360 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1649977179
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_369
timestamp 1649977179
transform 1 0 35052 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_409
timestamp 1649977179
transform 1 0 38732 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_421
timestamp 1649977179
transform 1 0 39836 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_433
timestamp 1649977179
transform 1 0 40940 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_445
timestamp 1649977179
transform 1 0 42044 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1649977179
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_21
timestamp 1649977179
transform 1 0 3036 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1649977179
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_37
timestamp 1649977179
transform 1 0 4508 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_45
timestamp 1649977179
transform 1 0 5244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_57
timestamp 1649977179
transform 1 0 6348 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_93
timestamp 1649977179
transform 1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_101
timestamp 1649977179
transform 1 0 10396 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_110
timestamp 1649977179
transform 1 0 11224 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_116
timestamp 1649977179
transform 1 0 11776 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_128
timestamp 1649977179
transform 1 0 12880 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_136
timestamp 1649977179
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_151
timestamp 1649977179
transform 1 0 14996 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_159
timestamp 1649977179
transform 1 0 15732 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_166
timestamp 1649977179
transform 1 0 16376 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_174
timestamp 1649977179
transform 1 0 17112 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_184
timestamp 1649977179
transform 1 0 18032 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_214
timestamp 1649977179
transform 1 0 20792 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_226
timestamp 1649977179
transform 1 0 21896 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_230
timestamp 1649977179
transform 1 0 22264 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_236
timestamp 1649977179
transform 1 0 22816 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1649977179
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_256
timestamp 1649977179
transform 1 0 24656 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_268
timestamp 1649977179
transform 1 0 25760 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_288
timestamp 1649977179
transform 1 0 27600 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_300
timestamp 1649977179
transform 1 0 28704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_342
timestamp 1649977179
transform 1 0 32568 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_350
timestamp 1649977179
transform 1 0 33304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_353
timestamp 1649977179
transform 1 0 33580 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_361
timestamp 1649977179
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_371
timestamp 1649977179
transform 1 0 35236 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_374
timestamp 1649977179
transform 1 0 35512 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_386
timestamp 1649977179
transform 1 0 36616 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_398
timestamp 1649977179
transform 1 0 37720 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_410
timestamp 1649977179
transform 1 0 38824 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_418
timestamp 1649977179
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_31
timestamp 1649977179
transform 1 0 3956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_43
timestamp 1649977179
transform 1 0 5060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1649977179
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_59
timestamp 1649977179
transform 1 0 6532 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_65
timestamp 1649977179
transform 1 0 7084 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_82
timestamp 1649977179
transform 1 0 8648 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_104
timestamp 1649977179
transform 1 0 10672 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_119
timestamp 1649977179
transform 1 0 12052 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_127
timestamp 1649977179
transform 1 0 12788 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_139
timestamp 1649977179
transform 1 0 13892 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_151
timestamp 1649977179
transform 1 0 14996 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_163
timestamp 1649977179
transform 1 0 16100 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_185
timestamp 1649977179
transform 1 0 18124 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_201
timestamp 1649977179
transform 1 0 19596 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_208
timestamp 1649977179
transform 1 0 20240 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1649977179
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_254
timestamp 1649977179
transform 1 0 24472 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_263
timestamp 1649977179
transform 1 0 25300 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_275
timestamp 1649977179
transform 1 0 26404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_284
timestamp 1649977179
transform 1 0 27232 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_297
timestamp 1649977179
transform 1 0 28428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_307
timestamp 1649977179
transform 1 0 29348 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_313
timestamp 1649977179
transform 1 0 29900 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_327
timestamp 1649977179
transform 1 0 31188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_345
timestamp 1649977179
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_33
timestamp 1649977179
transform 1 0 4140 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_39
timestamp 1649977179
transform 1 0 4692 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_45
timestamp 1649977179
transform 1 0 5244 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_58
timestamp 1649977179
transform 1 0 6440 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_66
timestamp 1649977179
transform 1 0 7176 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_72
timestamp 1649977179
transform 1 0 7728 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_101
timestamp 1649977179
transform 1 0 10396 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_118
timestamp 1649977179
transform 1 0 11960 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_129
timestamp 1649977179
transform 1 0 12972 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_137
timestamp 1649977179
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_176
timestamp 1649977179
transform 1 0 17296 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_185
timestamp 1649977179
transform 1 0 18124 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_193
timestamp 1649977179
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_201
timestamp 1649977179
transform 1 0 19596 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_207
timestamp 1649977179
transform 1 0 20148 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_228
timestamp 1649977179
transform 1 0 22080 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1649977179
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_282
timestamp 1649977179
transform 1 0 27048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_294
timestamp 1649977179
transform 1 0 28152 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 1649977179
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_320
timestamp 1649977179
transform 1 0 30544 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_340
timestamp 1649977179
transform 1 0 32384 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_348
timestamp 1649977179
transform 1 0 33120 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_359
timestamp 1649977179
transform 1 0 34132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_617
timestamp 1649977179
transform 1 0 57868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1649977179
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_34
timestamp 1649977179
transform 1 0 4232 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_46
timestamp 1649977179
transform 1 0 5336 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1649977179
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_59
timestamp 1649977179
transform 1 0 6532 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_71
timestamp 1649977179
transform 1 0 7636 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_83
timestamp 1649977179
transform 1 0 8740 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_95
timestamp 1649977179
transform 1 0 9844 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_106
timestamp 1649977179
transform 1 0 10856 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_119
timestamp 1649977179
transform 1 0 12052 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_131
timestamp 1649977179
transform 1 0 13156 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_172
timestamp 1649977179
transform 1 0 16928 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_178
timestamp 1649977179
transform 1 0 17480 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_190
timestamp 1649977179
transform 1 0 18584 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_198
timestamp 1649977179
transform 1 0 19320 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_203
timestamp 1649977179
transform 1 0 19780 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_215
timestamp 1649977179
transform 1 0 20884 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_230
timestamp 1649977179
transform 1 0 22264 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_242
timestamp 1649977179
transform 1 0 23368 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_248
timestamp 1649977179
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_254
timestamp 1649977179
transform 1 0 24472 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_266
timestamp 1649977179
transform 1 0 25576 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_278
timestamp 1649977179
transform 1 0 26680 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_301
timestamp 1649977179
transform 1 0 28796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_310
timestamp 1649977179
transform 1 0 29624 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_318
timestamp 1649977179
transform 1 0 30360 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_346
timestamp 1649977179
transform 1 0 32936 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_366
timestamp 1649977179
transform 1 0 34776 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_386
timestamp 1649977179
transform 1 0 36616 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_70
timestamp 1649977179
transform 1 0 7544 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_79
timestamp 1649977179
transform 1 0 8372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_106
timestamp 1649977179
transform 1 0 10856 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_112
timestamp 1649977179
transform 1 0 11408 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 1649977179
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_149
timestamp 1649977179
transform 1 0 14812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_155
timestamp 1649977179
transform 1 0 15364 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_161
timestamp 1649977179
transform 1 0 15916 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_170
timestamp 1649977179
transform 1 0 16744 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_181
timestamp 1649977179
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_193
timestamp 1649977179
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_213
timestamp 1649977179
transform 1 0 20700 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_216
timestamp 1649977179
transform 1 0 20976 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_228
timestamp 1649977179
transform 1 0 22080 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_232
timestamp 1649977179
transform 1 0 22448 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_235
timestamp 1649977179
transform 1 0 22724 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_246
timestamp 1649977179
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_258
timestamp 1649977179
transform 1 0 24840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_270
timestamp 1649977179
transform 1 0 25944 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_278
timestamp 1649977179
transform 1 0 26680 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_284
timestamp 1649977179
transform 1 0 27232 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_296
timestamp 1649977179
transform 1 0 28336 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_319
timestamp 1649977179
transform 1 0 30452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_328
timestamp 1649977179
transform 1 0 31280 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_356
timestamp 1649977179
transform 1 0 33856 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_373
timestamp 1649977179
transform 1 0 35420 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_385
timestamp 1649977179
transform 1 0 36524 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_388
timestamp 1649977179
transform 1 0 36800 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_412
timestamp 1649977179
transform 1 0 39008 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_617
timestamp 1649977179
transform 1 0 57868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1649977179
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_24
timestamp 1649977179
transform 1 0 3312 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_36
timestamp 1649977179
transform 1 0 4416 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1649977179
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_60
timestamp 1649977179
transform 1 0 6624 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_72
timestamp 1649977179
transform 1 0 7728 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_84
timestamp 1649977179
transform 1 0 8832 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_101
timestamp 1649977179
transform 1 0 10396 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 1649977179
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_121
timestamp 1649977179
transform 1 0 12236 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_129
timestamp 1649977179
transform 1 0 12972 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_136
timestamp 1649977179
transform 1 0 13616 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_144
timestamp 1649977179
transform 1 0 14352 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_150
timestamp 1649977179
transform 1 0 14904 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_162
timestamp 1649977179
transform 1 0 16008 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_173
timestamp 1649977179
transform 1 0 17020 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_182
timestamp 1649977179
transform 1 0 17848 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_188
timestamp 1649977179
transform 1 0 18400 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_208
timestamp 1649977179
transform 1 0 20240 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1649977179
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_233
timestamp 1649977179
transform 1 0 22540 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_244
timestamp 1649977179
transform 1 0 23552 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_252
timestamp 1649977179
transform 1 0 24288 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_270
timestamp 1649977179
transform 1 0 25944 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1649977179
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_285
timestamp 1649977179
transform 1 0 27324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_297
timestamp 1649977179
transform 1 0 28428 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_303
timestamp 1649977179
transform 1 0 28980 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_315
timestamp 1649977179
transform 1 0 30084 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_327
timestamp 1649977179
transform 1 0 31188 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_356
timestamp 1649977179
transform 1 0 33856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_362
timestamp 1649977179
transform 1 0 34408 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_368
timestamp 1649977179
transform 1 0 34960 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_380
timestamp 1649977179
transform 1 0 36064 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1649977179
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1649977179
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_37
timestamp 1649977179
transform 1 0 4508 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_43
timestamp 1649977179
transform 1 0 5060 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_63
timestamp 1649977179
transform 1 0 6900 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_75
timestamp 1649977179
transform 1 0 8004 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_104
timestamp 1649977179
transform 1 0 10672 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_122
timestamp 1649977179
transform 1 0 12328 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_134
timestamp 1649977179
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_157
timestamp 1649977179
transform 1 0 15548 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_173
timestamp 1649977179
transform 1 0 17020 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_181
timestamp 1649977179
transform 1 0 17756 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1649977179
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1649977179
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_222
timestamp 1649977179
transform 1 0 21528 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_236
timestamp 1649977179
transform 1 0 22816 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1649977179
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_269
timestamp 1649977179
transform 1 0 25852 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_281
timestamp 1649977179
transform 1 0 26956 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_287
timestamp 1649977179
transform 1 0 27508 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1649977179
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_341
timestamp 1649977179
transform 1 0 32476 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_353
timestamp 1649977179
transform 1 0 33580 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1649977179
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_11
timestamp 1649977179
transform 1 0 2116 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_21
timestamp 1649977179
transform 1 0 3036 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_45
timestamp 1649977179
transform 1 0 5244 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_65
timestamp 1649977179
transform 1 0 7084 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_74
timestamp 1649977179
transform 1 0 7912 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_85
timestamp 1649977179
transform 1 0 8924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_97
timestamp 1649977179
transform 1 0 10028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_109
timestamp 1649977179
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_141
timestamp 1649977179
transform 1 0 14076 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_159
timestamp 1649977179
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1649977179
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_197
timestamp 1649977179
transform 1 0 19228 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_209
timestamp 1649977179
transform 1 0 20332 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_215
timestamp 1649977179
transform 1 0 20884 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_245
timestamp 1649977179
transform 1 0 23644 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_251
timestamp 1649977179
transform 1 0 24196 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_271
timestamp 1649977179
transform 1 0 26036 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_315
timestamp 1649977179
transform 1 0 30084 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_345
timestamp 1649977179
transform 1 0 32844 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_351
timestamp 1649977179
transform 1 0 33396 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_360
timestamp 1649977179
transform 1 0 34224 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_369
timestamp 1649977179
transform 1 0 35052 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_381
timestamp 1649977179
transform 1 0 36156 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_389
timestamp 1649977179
transform 1 0 36892 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_621
timestamp 1649977179
transform 1 0 58236 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_23
timestamp 1649977179
transform 1 0 3220 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_45
timestamp 1649977179
transform 1 0 5244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_54
timestamp 1649977179
transform 1 0 6072 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_68
timestamp 1649977179
transform 1 0 7360 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1649977179
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_66_96
timestamp 1649977179
transform 1 0 9936 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_108
timestamp 1649977179
transform 1 0 11040 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_116
timestamp 1649977179
transform 1 0 11776 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_132
timestamp 1649977179
transform 1 0 13248 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_160
timestamp 1649977179
transform 1 0 15824 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_172
timestamp 1649977179
transform 1 0 16928 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_181
timestamp 1649977179
transform 1 0 17756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_193
timestamp 1649977179
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_201
timestamp 1649977179
transform 1 0 19596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_213
timestamp 1649977179
transform 1 0 20700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_225
timestamp 1649977179
transform 1 0 21804 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_231
timestamp 1649977179
transform 1 0 22356 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_237
timestamp 1649977179
transform 1 0 22908 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1649977179
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_255
timestamp 1649977179
transform 1 0 24564 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_267
timestamp 1649977179
transform 1 0 25668 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_279
timestamp 1649977179
transform 1 0 26772 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_315
timestamp 1649977179
transform 1 0 30084 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_327
timestamp 1649977179
transform 1 0 31188 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_336
timestamp 1649977179
transform 1 0 32016 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_351
timestamp 1649977179
transform 1 0 33396 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_360
timestamp 1649977179
transform 1 0 34224 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_381
timestamp 1649977179
transform 1 0 36156 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_393
timestamp 1649977179
transform 1 0 37260 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_405
timestamp 1649977179
transform 1 0 38364 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_417
timestamp 1649977179
transform 1 0 39468 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_23
timestamp 1649977179
transform 1 0 3220 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_26
timestamp 1649977179
transform 1 0 3496 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_38
timestamp 1649977179
transform 1 0 4600 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_43
timestamp 1649977179
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_115
timestamp 1649977179
transform 1 0 11684 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_127
timestamp 1649977179
transform 1 0 12788 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_140
timestamp 1649977179
transform 1 0 13984 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_152
timestamp 1649977179
transform 1 0 15088 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_164
timestamp 1649977179
transform 1 0 16192 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_201
timestamp 1649977179
transform 1 0 19596 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_213
timestamp 1649977179
transform 1 0 20700 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_221
timestamp 1649977179
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_227
timestamp 1649977179
transform 1 0 21988 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_239
timestamp 1649977179
transform 1 0 23092 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_248
timestamp 1649977179
transform 1 0 23920 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_260
timestamp 1649977179
transform 1 0 25024 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_272
timestamp 1649977179
transform 1 0 26128 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_285
timestamp 1649977179
transform 1 0 27324 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_297
timestamp 1649977179
transform 1 0 28428 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_306
timestamp 1649977179
transform 1 0 29256 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_314
timestamp 1649977179
transform 1 0 29992 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1649977179
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_345
timestamp 1649977179
transform 1 0 32844 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_359
timestamp 1649977179
transform 1 0 34132 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_379
timestamp 1649977179
transform 1 0 35972 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_621
timestamp 1649977179
transform 1 0 58236 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1649977179
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_34
timestamp 1649977179
transform 1 0 4232 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_58
timestamp 1649977179
transform 1 0 6440 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_70
timestamp 1649977179
transform 1 0 7544 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_82
timestamp 1649977179
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_96
timestamp 1649977179
transform 1 0 9936 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_105
timestamp 1649977179
transform 1 0 10764 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_111
timestamp 1649977179
transform 1 0 11316 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_123
timestamp 1649977179
transform 1 0 12420 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_135
timestamp 1649977179
transform 1 0 13524 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1649977179
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_207
timestamp 1649977179
transform 1 0 20148 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_213
timestamp 1649977179
transform 1 0 20700 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_229
timestamp 1649977179
transform 1 0 22172 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_241
timestamp 1649977179
transform 1 0 23276 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1649977179
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_299
timestamp 1649977179
transform 1 0 28612 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_314
timestamp 1649977179
transform 1 0 29992 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_320
timestamp 1649977179
transform 1 0 30544 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_68_330
timestamp 1649977179
transform 1 0 31464 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_350
timestamp 1649977179
transform 1 0 33304 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_356
timestamp 1649977179
transform 1 0 33856 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_41
timestamp 1649977179
transform 1 0 4876 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1649977179
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_65
timestamp 1649977179
transform 1 0 7084 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_71
timestamp 1649977179
transform 1 0 7636 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_95
timestamp 1649977179
transform 1 0 9844 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_107
timestamp 1649977179
transform 1 0 10948 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_115
timestamp 1649977179
transform 1 0 11684 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_121
timestamp 1649977179
transform 1 0 12236 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_130
timestamp 1649977179
transform 1 0 13064 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_136
timestamp 1649977179
transform 1 0 13616 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_148
timestamp 1649977179
transform 1 0 14720 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_160
timestamp 1649977179
transform 1 0 15824 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_171
timestamp 1649977179
transform 1 0 16836 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_183
timestamp 1649977179
transform 1 0 17940 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_189
timestamp 1649977179
transform 1 0 18492 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_195
timestamp 1649977179
transform 1 0 19044 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_203
timestamp 1649977179
transform 1 0 19780 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1649977179
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_239
timestamp 1649977179
transform 1 0 23092 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_259
timestamp 1649977179
transform 1 0 24932 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_271
timestamp 1649977179
transform 1 0 26036 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_285
timestamp 1649977179
transform 1 0 27324 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_302
timestamp 1649977179
transform 1 0 28888 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_318
timestamp 1649977179
transform 1 0 30360 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_327
timestamp 1649977179
transform 1 0 31188 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_35
timestamp 1649977179
transform 1 0 4324 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_44
timestamp 1649977179
transform 1 0 5152 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_64
timestamp 1649977179
transform 1 0 6992 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_72
timestamp 1649977179
transform 1 0 7728 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_80
timestamp 1649977179
transform 1 0 8464 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_101
timestamp 1649977179
transform 1 0 10396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_129
timestamp 1649977179
transform 1 0 12972 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_137
timestamp 1649977179
transform 1 0 13708 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_149
timestamp 1649977179
transform 1 0 14812 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_166
timestamp 1649977179
transform 1 0 16376 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_190
timestamp 1649977179
transform 1 0 18584 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_213
timestamp 1649977179
transform 1 0 20700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_225
timestamp 1649977179
transform 1 0 21804 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_231
timestamp 1649977179
transform 1 0 22356 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1649977179
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_269
timestamp 1649977179
transform 1 0 25852 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_281
timestamp 1649977179
transform 1 0 26956 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_286
timestamp 1649977179
transform 1 0 27416 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_298
timestamp 1649977179
transform 1 0 28520 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_304
timestamp 1649977179
transform 1 0 29072 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_329
timestamp 1649977179
transform 1 0 31372 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_341
timestamp 1649977179
transform 1 0 32476 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_353
timestamp 1649977179
transform 1 0 33580 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_361
timestamp 1649977179
transform 1 0 34316 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_617
timestamp 1649977179
transform 1 0 57868 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_621
timestamp 1649977179
transform 1 0 58236 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_43
timestamp 1649977179
transform 1 0 5060 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_49
timestamp 1649977179
transform 1 0 5612 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_77
timestamp 1649977179
transform 1 0 8188 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_83
timestamp 1649977179
transform 1 0 8740 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_92
timestamp 1649977179
transform 1 0 9568 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_98
timestamp 1649977179
transform 1 0 10120 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_102
timestamp 1649977179
transform 1 0 10488 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_108
timestamp 1649977179
transform 1 0 11040 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_129
timestamp 1649977179
transform 1 0 12972 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_135
timestamp 1649977179
transform 1 0 13524 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_152
timestamp 1649977179
transform 1 0 15088 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_164
timestamp 1649977179
transform 1 0 16192 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_171
timestamp 1649977179
transform 1 0 16836 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_187
timestamp 1649977179
transform 1 0 18308 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_207
timestamp 1649977179
transform 1 0 20148 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_219
timestamp 1649977179
transform 1 0 21252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_241
timestamp 1649977179
transform 1 0 23276 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_253
timestamp 1649977179
transform 1 0 24380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_265
timestamp 1649977179
transform 1 0 25484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_277
timestamp 1649977179
transform 1 0 26588 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_46
timestamp 1649977179
transform 1 0 5336 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_58
timestamp 1649977179
transform 1 0 6440 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_70
timestamp 1649977179
transform 1 0 7544 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_82
timestamp 1649977179
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_115
timestamp 1649977179
transform 1 0 11684 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_129
timestamp 1649977179
transform 1 0 12972 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_137
timestamp 1649977179
transform 1 0 13708 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_149
timestamp 1649977179
transform 1 0 14812 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_155
timestamp 1649977179
transform 1 0 15364 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_172
timestamp 1649977179
transform 1 0 16928 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_180
timestamp 1649977179
transform 1 0 17664 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_183
timestamp 1649977179
transform 1 0 17940 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_192
timestamp 1649977179
transform 1 0 18768 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_205
timestamp 1649977179
transform 1 0 19964 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_211
timestamp 1649977179
transform 1 0 20516 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_223
timestamp 1649977179
transform 1 0 21620 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_235
timestamp 1649977179
transform 1 0 22724 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_247
timestamp 1649977179
transform 1 0 23828 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_617
timestamp 1649977179
transform 1 0 57868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1649977179
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_119
timestamp 1649977179
transform 1 0 12052 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_131
timestamp 1649977179
transform 1 0 13156 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_143
timestamp 1649977179
transform 1 0 14260 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_152
timestamp 1649977179
transform 1 0 15088 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_164
timestamp 1649977179
transform 1 0 16192 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_171
timestamp 1649977179
transform 1 0 16836 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_183
timestamp 1649977179
transform 1 0 17940 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_73_191
timestamp 1649977179
transform 1 0 18676 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_203
timestamp 1649977179
transform 1 0 19780 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_207
timestamp 1649977179
transform 1 0 20148 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_219
timestamp 1649977179
transform 1 0 21252 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_129
timestamp 1649977179
transform 1 0 12972 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_74_151
timestamp 1649977179
transform 1 0 14996 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_155
timestamp 1649977179
transform 1 0 15364 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_161
timestamp 1649977179
transform 1 0 15916 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_173
timestamp 1649977179
transform 1 0 17020 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_185
timestamp 1649977179
transform 1 0 18124 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_193
timestamp 1649977179
transform 1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_621
timestamp 1649977179
transform 1 0 58236 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_621
timestamp 1649977179
transform 1 0 58236 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_617
timestamp 1649977179
transform 1 0 57868 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_621
timestamp 1649977179
transform 1 0 58236 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_617
timestamp 1649977179
transform 1 0 57868 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_621
timestamp 1649977179
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_621
timestamp 1649977179
transform 1 0 58236 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_621
timestamp 1649977179
transform 1 0 58236 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_617
timestamp 1649977179
transform 1 0 57868 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_621
timestamp 1649977179
transform 1 0 58236 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_617
timestamp 1649977179
transform 1 0 57868 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_621
timestamp 1649977179
transform 1 0 58236 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_621
timestamp 1649977179
transform 1 0 58236 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_621
timestamp 1649977179
transform 1 0 58236 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1649977179
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_621
timestamp 1649977179
transform 1 0 58236 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1649977179
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1649977179
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1649977179
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_301
timestamp 1649977179
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_457
timestamp 1649977179
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_469
timestamp 1649977179
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_475
timestamp 1649977179
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_609
timestamp 1649977179
transform 1 0 57132 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_614
timestamp 1649977179
transform 1 0 57592 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1649977179
transform 1 0 58236 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_7
timestamp 1649977179
transform 1 0 1748 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_11
timestamp 1649977179
transform 1 0 2116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_23
timestamp 1649977179
transform 1 0 3220 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1649977179
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_32
timestamp 1649977179
transform 1 0 4048 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_40
timestamp 1649977179
transform 1 0 4784 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_45
timestamp 1649977179
transform 1 0 5244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1649977179
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_62
timestamp 1649977179
transform 1 0 6808 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_74
timestamp 1649977179
transform 1 0 7912 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_79
timestamp 1649977179
transform 1 0 8372 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_83
timestamp 1649977179
transform 1 0 8740 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_96
timestamp 1649977179
transform 1 0 9936 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_108
timestamp 1649977179
transform 1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_116
timestamp 1649977179
transform 1 0 11776 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_124
timestamp 1649977179
transform 1 0 12512 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_130
timestamp 1649977179
transform 1 0 13064 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_138
timestamp 1649977179
transform 1 0 13800 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_147
timestamp 1649977179
transform 1 0 14628 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_159
timestamp 1649977179
transform 1 0 15732 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_164
timestamp 1649977179
transform 1 0 16192 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_169
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_177
timestamp 1649977179
transform 1 0 17388 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_181
timestamp 1649977179
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_193
timestamp 1649977179
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_200
timestamp 1649977179
transform 1 0 19504 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_215
timestamp 1649977179
transform 1 0 20884 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1649977179
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_232
timestamp 1649977179
transform 1 0 22448 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_244
timestamp 1649977179
transform 1 0 23552 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_101_256
timestamp 1649977179
transform 1 0 24656 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_262
timestamp 1649977179
transform 1 0 25208 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_266
timestamp 1649977179
transform 1 0 25576 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_278
timestamp 1649977179
transform 1 0 26680 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_284
timestamp 1649977179
transform 1 0 27232 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_296
timestamp 1649977179
transform 1 0 28336 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_300
timestamp 1649977179
transform 1 0 28704 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_313
timestamp 1649977179
transform 1 0 29900 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_317
timestamp 1649977179
transform 1 0 30268 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_329
timestamp 1649977179
transform 1 0 31372 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_335
timestamp 1649977179
transform 1 0 31924 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_340
timestamp 1649977179
transform 1 0 32384 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_351
timestamp 1649977179
transform 1 0 33396 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_363
timestamp 1649977179
transform 1 0 34500 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_368
timestamp 1649977179
transform 1 0 34960 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_380
timestamp 1649977179
transform 1 0 36064 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_385
timestamp 1649977179
transform 1 0 36524 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_391
timestamp 1649977179
transform 1 0 37076 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_402
timestamp 1649977179
transform 1 0 38088 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_414
timestamp 1649977179
transform 1 0 39192 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_101_424
timestamp 1649977179
transform 1 0 40112 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_432
timestamp 1649977179
transform 1 0 40848 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_436
timestamp 1649977179
transform 1 0 41216 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_453
timestamp 1649977179
transform 1 0 42780 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_465
timestamp 1649977179
transform 1 0 43884 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_101_470
timestamp 1649977179
transform 1 0 44344 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_477
timestamp 1649977179
transform 1 0 44988 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_483
timestamp 1649977179
transform 1 0 45540 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_487
timestamp 1649977179
transform 1 0 45908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_499
timestamp 1649977179
transform 1 0 47012 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_503
timestamp 1649977179
transform 1 0 47380 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_508
timestamp 1649977179
transform 1 0 47840 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_516
timestamp 1649977179
transform 1 0 48576 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_521
timestamp 1649977179
transform 1 0 49036 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1649977179
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1649977179
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_538
timestamp 1649977179
transform 1 0 50600 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_550
timestamp 1649977179
transform 1 0 51704 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_555
timestamp 1649977179
transform 1 0 52164 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1649977179
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_572
timestamp 1649977179
transform 1 0 53728 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_584
timestamp 1649977179
transform 1 0 54832 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_592
timestamp 1649977179
transform 1 0 55568 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_600
timestamp 1649977179
transform 1 0 56304 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_606
timestamp 1649977179
transform 1 0 56856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1649977179
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1649977179
transform 1 0 58236 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0855_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0856_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0857_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0858_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 1649977179
transform -1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1649977179
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0862_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0863_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14996 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0864_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0865_
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0866_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0867_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4508 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0868_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0869_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0870_
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0871_
timestamp 1649977179
transform -1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1649977179
transform 1 0 4232 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1649977179
transform 1 0 2944 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0874_
timestamp 1649977179
transform 1 0 2116 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 1649977179
transform 1 0 2208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp 1649977179
transform 1 0 3496 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1649977179
transform -1 0 2852 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1649977179
transform -1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1649977179
transform -1 0 8004 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1649977179
transform -1 0 4232 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0888_
timestamp 1649977179
transform -1 0 3312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1649977179
transform -1 0 4692 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 1649977179
transform 1 0 5152 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1649977179
transform -1 0 4508 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0892_
timestamp 1649977179
transform -1 0 3312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0897_
timestamp 1649977179
transform -1 0 12696 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 1649977179
transform -1 0 11868 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1649977179
transform -1 0 12880 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1649977179
transform -1 0 13616 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1649977179
transform -1 0 3128 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1649977179
transform 1 0 2392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0905_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7636 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0909_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0910_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0911_
timestamp 1649977179
transform 1 0 17020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_4  _0912_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11132 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0913_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0914_
timestamp 1649977179
transform 1 0 11408 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0915_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12788 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0916_
timestamp 1649977179
transform -1 0 7360 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1649977179
transform -1 0 12420 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0919_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6072 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1649977179
transform 1 0 3956 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0921_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0922_
timestamp 1649977179
transform -1 0 8556 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1649977179
transform -1 0 3312 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0924_
timestamp 1649977179
transform 1 0 2300 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0925_
timestamp 1649977179
transform -1 0 5888 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 1649977179
transform -1 0 4232 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0927_
timestamp 1649977179
transform 1 0 2576 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0928_
timestamp 1649977179
transform -1 0 7268 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1649977179
transform -1 0 5612 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0930_
timestamp 1649977179
transform -1 0 5152 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0931_
timestamp 1649977179
transform -1 0 7268 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1649977179
transform 1 0 5428 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0933_
timestamp 1649977179
transform -1 0 7084 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0934_
timestamp 1649977179
transform -1 0 26588 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0935_
timestamp 1649977179
transform 1 0 13064 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1649977179
transform -1 0 12236 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1649977179
transform 1 0 13800 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0938_
timestamp 1649977179
transform 1 0 12052 0 1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0939_
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1649977179
transform -1 0 22724 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1649977179
transform 1 0 14628 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0942_
timestamp 1649977179
transform -1 0 16192 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1649977179
transform -1 0 23092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 1649977179
transform 1 0 15456 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1649977179
transform 1 0 15456 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0946_
timestamp 1649977179
transform -1 0 22632 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0947_
timestamp 1649977179
transform 1 0 11224 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0948_
timestamp 1649977179
transform 1 0 12420 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0949_
timestamp 1649977179
transform -1 0 22816 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1649977179
transform -1 0 11040 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1649977179
transform 1 0 12328 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1649977179
transform -1 0 17020 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0953_
timestamp 1649977179
transform 1 0 12696 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1649977179
transform 1 0 12420 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0955_
timestamp 1649977179
transform 1 0 12512 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1649977179
transform -1 0 14996 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1649977179
transform 1 0 13156 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1649977179
transform -1 0 14260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0959_
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1649977179
transform -1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0961_
timestamp 1649977179
transform 1 0 29348 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0962_
timestamp 1649977179
transform 1 0 29808 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0963_
timestamp 1649977179
transform 1 0 30728 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0964_
timestamp 1649977179
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0965_
timestamp 1649977179
transform 1 0 29716 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1649977179
transform -1 0 31188 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1649977179
transform -1 0 28980 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0968_
timestamp 1649977179
transform 1 0 27600 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1649977179
transform -1 0 28428 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0970_
timestamp 1649977179
transform 1 0 27416 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0971_
timestamp 1649977179
transform -1 0 29624 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0972_
timestamp 1649977179
transform 1 0 27692 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1649977179
transform 1 0 32108 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0974_
timestamp 1649977179
transform 1 0 12696 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0975_
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0976_
timestamp 1649977179
transform 1 0 29624 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1649977179
transform -1 0 31280 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1649977179
transform 1 0 29808 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0979_
timestamp 1649977179
transform 1 0 35236 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1649977179
transform -1 0 34960 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0981_
timestamp 1649977179
transform 1 0 35788 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0982_
timestamp 1649977179
transform -1 0 36616 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0983_
timestamp 1649977179
transform 1 0 35604 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0984_
timestamp 1649977179
transform -1 0 36616 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0985_
timestamp 1649977179
transform 1 0 35052 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0986_
timestamp 1649977179
transform -1 0 36524 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0988_
timestamp 1649977179
transform 1 0 28612 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0989_
timestamp 1649977179
transform -1 0 36248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0990_
timestamp 1649977179
transform 1 0 35328 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0991_
timestamp 1649977179
transform -1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0992_
timestamp 1649977179
transform 1 0 34500 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0993_
timestamp 1649977179
transform -1 0 35420 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1649977179
transform -1 0 34224 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0995_
timestamp 1649977179
transform -1 0 33396 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _0996_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0998_
timestamp 1649977179
transform -1 0 30176 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1649977179
transform 1 0 30544 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1000_
timestamp 1649977179
transform -1 0 30452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1649977179
transform 1 0 29716 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1002_
timestamp 1649977179
transform -1 0 31372 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1649977179
transform -1 0 28888 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 1649977179
transform 1 0 28244 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1649977179
transform -1 0 29256 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1006_
timestamp 1649977179
transform -1 0 31372 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1007_
timestamp 1649977179
transform 1 0 27692 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1649977179
transform -1 0 29992 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1649977179
transform 1 0 27784 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1649977179
transform -1 0 31188 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1649977179
transform -1 0 30360 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1649977179
transform 1 0 31556 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1013_
timestamp 1649977179
transform 1 0 30452 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1014_
timestamp 1649977179
transform 1 0 33212 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1649977179
transform -1 0 33212 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1649977179
transform -1 0 32844 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1649977179
transform 1 0 32476 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1019_
timestamp 1649977179
transform 1 0 32476 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1020_
timestamp 1649977179
transform -1 0 35420 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1649977179
transform 1 0 33396 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1649977179
transform -1 0 34316 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1649977179
transform -1 0 34224 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1024_
timestamp 1649977179
transform -1 0 34224 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1649977179
transform 1 0 34592 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1026_
timestamp 1649977179
transform -1 0 34132 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1649977179
transform 1 0 33764 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1028_
timestamp 1649977179
transform -1 0 34868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1029_
timestamp 1649977179
transform -1 0 31648 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1030_
timestamp 1649977179
transform 1 0 29900 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1649977179
transform -1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1032_
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1649977179
transform -1 0 13616 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1034_
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1035_
timestamp 1649977179
transform -1 0 13708 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1036_
timestamp 1649977179
transform -1 0 10120 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1037_
timestamp 1649977179
transform 1 0 14720 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1038_
timestamp 1649977179
transform -1 0 17204 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1649977179
transform 1 0 7176 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1040_
timestamp 1649977179
transform 1 0 6348 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1041_
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1649977179
transform -1 0 5244 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1649977179
transform 1 0 4232 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1649977179
transform 1 0 4324 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1649977179
transform -1 0 4416 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1047_
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1649977179
transform 1 0 7268 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1049_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1050_
timestamp 1649977179
transform 1 0 22448 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1052_
timestamp 1649977179
transform 1 0 7452 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1053_
timestamp 1649977179
transform 1 0 17572 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1054_
timestamp 1649977179
transform -1 0 17848 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 1649977179
transform 1 0 19136 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1056_
timestamp 1649977179
transform -1 0 20148 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1649977179
transform 1 0 18308 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1058_
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1649977179
transform -1 0 19044 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1649977179
transform -1 0 18308 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 1649977179
transform -1 0 20332 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1649977179
transform 1 0 19136 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1064_
timestamp 1649977179
transform -1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1649977179
transform -1 0 19780 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1649977179
transform 1 0 17940 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1649977179
transform 1 0 15732 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1069_
timestamp 1649977179
transform 1 0 15456 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 1649977179
transform -1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1649977179
transform -1 0 18584 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1073_
timestamp 1649977179
transform -1 0 16468 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1074_
timestamp 1649977179
transform 1 0 16928 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1649977179
transform 1 0 16928 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1649977179
transform 1 0 9660 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1077_
timestamp 1649977179
transform 1 0 9568 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1649977179
transform 1 0 9476 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1649977179
transform 1 0 10304 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1649977179
transform 1 0 10948 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1081_
timestamp 1649977179
transform 1 0 23828 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1649977179
transform 1 0 11776 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1649977179
transform -1 0 13708 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1649977179
transform -1 0 15640 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1649977179
transform 1 0 14720 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1649977179
transform 1 0 24656 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1649977179
transform -1 0 23920 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1649977179
transform 1 0 25484 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1090_
timestamp 1649977179
transform -1 0 23920 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1649977179
transform -1 0 24840 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1649977179
transform -1 0 25116 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1093_
timestamp 1649977179
transform -1 0 23644 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1649977179
transform 1 0 24840 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1097_
timestamp 1649977179
transform -1 0 25760 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1649977179
transform -1 0 24656 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1649977179
transform -1 0 24840 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1649977179
transform -1 0 25116 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1649977179
transform -1 0 25208 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1649977179
transform 1 0 24748 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1103_
timestamp 1649977179
transform -1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1104_
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1105_
timestamp 1649977179
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1649977179
transform -1 0 20056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1107_
timestamp 1649977179
transform 1 0 20792 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1109_
timestamp 1649977179
transform 1 0 27600 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1649977179
transform -1 0 24012 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1649977179
transform 1 0 25300 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1113_
timestamp 1649977179
transform 1 0 24380 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1649977179
transform -1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1115_
timestamp 1649977179
transform 1 0 15364 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1649977179
transform -1 0 25944 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1649977179
transform 1 0 23184 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1649977179
transform -1 0 24840 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1120_
timestamp 1649977179
transform 1 0 24288 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1649977179
transform 1 0 27968 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1649977179
transform 1 0 27232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1124_
timestamp 1649977179
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1649977179
transform 1 0 27324 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1126_
timestamp 1649977179
transform -1 0 29072 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1649977179
transform 1 0 30452 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1128_
timestamp 1649977179
transform 1 0 28152 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1129_
timestamp 1649977179
transform 1 0 27600 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1649977179
transform 1 0 31648 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1131_
timestamp 1649977179
transform 1 0 32476 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1649977179
transform 1 0 32752 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1134_
timestamp 1649977179
transform 1 0 30084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1649977179
transform 1 0 31188 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1649977179
transform -1 0 32844 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1137_
timestamp 1649977179
transform 1 0 29992 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1649977179
transform -1 0 31648 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1139_
timestamp 1649977179
transform -1 0 31096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1649977179
transform 1 0 26956 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1649977179
transform 1 0 31556 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1649977179
transform -1 0 32844 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1143_
timestamp 1649977179
transform 1 0 27140 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1145_
timestamp 1649977179
transform 1 0 29440 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1146_
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1649977179
transform -1 0 22816 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1148_
timestamp 1649977179
transform -1 0 25116 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1150_
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1151_
timestamp 1649977179
transform -1 0 24932 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1152_
timestamp 1649977179
transform 1 0 23184 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1649977179
transform -1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1649977179
transform -1 0 19504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1156_
timestamp 1649977179
transform -1 0 19504 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1157_
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1158_
timestamp 1649977179
transform -1 0 20148 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1649977179
transform 1 0 19136 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 1649977179
transform 1 0 13156 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 1649977179
transform 1 0 14168 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1649977179
transform -1 0 15732 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1166_
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1168_
timestamp 1649977179
transform 1 0 25668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1169_
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1170_
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1171_
timestamp 1649977179
transform 1 0 17480 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1172_
timestamp 1649977179
transform 1 0 27508 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1173_
timestamp 1649977179
transform -1 0 27232 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1649977179
transform 1 0 29348 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1175_
timestamp 1649977179
transform -1 0 30544 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1649977179
transform 1 0 29624 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1177_
timestamp 1649977179
transform -1 0 30820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1178_
timestamp 1649977179
transform 1 0 28612 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1179_
timestamp 1649977179
transform -1 0 30360 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1649977179
transform 1 0 27692 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1181_
timestamp 1649977179
transform -1 0 27048 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1649977179
transform 1 0 27600 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1649977179
transform 1 0 27508 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1184_
timestamp 1649977179
transform 1 0 27692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1186_
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1649977179
transform -1 0 20700 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1188_
timestamp 1649977179
transform -1 0 20976 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1189_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1649977179
transform 1 0 23092 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1191_
timestamp 1649977179
transform -1 0 34684 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1192_
timestamp 1649977179
transform 1 0 34868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_
timestamp 1649977179
transform -1 0 38548 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1649977179
transform 1 0 34592 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1195_
timestamp 1649977179
transform -1 0 36340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1649977179
transform -1 0 35328 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1199_
timestamp 1649977179
transform 1 0 36156 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1200_
timestamp 1649977179
transform -1 0 37904 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1649977179
transform 1 0 36984 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1202_
timestamp 1649977179
transform -1 0 37996 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1203_
timestamp 1649977179
transform -1 0 38272 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1204_
timestamp 1649977179
transform -1 0 38180 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1206_
timestamp 1649977179
transform -1 0 39376 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1207_
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1649977179
transform -1 0 37536 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1649977179
transform -1 0 37168 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1210_
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1212_
timestamp 1649977179
transform 1 0 32752 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1213_
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1215_
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1216_
timestamp 1649977179
transform 1 0 38640 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1217_
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1218_
timestamp 1649977179
transform -1 0 41124 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1649977179
transform -1 0 41032 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1649977179
transform 1 0 37628 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_
timestamp 1649977179
transform -1 0 38916 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1649977179
transform 1 0 34960 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1224_
timestamp 1649977179
transform -1 0 35880 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1226_
timestamp 1649977179
transform -1 0 22724 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1227_
timestamp 1649977179
transform 1 0 33304 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1228_
timestamp 1649977179
transform 1 0 35512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1229_
timestamp 1649977179
transform -1 0 37352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1230_
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1231_
timestamp 1649977179
transform -1 0 36616 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1649977179
transform -1 0 35144 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1649977179
transform 1 0 34224 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1649977179
transform -1 0 35144 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1235_
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1236_
timestamp 1649977179
transform 1 0 35604 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1237_
timestamp 1649977179
transform -1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1238_
timestamp 1649977179
transform -1 0 36892 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1649977179
transform -1 0 36800 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1241_
timestamp 1649977179
transform 1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1242_
timestamp 1649977179
transform 1 0 37076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1243_
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1244_
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1649977179
transform 1 0 36432 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1246_
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1247_
timestamp 1649977179
transform 1 0 39008 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1248_
timestamp 1649977179
transform -1 0 38640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1249_
timestamp 1649977179
transform -1 0 38732 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1250_
timestamp 1649977179
transform -1 0 38640 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1251_
timestamp 1649977179
transform 1 0 36340 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1252_
timestamp 1649977179
transform -1 0 38180 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1253_
timestamp 1649977179
transform 1 0 38548 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1254_
timestamp 1649977179
transform -1 0 40204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1255_
timestamp 1649977179
transform 1 0 38640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1649977179
transform 1 0 36800 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1257_
timestamp 1649977179
transform -1 0 38180 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1649977179
transform -1 0 35604 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1649977179
transform -1 0 35512 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1260_
timestamp 1649977179
transform -1 0 22724 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1261_
timestamp 1649977179
transform -1 0 24104 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1262_
timestamp 1649977179
transform -1 0 26680 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1263_
timestamp 1649977179
transform -1 0 27876 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1649977179
transform -1 0 27140 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1649977179
transform -1 0 26496 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1649977179
transform -1 0 25392 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1267_
timestamp 1649977179
transform 1 0 25760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1268_
timestamp 1649977179
transform 1 0 25576 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1269_
timestamp 1649977179
transform 1 0 25760 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1270_
timestamp 1649977179
transform 1 0 25852 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1271_
timestamp 1649977179
transform -1 0 33304 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1272_
timestamp 1649977179
transform 1 0 26956 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1649977179
transform -1 0 28796 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1649977179
transform 1 0 28060 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1649977179
transform -1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1649977179
transform 1 0 30084 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1278_
timestamp 1649977179
transform -1 0 29808 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1649977179
transform -1 0 31188 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1280_
timestamp 1649977179
transform -1 0 31372 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1281_
timestamp 1649977179
transform 1 0 32568 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1282_
timestamp 1649977179
transform -1 0 33396 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1649977179
transform -1 0 32568 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1284_
timestamp 1649977179
transform 1 0 13156 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1649977179
transform 1 0 25668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1286_
timestamp 1649977179
transform -1 0 32752 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1287_
timestamp 1649977179
transform 1 0 33120 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1288_
timestamp 1649977179
transform -1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1649977179
transform 1 0 32568 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1290_
timestamp 1649977179
transform -1 0 33764 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1649977179
transform -1 0 27232 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1292_
timestamp 1649977179
transform -1 0 27508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1649977179
transform -1 0 26404 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1294_
timestamp 1649977179
transform 1 0 25668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1295_
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1296_
timestamp 1649977179
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 1649977179
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1298_
timestamp 1649977179
transform -1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1299_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10396 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1300_
timestamp 1649977179
transform -1 0 7268 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1649977179
transform -1 0 17848 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1649977179
transform 1 0 6256 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1303_
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1304_
timestamp 1649977179
transform -1 0 5888 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1305_
timestamp 1649977179
transform -1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1306_
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1307_
timestamp 1649977179
transform -1 0 3588 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1308_
timestamp 1649977179
transform 1 0 2576 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1309_
timestamp 1649977179
transform 1 0 3864 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1649977179
transform -1 0 2760 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1649977179
transform 1 0 2852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1312_
timestamp 1649977179
transform 1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1649977179
transform 1 0 5428 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1314_
timestamp 1649977179
transform -1 0 7084 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1315_
timestamp 1649977179
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1649977179
transform 1 0 7452 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1317_
timestamp 1649977179
transform -1 0 5244 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1318_
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1319_
timestamp 1649977179
transform 1 0 19872 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1320_
timestamp 1649977179
transform -1 0 20056 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1649977179
transform 1 0 22448 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1322_
timestamp 1649977179
transform -1 0 23000 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1649977179
transform -1 0 23092 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1324_
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1649977179
transform 1 0 23460 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1326_
timestamp 1649977179
transform -1 0 23276 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1327_
timestamp 1649977179
transform 1 0 25576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1649977179
transform 1 0 21712 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1329_
timestamp 1649977179
transform -1 0 23092 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1330_
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1649977179
transform -1 0 22264 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1332_
timestamp 1649977179
transform 1 0 21344 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1333_
timestamp 1649977179
transform -1 0 24012 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1649977179
transform 1 0 20884 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1335_
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1336_
timestamp 1649977179
transform 1 0 12696 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1649977179
transform -1 0 20056 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1649977179
transform 1 0 16744 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1339_
timestamp 1649977179
transform 1 0 17848 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1340_
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1649977179
transform -1 0 19964 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1649977179
transform -1 0 19964 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _1343_
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1649977179
transform 1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1345_
timestamp 1649977179
transform 1 0 20516 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1649977179
transform -1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1347_
timestamp 1649977179
transform -1 0 17848 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1348_
timestamp 1649977179
transform 1 0 17020 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1349_
timestamp 1649977179
transform 1 0 18216 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1351_
timestamp 1649977179
transform -1 0 17112 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1352_
timestamp 1649977179
transform -1 0 16192 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1649977179
transform 1 0 18032 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1649977179
transform -1 0 17664 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1649977179
transform -1 0 15548 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1356_
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp 1649977179
transform -1 0 16192 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1358_
timestamp 1649977179
transform 1 0 15364 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1359_
timestamp 1649977179
transform 1 0 15088 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1649977179
transform -1 0 17112 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1361_
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1649977179
transform 1 0 23552 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1649977179
transform -1 0 24656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1649977179
transform -1 0 26404 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1365_
timestamp 1649977179
transform -1 0 25392 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1649977179
transform -1 0 25760 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1367_
timestamp 1649977179
transform -1 0 25484 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1649977179
transform -1 0 26312 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1369_
timestamp 1649977179
transform -1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1649977179
transform -1 0 26036 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1371_
timestamp 1649977179
transform -1 0 12880 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1372_
timestamp 1649977179
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1373_
timestamp 1649977179
transform -1 0 24932 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1649977179
transform -1 0 26220 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1375_
timestamp 1649977179
transform -1 0 25576 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1649977179
transform -1 0 22908 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1377_
timestamp 1649977179
transform -1 0 21988 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 1649977179
transform -1 0 24196 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1379_
timestamp 1649977179
transform 1 0 22172 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1649977179
transform -1 0 10672 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1649977179
transform -1 0 11040 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1382_
timestamp 1649977179
transform -1 0 10028 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1383_
timestamp 1649977179
transform -1 0 9568 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1384_
timestamp 1649977179
transform 1 0 11776 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1385_
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1386_
timestamp 1649977179
transform 1 0 7360 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1387_
timestamp 1649977179
transform 1 0 5888 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1388_
timestamp 1649977179
transform 1 0 6716 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1649977179
transform -1 0 4232 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1390_
timestamp 1649977179
transform 1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1391_
timestamp 1649977179
transform 1 0 3128 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1649977179
transform -1 0 3312 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1393_
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1395_
timestamp 1649977179
transform 1 0 6900 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1649977179
transform 1 0 6532 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1397_
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1398_
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1399_
timestamp 1649977179
transform -1 0 14260 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1649977179
transform -1 0 13616 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1649977179
transform 1 0 12420 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1649977179
transform -1 0 14904 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1403_
timestamp 1649977179
transform 1 0 13248 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1404_
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1649977179
transform -1 0 17020 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1406_
timestamp 1649977179
transform -1 0 16744 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1649977179
transform -1 0 17756 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1408_
timestamp 1649977179
transform -1 0 17848 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1649977179
transform 1 0 17664 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1410_
timestamp 1649977179
transform 1 0 16560 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1411_
timestamp 1649977179
transform 1 0 14996 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1412_
timestamp 1649977179
transform -1 0 14628 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1649977179
transform -1 0 13064 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1649977179
transform 1 0 10488 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1415_
timestamp 1649977179
transform -1 0 12236 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1416_
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1417_
timestamp 1649977179
transform -1 0 11040 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1418_
timestamp 1649977179
transform 1 0 9108 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1419_
timestamp 1649977179
transform -1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1420_
timestamp 1649977179
transform -1 0 9936 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1421_
timestamp 1649977179
transform -1 0 9108 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1649977179
transform 1 0 2760 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1423_
timestamp 1649977179
transform 1 0 2576 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1424_
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1425_
timestamp 1649977179
transform 1 0 2668 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1649977179
transform -1 0 4232 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1427_
timestamp 1649977179
transform 1 0 2576 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1428_
timestamp 1649977179
transform -1 0 6440 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1429_
timestamp 1649977179
transform 1 0 5612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1649977179
transform -1 0 8372 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1431_
timestamp 1649977179
transform -1 0 10672 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1649977179
transform 1 0 6900 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1433_
timestamp 1649977179
transform 1 0 9568 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1434_
timestamp 1649977179
transform -1 0 9384 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1435_
timestamp 1649977179
transform -1 0 8464 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1436_
timestamp 1649977179
transform 1 0 8832 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1649977179
transform 1 0 9476 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1438_
timestamp 1649977179
transform 1 0 9200 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1649977179
transform 1 0 10304 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1440_
timestamp 1649977179
transform 1 0 10212 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1441_
timestamp 1649977179
transform 1 0 10212 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1442_
timestamp 1649977179
transform 1 0 10120 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1443_
timestamp 1649977179
transform 1 0 10396 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1444_
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1445_
timestamp 1649977179
transform -1 0 11592 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1446_
timestamp 1649977179
transform -1 0 11224 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1649977179
transform 1 0 9752 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1448_
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1649977179
transform 1 0 9752 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1450_
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1451_
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1452_
timestamp 1649977179
transform -1 0 13616 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1453_
timestamp 1649977179
transform 1 0 13432 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1454_
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1455_
timestamp 1649977179
transform 1 0 14444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1456_
timestamp 1649977179
transform 1 0 14996 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1649977179
transform 1 0 15824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 1649977179
transform -1 0 10488 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1649977179
transform -1 0 11960 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1461_
timestamp 1649977179
transform 1 0 10120 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1649977179
transform 1 0 10580 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1463_
timestamp 1649977179
transform 1 0 12696 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1464_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1465_
timestamp 1649977179
transform -1 0 13248 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1466_
timestamp 1649977179
transform 1 0 12420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1467_
timestamp 1649977179
transform -1 0 15824 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1468_
timestamp 1649977179
transform -1 0 14628 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1469_
timestamp 1649977179
transform 1 0 17848 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1649977179
transform -1 0 18400 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1471_
timestamp 1649977179
transform -1 0 22264 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1472_
timestamp 1649977179
transform -1 0 21344 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1473_
timestamp 1649977179
transform -1 0 20424 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1474_
timestamp 1649977179
transform -1 0 19596 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1475_
timestamp 1649977179
transform -1 0 24748 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1476_
timestamp 1649977179
transform 1 0 19780 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1477_
timestamp 1649977179
transform -1 0 21896 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1479_
timestamp 1649977179
transform -1 0 22540 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 1649977179
transform 1 0 18952 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1481_
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1649977179
transform 1 0 18952 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1483_
timestamp 1649977179
transform -1 0 18768 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1649977179
transform 1 0 17204 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1485_
timestamp 1649977179
transform -1 0 18584 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1486_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7728 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1487_
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1488_
timestamp 1649977179
transform -1 0 19504 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1649977179
transform -1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1490_
timestamp 1649977179
transform -1 0 19412 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1649977179
transform -1 0 19688 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1649977179
transform -1 0 17112 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1649977179
transform -1 0 18032 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1495_
timestamp 1649977179
transform 1 0 15364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1496_
timestamp 1649977179
transform -1 0 16928 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1497_
timestamp 1649977179
transform 1 0 14536 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 1649977179
transform -1 0 17112 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1499_
timestamp 1649977179
transform -1 0 15916 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1649977179
transform 1 0 18308 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1649977179
transform -1 0 20332 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1649977179
transform 1 0 19320 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1649977179
transform -1 0 19228 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1504_
timestamp 1649977179
transform 1 0 25576 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1505_
timestamp 1649977179
transform 1 0 22448 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1649977179
transform 1 0 31096 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1507_
timestamp 1649977179
transform 1 0 24932 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1508_
timestamp 1649977179
transform -1 0 30728 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1649977179
transform 1 0 29808 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1510_
timestamp 1649977179
transform -1 0 30912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 1649977179
transform 1 0 29256 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1512_
timestamp 1649977179
transform -1 0 30820 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1513_
timestamp 1649977179
transform -1 0 28152 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1514_
timestamp 1649977179
transform 1 0 26956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1515_
timestamp 1649977179
transform -1 0 28060 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1516_
timestamp 1649977179
transform 1 0 26496 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1517_
timestamp 1649977179
transform -1 0 18768 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1518_
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1519_
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 1649977179
transform -1 0 22264 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1521_
timestamp 1649977179
transform 1 0 19780 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1522_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8004 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1523_
timestamp 1649977179
transform -1 0 8096 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1524_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1525_
timestamp 1649977179
transform -1 0 7268 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1526_
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1527_
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1528_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_2  _1529_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1530_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1531_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 34960 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1649977179
transform 1 0 23276 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1649977179
transform 1 0 22448 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1534_
timestamp 1649977179
transform -1 0 28980 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1535_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1536_
timestamp 1649977179
transform 1 0 4692 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1537_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6716 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1538_
timestamp 1649977179
transform 1 0 9384 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1539_
timestamp 1649977179
transform 1 0 9936 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1540_
timestamp 1649977179
transform -1 0 10672 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1541_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5888 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1542_
timestamp 1649977179
transform -1 0 35052 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1649977179
transform 1 0 22264 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1649977179
transform 1 0 22356 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 1649977179
transform -1 0 28980 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1546_
timestamp 1649977179
transform -1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1649977179
transform 1 0 4048 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1548_
timestamp 1649977179
transform 1 0 4692 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1549_
timestamp 1649977179
transform 1 0 9200 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1550_
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1649977179
transform -1 0 7820 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1552_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1553_
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1554_
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1555_
timestamp 1649977179
transform -1 0 36064 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1556_
timestamp 1649977179
transform 1 0 23000 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1557_
timestamp 1649977179
transform 1 0 22172 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1558_
timestamp 1649977179
transform -1 0 29072 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1559_
timestamp 1649977179
transform -1 0 24840 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1560_
timestamp 1649977179
transform 1 0 4048 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1561_
timestamp 1649977179
transform 1 0 4784 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1649977179
transform -1 0 11960 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1563_
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1564_
timestamp 1649977179
transform -1 0 7452 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1565_
timestamp 1649977179
transform -1 0 6440 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1566_
timestamp 1649977179
transform 1 0 5152 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1567_
timestamp 1649977179
transform 1 0 6164 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1568_
timestamp 1649977179
transform 1 0 35052 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1569_
timestamp 1649977179
transform -1 0 36432 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1570_
timestamp 1649977179
transform 1 0 33764 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1571_
timestamp 1649977179
transform -1 0 36248 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1649977179
transform -1 0 36800 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1573_
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1574_
timestamp 1649977179
transform 1 0 28796 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1649977179
transform 1 0 22448 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1576_
timestamp 1649977179
transform 1 0 30084 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1578_
timestamp 1649977179
transform 1 0 20424 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1580_
timestamp 1649977179
transform 1 0 19412 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1581_
timestamp 1649977179
transform 1 0 29532 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1649977179
transform -1 0 30176 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1583_
timestamp 1649977179
transform 1 0 31372 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1584_
timestamp 1649977179
transform 1 0 32108 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1585_
timestamp 1649977179
transform 1 0 30544 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1586_
timestamp 1649977179
transform -1 0 33028 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1587_
timestamp 1649977179
transform -1 0 31832 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1588_
timestamp 1649977179
transform -1 0 29716 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1589_
timestamp 1649977179
transform 1 0 11592 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1590_
timestamp 1649977179
transform -1 0 12604 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1591_
timestamp 1649977179
transform 1 0 11040 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1592_
timestamp 1649977179
transform -1 0 12328 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1593_
timestamp 1649977179
transform 1 0 7268 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1594_
timestamp 1649977179
transform 1 0 8648 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1595_
timestamp 1649977179
transform 1 0 19780 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1596_
timestamp 1649977179
transform 1 0 23000 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1597_
timestamp 1649977179
transform 1 0 20424 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1598_
timestamp 1649977179
transform 1 0 22724 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1599_
timestamp 1649977179
transform -1 0 14720 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1600_
timestamp 1649977179
transform -1 0 13616 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1601_
timestamp 1649977179
transform -1 0 9476 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1602_
timestamp 1649977179
transform 1 0 5060 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1603_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1604_
timestamp 1649977179
transform -1 0 8004 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1649977179
transform -1 0 37444 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1606_
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1649977179
transform -1 0 31464 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 1649977179
transform -1 0 32844 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1609_
timestamp 1649977179
transform -1 0 30820 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1610_
timestamp 1649977179
transform -1 0 15640 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1611_
timestamp 1649977179
transform -1 0 16376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1612_
timestamp 1649977179
transform 1 0 8280 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1613_
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1614_
timestamp 1649977179
transform 1 0 19780 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1615_
timestamp 1649977179
transform -1 0 17480 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1616_
timestamp 1649977179
transform 1 0 15180 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1617_
timestamp 1649977179
transform 1 0 15456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1618_
timestamp 1649977179
transform -1 0 10120 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1619_
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1620_
timestamp 1649977179
transform -1 0 7636 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1621_
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1622_
timestamp 1649977179
transform -1 0 36340 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1649977179
transform 1 0 29716 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1624_
timestamp 1649977179
transform 1 0 31004 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1649977179
transform -1 0 32936 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1626_
timestamp 1649977179
transform -1 0 32660 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1627_
timestamp 1649977179
transform 1 0 12604 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1628_
timestamp 1649977179
transform 1 0 13340 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1649977179
transform 1 0 23092 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1649977179
transform -1 0 23828 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1631_
timestamp 1649977179
transform -1 0 14812 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1632_
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1633_
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1634_
timestamp 1649977179
transform -1 0 36248 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1649977179
transform 1 0 30728 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp 1649977179
transform 1 0 30820 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1637_
timestamp 1649977179
transform -1 0 33120 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1638_
timestamp 1649977179
transform -1 0 32476 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1639_
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp 1649977179
transform 1 0 17020 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1641_
timestamp 1649977179
transform -1 0 23552 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1642_
timestamp 1649977179
transform -1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1643_
timestamp 1649977179
transform -1 0 18768 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1644_
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1645_
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1646_
timestamp 1649977179
transform 1 0 8372 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1647_
timestamp 1649977179
transform -1 0 36248 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 1649977179
transform 1 0 30636 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1649977179
transform 1 0 31004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1650_
timestamp 1649977179
transform -1 0 33028 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1651_
timestamp 1649977179
transform -1 0 32660 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1652_
timestamp 1649977179
transform 1 0 15088 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1653_
timestamp 1649977179
transform 1 0 18492 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1649977179
transform -1 0 23828 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1655_
timestamp 1649977179
transform -1 0 23920 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1656_
timestamp 1649977179
transform -1 0 19688 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1657_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1658_
timestamp 1649977179
transform -1 0 10856 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1659_
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1649977179
transform -1 0 35696 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1649977179
transform 1 0 27876 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1649977179
transform 1 0 29440 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1663_
timestamp 1649977179
transform -1 0 34224 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1664_
timestamp 1649977179
transform -1 0 29900 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1665_
timestamp 1649977179
transform 1 0 11592 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1666_
timestamp 1649977179
transform 1 0 18032 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1667_
timestamp 1649977179
transform 1 0 22080 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1668_
timestamp 1649977179
transform -1 0 23644 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1669_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18768 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1670_
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1671_
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1649977179
transform -1 0 35512 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1673_
timestamp 1649977179
transform 1 0 27784 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1674_
timestamp 1649977179
transform 1 0 27600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1649977179
transform -1 0 34040 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1676_
timestamp 1649977179
transform -1 0 30084 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 1649977179
transform 1 0 12328 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1678_
timestamp 1649977179
transform 1 0 17296 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1679_
timestamp 1649977179
transform -1 0 21712 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1680_
timestamp 1649977179
transform -1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1681_
timestamp 1649977179
transform -1 0 19688 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1682_
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1683_
timestamp 1649977179
transform -1 0 12788 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1684_
timestamp 1649977179
transform -1 0 37536 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1685_
timestamp 1649977179
transform 1 0 23736 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1686_
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1687_
timestamp 1649977179
transform -1 0 34040 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1688_
timestamp 1649977179
transform -1 0 24932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1689_
timestamp 1649977179
transform 1 0 11684 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1690_
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1691_
timestamp 1649977179
transform 1 0 20424 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1692_
timestamp 1649977179
transform -1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1693_
timestamp 1649977179
transform -1 0 17940 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1694_
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1695_
timestamp 1649977179
transform -1 0 6164 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1696_
timestamp 1649977179
transform -1 0 36524 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1697_
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1698_
timestamp 1649977179
transform 1 0 22908 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1699_
timestamp 1649977179
transform -1 0 33028 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1700_
timestamp 1649977179
transform -1 0 25024 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1701_
timestamp 1649977179
transform 1 0 12420 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1702_
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1703_
timestamp 1649977179
transform -1 0 21436 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1704_
timestamp 1649977179
transform -1 0 20516 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1705_
timestamp 1649977179
transform -1 0 18768 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1706_
timestamp 1649977179
transform 1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1707_
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1708_
timestamp 1649977179
transform -1 0 2208 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1709_
timestamp 1649977179
transform -1 0 1932 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1710_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1649977179
transform 1 0 1840 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1649977179
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1649977179
transform 1 0 1840 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1649977179
transform 1 0 3404 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1649977179
transform 1 0 8280 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1649977179
transform -1 0 14996 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1649977179
transform 1 0 1840 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1649977179
transform 1 0 2116 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1649977179
transform 1 0 4968 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1649977179
transform -1 0 6992 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1649977179
transform -1 0 15088 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1649977179
transform -1 0 16928 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1649977179
transform 1 0 14904 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1649977179
transform -1 0 12972 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1649977179
transform -1 0 12972 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1649977179
transform -1 0 13064 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1649977179
transform -1 0 15548 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1649977179
transform 1 0 27600 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1649977179
transform 1 0 27324 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1649977179
transform 1 0 27324 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1649977179
transform 1 0 30268 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1649977179
transform 1 0 30912 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1649977179
transform -1 0 38456 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1649977179
transform -1 0 38548 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1649977179
transform -1 0 38732 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1649977179
transform -1 0 38732 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1649977179
transform -1 0 38732 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1649977179
transform -1 0 38732 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1649977179
transform 1 0 33120 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1649977179
transform 1 0 29532 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1649977179
transform 1 0 27416 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1649977179
transform 1 0 27692 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1649977179
transform 1 0 29900 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1649977179
transform 1 0 30176 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1649977179
transform 1 0 31832 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1649977179
transform -1 0 34776 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1649977179
transform -1 0 36616 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1649977179
transform -1 0 36156 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1649977179
transform -1 0 35972 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1649977179
transform -1 0 37168 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1649977179
transform 1 0 31556 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1649977179
transform 1 0 2760 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1649977179
transform 1 0 7176 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1649977179
transform 1 0 19872 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1649977179
transform -1 0 20148 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1649977179
transform -1 0 21528 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1649977179
transform -1 0 20792 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1649977179
transform 1 0 16100 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1649977179
transform 1 0 8464 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1649977179
transform 1 0 6992 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1649977179
transform -1 0 12972 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1649977179
transform 1 0 12144 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1649977179
transform 1 0 14812 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1649977179
transform -1 0 26036 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1649977179
transform -1 0 24472 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1649977179
transform -1 0 27600 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1649977179
transform -1 0 25852 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1649977179
transform -1 0 27048 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1649977179
transform -1 0 27324 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1649977179
transform 1 0 25576 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1649977179
transform 1 0 23276 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1649977179
transform -1 0 24564 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1649977179
transform 1 0 27416 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1649977179
transform 1 0 29808 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1649977179
transform -1 0 33304 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1649977179
transform -1 0 33580 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1649977179
transform -1 0 32936 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1649977179
transform -1 0 33580 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1649977179
transform -1 0 28704 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1649977179
transform 1 0 22632 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1649977179
transform -1 0 13248 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1649977179
transform -1 0 13524 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1649977179
transform -1 0 18124 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1649977179
transform -1 0 32384 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1649977179
transform -1 0 31648 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1649977179
transform -1 0 31004 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1649977179
transform -1 0 28888 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1649977179
transform -1 0 28796 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1649977179
transform -1 0 21252 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1649977179
transform 1 0 34500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1649977179
transform 1 0 37720 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1649977179
transform 1 0 37904 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1649977179
transform 1 0 38548 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1649977179
transform -1 0 39928 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1649977179
transform 1 0 35328 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1649977179
transform 1 0 38640 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1649977179
transform 1 0 38732 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1649977179
transform -1 0 40020 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1649977179
transform -1 0 40204 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1649977179
transform -1 0 40204 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1649977179
transform 1 0 32752 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1649977179
transform 1 0 33488 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1649977179
transform -1 0 37352 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1649977179
transform 1 0 36340 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1649977179
transform -1 0 40020 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1649977179
transform -1 0 37904 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1649977179
transform 1 0 40480 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1649977179
transform -1 0 40112 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1649977179
transform 1 0 37904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1649977179
transform -1 0 39376 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1649977179
transform -1 0 40112 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1649977179
transform -1 0 37352 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1649977179
transform -1 0 26404 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1649977179
transform -1 0 24932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1649977179
transform 1 0 29624 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1649977179
transform 1 0 28428 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1649977179
transform -1 0 32292 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1649977179
transform -1 0 34224 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1649977179
transform -1 0 34316 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1649977179
transform -1 0 35328 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1649977179
transform -1 0 36156 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1649977179
transform -1 0 26496 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1649977179
transform 1 0 4232 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1649977179
transform 1 0 2392 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1649977179
transform -1 0 3312 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1649977179
transform 1 0 6072 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1649977179
transform 1 0 5612 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1649977179
transform -1 0 23920 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1649977179
transform -1 0 24932 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1649977179
transform -1 0 25852 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1649977179
transform 1 0 22448 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1649977179
transform -1 0 21712 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1649977179
transform 1 0 16652 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1649977179
transform 1 0 17940 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1649977179
transform 1 0 15272 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1649977179
transform 1 0 25576 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1649977179
transform -1 0 27324 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1649977179
transform 1 0 26772 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1649977179
transform 1 0 24932 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1649977179
transform 1 0 24932 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1649977179
transform 1 0 21896 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1649977179
transform 1 0 22356 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1649977179
transform -1 0 7820 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1649977179
transform 1 0 2576 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1649977179
transform -1 0 4048 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1649977179
transform 1 0 6808 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1649977179
transform 1 0 6164 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1649977179
transform 1 0 11776 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1649977179
transform -1 0 20240 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1649977179
transform 1 0 11684 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1649977179
transform 1 0 2300 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1649977179
transform 1 0 2116 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1649977179
transform 1 0 1840 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1649977179
transform 1 0 5428 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1649977179
transform 1 0 6072 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1649977179
transform 1 0 6716 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1649977179
transform 1 0 8372 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1649977179
transform 1 0 8924 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1649977179
transform 1 0 10488 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1649977179
transform 1 0 9200 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1649977179
transform 1 0 8280 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1649977179
transform 1 0 7912 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1649977179
transform 1 0 9568 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1649977179
transform 1 0 12144 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1649977179
transform 1 0 14260 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1649977179
transform 1 0 21988 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1649977179
transform 1 0 22448 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1649977179
transform -1 0 19596 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1649977179
transform 1 0 15364 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1649977179
transform 1 0 19320 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1649977179
transform 1 0 30176 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1649977179
transform -1 0 32108 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1649977179
transform 1 0 30176 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1649977179
transform 1 0 27048 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1649977179
transform 1 0 26036 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1649977179
transform 1 0 19872 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1649977179
transform -1 0 8188 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1649977179
transform -1 0 8464 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1649977179
transform -1 0 7820 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1649977179
transform -1 0 11040 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1649977179
transform 1 0 9936 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1649977179
transform -1 0 13156 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1649977179
transform 1 0 3036 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1649977179
transform -1 0 8648 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1649977179
transform 1 0 1840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21068 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1649977179
transform -1 0 12236 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1649977179
transform 1 0 31188 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1649977179
transform 1 0 3128 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1649977179
transform 1 0 5704 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1649977179
transform 1 0 16100 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1649977179
transform 1 0 13064 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1649977179
transform -1 0 7268 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1649977179
transform 1 0 5704 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1649977179
transform -1 0 5244 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1649977179
transform 1 0 8924 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1649977179
transform -1 0 18584 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1649977179
transform 1 0 20240 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1649977179
transform 1 0 16008 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1649977179
transform -1 0 23276 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1649977179
transform 1 0 27324 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1649977179
transform 1 0 26772 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1649977179
transform 1 0 32016 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1649977179
transform -1 0 39008 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1649977179
transform 1 0 38916 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1649977179
transform 1 0 30360 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1649977179
transform -1 0 28152 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1649977179
transform 1 0 33948 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1649977179
transform 1 0 39560 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1649977179
transform 1 0 36432 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1649977179
transform -1 0 36984 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1649977179
transform -1 0 31096 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1649977179
transform -1 0 26864 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1649977179
transform 1 0 27416 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1649977179
transform -1 0 23644 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1649977179
transform 1 0 19596 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1649977179
transform 1 0 12696 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_32_wb_clk_i
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_33_wb_clk_i
timestamp 1649977179
transform 1 0 6624 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 2392 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1649977179
transform -1 0 7728 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1649977179
transform -1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1649977179
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform -1 0 5612 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform -1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1649977179
transform 1 0 8464 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input22
timestamp 1649977179
transform -1 0 10948 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1649977179
transform -1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 1932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform -1 0 2668 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform -1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1649977179
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform -1 0 10028 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_43 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 53728 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_44
timestamp 1649977179
transform -1 0 50600 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_45
timestamp 1649977179
transform -1 0 55568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_46
timestamp 1649977179
transform -1 0 41216 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_47
timestamp 1649977179
transform -1 0 42780 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_48
timestamp 1649977179
transform -1 0 44344 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_49
timestamp 1649977179
transform -1 0 45908 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_50
timestamp 1649977179
transform -1 0 47840 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_51
timestamp 1649977179
transform -1 0 49036 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_52
timestamp 1649977179
transform -1 0 13064 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_53
timestamp 1649977179
transform -1 0 14628 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_54
timestamp 1649977179
transform -1 0 16192 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_55
timestamp 1649977179
transform -1 0 17756 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_56
timestamp 1649977179
transform -1 0 19504 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_57
timestamp 1649977179
transform -1 0 20884 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_58
timestamp 1649977179
transform -1 0 22448 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_59
timestamp 1649977179
transform -1 0 24656 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_60
timestamp 1649977179
transform -1 0 25576 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_61
timestamp 1649977179
transform -1 0 27232 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_62
timestamp 1649977179
transform -1 0 28704 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_63
timestamp 1649977179
transform -1 0 30268 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_64
timestamp 1649977179
transform -1 0 32384 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_65
timestamp 1649977179
transform -1 0 33396 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_66
timestamp 1649977179
transform -1 0 34960 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_67
timestamp 1649977179
transform -1 0 36524 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_68
timestamp 1649977179
transform -1 0 38088 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_69
timestamp 1649977179
transform -1 0 40112 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_70
timestamp 1649977179
transform -1 0 52164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_71
timestamp 1649977179
transform -1 0 8372 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_72
timestamp 1649977179
transform -1 0 9936 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_73
timestamp 1649977179
transform -1 0 11776 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_74
timestamp 1649977179
transform -1 0 5244 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_75
timestamp 1649977179
transform -1 0 6808 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_76
timestamp 1649977179
transform -1 0 2116 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_77
timestamp 1649977179
transform -1 0 4048 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_78
timestamp 1649977179
transform -1 0 56856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_79
timestamp 1649977179
transform -1 0 58236 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_80
timestamp 1649977179
transform 1 0 57960 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_81
timestamp 1649977179
transform 1 0 57960 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_82
timestamp 1649977179
transform 1 0 57316 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_83
timestamp 1649977179
transform 1 0 57960 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_84
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_85
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_86
timestamp 1649977179
transform -1 0 51428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_87
timestamp 1649977179
transform -1 0 52440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_88
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_89
timestamp 1649977179
transform -1 0 52072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_90
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_91
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_92
timestamp 1649977179
transform -1 0 53728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_93
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_94
timestamp 1649977179
transform -1 0 52992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_95
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_96
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_97
timestamp 1649977179
transform -1 0 52440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_98
timestamp 1649977179
transform -1 0 53084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_99
timestamp 1649977179
transform -1 0 54372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_100
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_101
timestamp 1649977179
transform -1 0 53636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_102
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103
timestamp 1649977179
transform -1 0 53728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform -1 0 54280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform -1 0 54924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform -1 0 54372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform -1 0 55568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform -1 0 54004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform -1 0 54648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform -1 0 55568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform -1 0 56212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform -1 0 55292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform -1 0 56212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform 1 0 57960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform 1 0 57316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform 1 0 57960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform 1 0 57960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform 1 0 57960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform 1 0 57960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform 1 0 57960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform 1 0 57960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform 1 0 57960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform 1 0 57960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform 1 0 57960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform 1 0 57960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform 1 0 57960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform 1 0 57960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform 1 0 57960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform 1 0 57960 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform 1 0 57960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform 1 0 57960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform 1 0 57960 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform 1 0 57960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform 1 0 57960 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform 1 0 57960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform 1 0 57960 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform 1 0 57960 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform 1 0 57960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform 1 0 57960 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform 1 0 57960 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform 1 0 57960 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform 1 0 57960 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform 1 0 57960 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform 1 0 57960 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform 1 0 57960 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform 1 0 57960 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform 1 0 57960 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform 1 0 57960 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform 1 0 57960 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform 1 0 57960 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform 1 0 57960 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform -1 0 51796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform -1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform -1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform -1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform -1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform -1 0 19872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform -1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform -1 0 21528 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform -1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform -1 0 23736 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform 1 0 25392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform -1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform -1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform -1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform 1 0 29348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform -1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform 1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform -1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform -1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 33672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform -1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform -1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform -1 0 34960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform -1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform -1 0 35052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform -1 0 35696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform -1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform -1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform -1 0 36984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform -1 0 37812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform -1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform -1 0 42780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform -1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform -1 0 45264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform -1 0 45908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform -1 0 46552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform -1 0 47196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_278
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_279
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_280
timestamp 1649977179
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_281
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_282
timestamp 1649977179
transform -1 0 48668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_283
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_284
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_285
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_286
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_287
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_288
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_289
timestamp 1649977179
transform -1 0 50508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_290
timestamp 1649977179
transform -1 0 51152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_291
timestamp 1649977179
transform 1 0 57960 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_292
timestamp 1649977179
transform 1 0 57960 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_293
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_294
timestamp 1649977179
transform -1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_295
timestamp 1649977179
transform -1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_296
timestamp 1649977179
transform 1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_297
timestamp 1649977179
transform -1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_298
timestamp 1649977179
transform -1 0 11684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_299
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_300
timestamp 1649977179
transform -1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_301
timestamp 1649977179
transform 1 0 11592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_302
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_303
timestamp 1649977179
transform -1 0 13064 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_304
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_305
timestamp 1649977179
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_306
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_307
timestamp 1649977179
transform 1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_308
timestamp 1649977179
transform -1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_309
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_310
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_311
timestamp 1649977179
transform 1 0 13984 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_312
timestamp 1649977179
transform -1 0 15640 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 CMP_out_c
port 0 nsew signal tristate
flabel metal2 s 50250 59200 50306 60000 0 FreeSans 224 90 0 0 OTA_out_c
port 1 nsew signal tristate
flabel metal2 s 54942 59200 54998 60000 0 FreeSans 224 90 0 0 OTA_sh_c
port 2 nsew signal tristate
flabel metal2 s 40866 59200 40922 60000 0 FreeSans 224 90 0 0 Pd10_a
port 3 nsew signal tristate
flabel metal2 s 42430 59200 42486 60000 0 FreeSans 224 90 0 0 Pd10_b
port 4 nsew signal tristate
flabel metal2 s 43994 59200 44050 60000 0 FreeSans 224 90 0 0 Pd11_a
port 5 nsew signal tristate
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 Pd11_b
port 6 nsew signal tristate
flabel metal2 s 47122 59200 47178 60000 0 FreeSans 224 90 0 0 Pd12_a
port 7 nsew signal tristate
flabel metal2 s 48686 59200 48742 60000 0 FreeSans 224 90 0 0 Pd12_b
port 8 nsew signal tristate
flabel metal2 s 12714 59200 12770 60000 0 FreeSans 224 90 0 0 Pd1_a
port 9 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 Pd1_b
port 10 nsew signal tristate
flabel metal2 s 15842 59200 15898 60000 0 FreeSans 224 90 0 0 Pd2_a
port 11 nsew signal tristate
flabel metal2 s 17406 59200 17462 60000 0 FreeSans 224 90 0 0 Pd2_b
port 12 nsew signal tristate
flabel metal2 s 18970 59200 19026 60000 0 FreeSans 224 90 0 0 Pd3_a
port 13 nsew signal tristate
flabel metal2 s 20534 59200 20590 60000 0 FreeSans 224 90 0 0 Pd3_b
port 14 nsew signal tristate
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 Pd4_a
port 15 nsew signal tristate
flabel metal2 s 23662 59200 23718 60000 0 FreeSans 224 90 0 0 Pd4_b
port 16 nsew signal tristate
flabel metal2 s 25226 59200 25282 60000 0 FreeSans 224 90 0 0 Pd5_a
port 17 nsew signal tristate
flabel metal2 s 26790 59200 26846 60000 0 FreeSans 224 90 0 0 Pd5_b
port 18 nsew signal tristate
flabel metal2 s 28354 59200 28410 60000 0 FreeSans 224 90 0 0 Pd6_a
port 19 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 Pd6_b
port 20 nsew signal tristate
flabel metal2 s 31482 59200 31538 60000 0 FreeSans 224 90 0 0 Pd7_a
port 21 nsew signal tristate
flabel metal2 s 33046 59200 33102 60000 0 FreeSans 224 90 0 0 Pd7_b
port 22 nsew signal tristate
flabel metal2 s 34610 59200 34666 60000 0 FreeSans 224 90 0 0 Pd8_a
port 23 nsew signal tristate
flabel metal2 s 36174 59200 36230 60000 0 FreeSans 224 90 0 0 Pd8_b
port 24 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 Pd9_a
port 25 nsew signal tristate
flabel metal2 s 39302 59200 39358 60000 0 FreeSans 224 90 0 0 Pd9_b
port 26 nsew signal tristate
flabel metal2 s 51814 59200 51870 60000 0 FreeSans 224 90 0 0 SH_out_c
port 27 nsew signal tristate
flabel metal2 s 8022 59200 8078 60000 0 FreeSans 224 90 0 0 Sh
port 28 nsew signal tristate
flabel metal2 s 9586 59200 9642 60000 0 FreeSans 224 90 0 0 Sh_cmp
port 29 nsew signal tristate
flabel metal2 s 11150 59200 11206 60000 0 FreeSans 224 90 0 0 Sh_rst
port 30 nsew signal tristate
flabel metal2 s 4894 59200 4950 60000 0 FreeSans 224 90 0 0 Sw1
port 31 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 Sw2
port 32 nsew signal tristate
flabel metal2 s 1766 59200 1822 60000 0 FreeSans 224 90 0 0 Vd1
port 33 nsew signal tristate
flabel metal2 s 3330 59200 3386 60000 0 FreeSans 224 90 0 0 Vd2
port 34 nsew signal tristate
flabel metal2 s 56506 59200 56562 60000 0 FreeSans 224 90 0 0 Vref_cmp_c
port 35 nsew signal tristate
flabel metal2 s 58070 59200 58126 60000 0 FreeSans 224 90 0 0 Vref_sel_c
port 36 nsew signal tristate
flabel metal3 s 59200 52368 60000 52488 0 FreeSans 480 0 0 0 clk_o
port 37 nsew signal tristate
flabel metal3 s 59200 59168 60000 59288 0 FreeSans 480 0 0 0 counter_rst
port 38 nsew signal tristate
flabel metal3 s 59200 57808 60000 57928 0 FreeSans 480 0 0 0 data_o
port 39 nsew signal tristate
flabel metal3 s 59200 55088 60000 55208 0 FreeSans 480 0 0 0 done_o
port 40 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 io_in[0]
port 41 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_in[10]
port 42 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[11]
port 43 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 io_in[12]
port 44 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 io_in[13]
port 45 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 io_in[14]
port 46 nsew signal input
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 io_in[15]
port 47 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_in[16]
port 48 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 io_in[17]
port 49 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 io_in[18]
port 50 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_in[19]
port 51 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_in[1]
port 52 nsew signal input
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 io_in[20]
port 53 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 io_in[21]
port 54 nsew signal input
flabel metal3 s 0 35096 800 35216 0 FreeSans 480 0 0 0 io_in[22]
port 55 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 io_in[23]
port 56 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_in[24]
port 57 nsew signal input
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 io_in[25]
port 58 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 io_in[26]
port 59 nsew signal input
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 io_in[27]
port 60 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 io_in[28]
port 61 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_in[29]
port 62 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_in[2]
port 63 nsew signal input
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 io_in[30]
port 64 nsew signal input
flabel metal3 s 0 48560 800 48680 0 FreeSans 480 0 0 0 io_in[31]
port 65 nsew signal input
flabel metal3 s 0 50056 800 50176 0 FreeSans 480 0 0 0 io_in[32]
port 66 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 io_in[33]
port 67 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 io_in[34]
port 68 nsew signal input
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 io_in[35]
port 69 nsew signal input
flabel metal3 s 0 56040 800 56160 0 FreeSans 480 0 0 0 io_in[36]
port 70 nsew signal input
flabel metal3 s 0 57536 800 57656 0 FreeSans 480 0 0 0 io_in[37]
port 71 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 io_in[3]
port 72 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_in[4]
port 73 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[5]
port 74 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_in[6]
port 75 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_in[7]
port 76 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_in[8]
port 77 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_in[9]
port 78 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 79 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 80 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 81 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 82 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 83 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 84 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 85 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 86 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 87 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 88 nsew signal tristate
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 89 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 90 nsew signal tristate
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 91 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 92 nsew signal tristate
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 93 nsew signal tristate
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 94 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 95 nsew signal tristate
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 96 nsew signal tristate
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 97 nsew signal tristate
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 98 nsew signal tristate
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 99 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 100 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 101 nsew signal tristate
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 102 nsew signal tristate
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 103 nsew signal tristate
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 104 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 105 nsew signal tristate
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 106 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 107 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 108 nsew signal tristate
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 109 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 110 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 111 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 112 nsew signal tristate
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 113 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 114 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 115 nsew signal tristate
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 116 nsew signal tristate
flabel metal3 s 59200 688 60000 808 0 FreeSans 480 0 0 0 io_out[0]
port 117 nsew signal tristate
flabel metal3 s 59200 14288 60000 14408 0 FreeSans 480 0 0 0 io_out[10]
port 118 nsew signal tristate
flabel metal3 s 59200 15648 60000 15768 0 FreeSans 480 0 0 0 io_out[11]
port 119 nsew signal tristate
flabel metal3 s 59200 17008 60000 17128 0 FreeSans 480 0 0 0 io_out[12]
port 120 nsew signal tristate
flabel metal3 s 59200 18368 60000 18488 0 FreeSans 480 0 0 0 io_out[13]
port 121 nsew signal tristate
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 io_out[14]
port 122 nsew signal tristate
flabel metal3 s 59200 21088 60000 21208 0 FreeSans 480 0 0 0 io_out[15]
port 123 nsew signal tristate
flabel metal3 s 59200 22448 60000 22568 0 FreeSans 480 0 0 0 io_out[16]
port 124 nsew signal tristate
flabel metal3 s 59200 23808 60000 23928 0 FreeSans 480 0 0 0 io_out[17]
port 125 nsew signal tristate
flabel metal3 s 59200 25168 60000 25288 0 FreeSans 480 0 0 0 io_out[18]
port 126 nsew signal tristate
flabel metal3 s 59200 26528 60000 26648 0 FreeSans 480 0 0 0 io_out[19]
port 127 nsew signal tristate
flabel metal3 s 59200 2048 60000 2168 0 FreeSans 480 0 0 0 io_out[1]
port 128 nsew signal tristate
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 io_out[20]
port 129 nsew signal tristate
flabel metal3 s 59200 29248 60000 29368 0 FreeSans 480 0 0 0 io_out[21]
port 130 nsew signal tristate
flabel metal3 s 59200 30608 60000 30728 0 FreeSans 480 0 0 0 io_out[22]
port 131 nsew signal tristate
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 io_out[23]
port 132 nsew signal tristate
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 io_out[24]
port 133 nsew signal tristate
flabel metal3 s 59200 34688 60000 34808 0 FreeSans 480 0 0 0 io_out[25]
port 134 nsew signal tristate
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 io_out[26]
port 135 nsew signal tristate
flabel metal3 s 59200 37408 60000 37528 0 FreeSans 480 0 0 0 io_out[27]
port 136 nsew signal tristate
flabel metal3 s 59200 38768 60000 38888 0 FreeSans 480 0 0 0 io_out[28]
port 137 nsew signal tristate
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 io_out[29]
port 138 nsew signal tristate
flabel metal3 s 59200 3408 60000 3528 0 FreeSans 480 0 0 0 io_out[2]
port 139 nsew signal tristate
flabel metal3 s 59200 41488 60000 41608 0 FreeSans 480 0 0 0 io_out[30]
port 140 nsew signal tristate
flabel metal3 s 59200 42848 60000 42968 0 FreeSans 480 0 0 0 io_out[31]
port 141 nsew signal tristate
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 io_out[32]
port 142 nsew signal tristate
flabel metal3 s 59200 45568 60000 45688 0 FreeSans 480 0 0 0 io_out[33]
port 143 nsew signal tristate
flabel metal3 s 59200 46928 60000 47048 0 FreeSans 480 0 0 0 io_out[34]
port 144 nsew signal tristate
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 io_out[35]
port 145 nsew signal tristate
flabel metal3 s 59200 49648 60000 49768 0 FreeSans 480 0 0 0 io_out[36]
port 146 nsew signal tristate
flabel metal3 s 59200 51008 60000 51128 0 FreeSans 480 0 0 0 io_out[37]
port 147 nsew signal tristate
flabel metal3 s 59200 4768 60000 4888 0 FreeSans 480 0 0 0 io_out[3]
port 148 nsew signal tristate
flabel metal3 s 59200 6128 60000 6248 0 FreeSans 480 0 0 0 io_out[4]
port 149 nsew signal tristate
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 150 nsew signal tristate
flabel metal3 s 59200 8848 60000 8968 0 FreeSans 480 0 0 0 io_out[6]
port 151 nsew signal tristate
flabel metal3 s 59200 10208 60000 10328 0 FreeSans 480 0 0 0 io_out[7]
port 152 nsew signal tristate
flabel metal3 s 59200 11568 60000 11688 0 FreeSans 480 0 0 0 io_out[8]
port 153 nsew signal tristate
flabel metal3 s 59200 12928 60000 13048 0 FreeSans 480 0 0 0 io_out[9]
port 154 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 irq[0]
port 155 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 irq[1]
port 156 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 irq[2]
port 157 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 158 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 159 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 160 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 161 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 162 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 163 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 164 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 165 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 166 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 167 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 168 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 169 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 170 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 171 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 172 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 173 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 174 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 175 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 176 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 177 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 178 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 179 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 180 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 181 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 182 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 183 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 184 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 185 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 186 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 187 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 188 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 189 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 190 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 191 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 192 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 193 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 194 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 195 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 196 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 197 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 198 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 199 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 200 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 201 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 202 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 203 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 204 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 205 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 206 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 207 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 208 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 209 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 210 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 211 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 212 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 213 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 214 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 215 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 216 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 217 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 218 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 219 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 220 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 221 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 222 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 223 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 224 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 225 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 226 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 227 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 228 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 229 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 230 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 231 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 232 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 233 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 234 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 235 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 236 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 237 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 238 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 239 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 240 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 241 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 242 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 243 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 244 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 245 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 246 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 247 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 248 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 249 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 250 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 251 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 252 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 253 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 254 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 255 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 256 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 257 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 258 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 259 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 260 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 261 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 262 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 263 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 264 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 265 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 266 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 267 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 268 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 269 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 270 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 271 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 272 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 273 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 274 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 275 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 276 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 277 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 278 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 279 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 280 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 281 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 282 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 283 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 284 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 285 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 286 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 287 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 288 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 289 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 290 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 291 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 292 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 293 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 294 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 295 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 296 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 297 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 298 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 299 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 300 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 301 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 302 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 303 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 304 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 305 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 306 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 307 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 308 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 309 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 310 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 311 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 312 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 313 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 314 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 315 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 316 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 317 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 318 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 319 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 320 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 321 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 322 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 323 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 324 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 325 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 326 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 327 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 328 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 329 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 330 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 331 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 332 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 333 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 334 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 335 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 336 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 337 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 338 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 339 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 340 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 341 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 342 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 343 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 344 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 345 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 346 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 347 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 348 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 349 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 350 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 351 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 352 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 353 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 354 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 355 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 356 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 357 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 358 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 359 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 360 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 361 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 362 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 363 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 364 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 365 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 366 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 367 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 368 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 369 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 370 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 371 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 372 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 373 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 374 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 375 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 376 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 377 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 378 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 379 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 380 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 381 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 382 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 383 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 384 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 385 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 386 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 387 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 388 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 389 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 390 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 391 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 392 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 393 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 394 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 395 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 396 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 397 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 398 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 399 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 400 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 401 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 402 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 403 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 404 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 405 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 406 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 407 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 408 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 409 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 410 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 411 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 412 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 413 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 414 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 415 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 416 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 417 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 418 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 419 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 420 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 421 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 422 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 423 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 424 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 425 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 426 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 427 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 428 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 429 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 430 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 431 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 432 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 433 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 434 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 435 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 436 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 437 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 438 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 439 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 440 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 441 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 442 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 443 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 444 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 445 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 446 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 447 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 448 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 449 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 450 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 451 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 452 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 453 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 454 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 455 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 456 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 457 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 458 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 459 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 460 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 461 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 462 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 463 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 464 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 465 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 466 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 467 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 468 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 469 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 470 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 471 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 472 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 473 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 474 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 475 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 476 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 477 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 478 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 479 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 480 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 481 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 482 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 483 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 484 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 485 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 486 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 487 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 488 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 489 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 490 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 491 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 492 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 493 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 494 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 495 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 496 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 497 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 498 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 499 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 500 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 501 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 502 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 503 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 504 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 505 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 506 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 507 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 508 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 509 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 510 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 511 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 512 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 513 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 514 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 515 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 516 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 517 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 518 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 519 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 520 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 521 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 522 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 523 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 524 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 525 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 526 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 527 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 528 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 529 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 530 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 531 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 532 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 533 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 534 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 535 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 536 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 537 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 538 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 539 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 540 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 541 nsew signal input
flabel metal3 s 59200 53728 60000 53848 0 FreeSans 480 0 0 0 rst_o
port 542 nsew signal tristate
flabel metal3 s 59200 56448 60000 56568 0 FreeSans 480 0 0 0 start_o
port 543 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 544 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 544 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 545 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 545 nsew ground bidirectional
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wb_clk_i
port 546 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wb_rst_i
port 547 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 548 nsew signal tristate
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 549 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 550 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 551 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 552 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 553 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 554 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 555 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 556 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 557 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 558 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 559 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 560 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 561 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 562 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 563 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 564 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 565 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 566 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 567 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 568 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 569 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 570 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 571 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 572 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 573 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 574 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 575 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 576 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 577 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 578 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 579 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 580 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 581 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 582 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 583 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 584 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 585 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 586 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 587 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 588 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 589 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 590 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 591 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 592 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 593 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 594 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 595 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 596 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 597 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 598 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 599 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 600 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 601 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 602 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 603 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 604 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 605 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 606 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 607 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 608 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 609 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 610 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 611 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 612 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 613 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 614 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 615 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 616 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 617 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 618 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 619 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 620 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 621 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 622 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 623 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 624 nsew signal tristate
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 625 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 626 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 627 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 628 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 629 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 630 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 631 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 632 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 633 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 634 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 635 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 636 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 637 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 638 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 639 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 640 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 641 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 642 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 643 nsew signal tristate
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 644 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 645 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 646 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 647 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 648 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 649 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 650 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_we_i
port 651 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
