magic
tech sky130B
magscale 1 2
timestamp 1668103035
<< viali >>
rect 12909 57545 12943 57579
rect 14473 57545 14507 57579
rect 16865 57545 16899 57579
rect 17693 57545 17727 57579
rect 19441 57545 19475 57579
rect 20821 57545 20855 57579
rect 22385 57545 22419 57579
rect 24593 57545 24627 57579
rect 25513 57545 25547 57579
rect 27169 57545 27203 57579
rect 28641 57545 28675 57579
rect 30205 57545 30239 57579
rect 32321 57545 32355 57579
rect 33333 57545 33367 57579
rect 34897 57545 34931 57579
rect 36461 57545 36495 57579
rect 38025 57545 38059 57579
rect 40049 57545 40083 57579
rect 41153 57545 41187 57579
rect 42717 57545 42751 57579
rect 44281 57545 44315 57579
rect 45845 57545 45879 57579
rect 47777 57545 47811 57579
rect 48973 57545 49007 57579
rect 50537 57545 50571 57579
rect 52101 57545 52135 57579
rect 53665 57545 53699 57579
rect 55505 57545 55539 57579
rect 56793 57545 56827 57579
rect 58081 57545 58115 57579
rect 1869 57409 1903 57443
rect 3801 57409 3835 57443
rect 4997 57409 5031 57443
rect 6561 57409 6595 57443
rect 8125 57409 8159 57443
rect 9689 57409 9723 57443
rect 11529 57409 11563 57443
rect 13093 57409 13127 57443
rect 14657 57409 14691 57443
rect 16681 57409 16715 57443
rect 17509 57409 17543 57443
rect 19257 57409 19291 57443
rect 20637 57409 20671 57443
rect 22201 57409 22235 57443
rect 24409 57409 24443 57443
rect 25329 57409 25363 57443
rect 26985 57409 27019 57443
rect 28457 57409 28491 57443
rect 30021 57409 30055 57443
rect 32137 57409 32171 57443
rect 33149 57409 33183 57443
rect 34713 57409 34747 57443
rect 36277 57409 36311 57443
rect 37841 57409 37875 57443
rect 39865 57409 39899 57443
rect 40969 57409 41003 57443
rect 42533 57409 42567 57443
rect 44097 57409 44131 57443
rect 45661 57409 45695 57443
rect 47593 57409 47627 57443
rect 48789 57409 48823 57443
rect 50353 57409 50387 57443
rect 51917 57409 51951 57443
rect 53481 57409 53515 57443
rect 55321 57409 55355 57443
rect 56609 57409 56643 57443
rect 57897 57409 57931 57443
rect 56057 57205 56091 57239
rect 40785 57001 40819 57035
rect 57529 57001 57563 57035
rect 42349 56933 42383 56967
rect 58173 56797 58207 56831
rect 16129 56661 16163 56695
rect 28089 56661 28123 56695
rect 29561 56661 29595 56695
rect 45385 56661 45419 56695
rect 13737 56457 13771 56491
rect 14841 56457 14875 56491
rect 15945 56457 15979 56491
rect 16865 56457 16899 56491
rect 18153 56457 18187 56491
rect 18797 56457 18831 56491
rect 22293 56457 22327 56491
rect 23305 56457 23339 56491
rect 27813 56457 27847 56491
rect 30389 56457 30423 56491
rect 32321 56457 32355 56491
rect 33793 56457 33827 56491
rect 36001 56457 36035 56491
rect 43085 56457 43119 56491
rect 43729 56457 43763 56491
rect 45017 56457 45051 56491
rect 46305 56457 46339 56491
rect 21097 56389 21131 56423
rect 13921 56321 13955 56355
rect 15025 56321 15059 56355
rect 15761 56321 15795 56355
rect 16681 56321 16715 56355
rect 17325 56321 17359 56355
rect 17969 56321 18003 56355
rect 18613 56321 18647 56355
rect 19257 56321 19291 56355
rect 20913 56321 20947 56355
rect 22109 56321 22143 56355
rect 23121 56321 23155 56355
rect 23765 56321 23799 56355
rect 27629 56321 27663 56355
rect 28273 56321 28307 56355
rect 29193 56321 29227 56355
rect 30205 56321 30239 56355
rect 31401 56321 31435 56355
rect 32137 56321 32171 56355
rect 32781 56321 32815 56355
rect 33609 56321 33643 56355
rect 34253 56321 34287 56355
rect 35817 56321 35851 56355
rect 36461 56321 36495 56355
rect 42901 56321 42935 56355
rect 43545 56321 43579 56355
rect 44189 56321 44223 56355
rect 44833 56321 44867 56355
rect 45477 56321 45511 56355
rect 46121 56321 46155 56355
rect 46765 56321 46799 56355
rect 58173 56321 58207 56355
rect 17509 56185 17543 56219
rect 19441 56185 19475 56219
rect 28457 56185 28491 56219
rect 29377 56185 29411 56219
rect 44373 56185 44407 56219
rect 46949 56185 46983 56219
rect 20361 56117 20395 56151
rect 27077 56117 27111 56151
rect 30849 56117 30883 56151
rect 31585 56117 31619 56151
rect 45661 56117 45695 56151
rect 17877 55913 17911 55947
rect 21189 55913 21223 55947
rect 21005 55709 21039 55743
rect 27629 55709 27663 55743
rect 28273 55709 28307 55743
rect 18429 55641 18463 55675
rect 14197 55573 14231 55607
rect 15117 55573 15151 55607
rect 16589 55573 16623 55607
rect 17233 55573 17267 55607
rect 19257 55573 19291 55607
rect 20453 55573 20487 55607
rect 21925 55573 21959 55607
rect 27813 55573 27847 55607
rect 30021 55573 30055 55607
rect 42809 55573 42843 55607
rect 43453 55573 43487 55607
rect 44005 55573 44039 55607
rect 45017 55573 45051 55607
rect 46029 55573 46063 55607
rect 46673 55573 46707 55607
rect 58173 55097 58207 55131
rect 58173 53941 58207 53975
rect 58173 52445 58207 52479
rect 43177 51357 43211 51391
rect 43821 51357 43855 51391
rect 58173 51357 58207 51391
rect 43361 51221 43395 51255
rect 58173 49725 58207 49759
rect 58173 48501 58207 48535
rect 58173 47005 58207 47039
rect 58173 45917 58207 45951
rect 56333 45441 56367 45475
rect 56977 45441 57011 45475
rect 56517 45305 56551 45339
rect 58173 44217 58207 44251
rect 58173 43061 58207 43095
rect 15853 42517 15887 42551
rect 12265 42177 12299 42211
rect 12449 42177 12483 42211
rect 15025 42177 15059 42211
rect 15209 42177 15243 42211
rect 15301 42177 15335 42211
rect 15439 42177 15473 42211
rect 12633 41973 12667 42007
rect 15669 41973 15703 42007
rect 16589 41769 16623 41803
rect 11529 41701 11563 41735
rect 18705 41701 18739 41735
rect 14657 41633 14691 41667
rect 15761 41633 15795 41667
rect 12633 41565 12667 41599
rect 12725 41565 12759 41599
rect 12817 41565 12851 41599
rect 13001 41565 13035 41599
rect 15117 41565 15151 41599
rect 15301 41565 15335 41599
rect 15393 41565 15427 41599
rect 15485 41565 15519 41599
rect 19533 41565 19567 41599
rect 19625 41565 19659 41599
rect 19717 41565 19751 41599
rect 19901 41565 19935 41599
rect 58173 41565 58207 41599
rect 11713 41497 11747 41531
rect 11897 41497 11931 41531
rect 13553 41497 13587 41531
rect 14289 41497 14323 41531
rect 14473 41497 14507 41531
rect 16221 41497 16255 41531
rect 16405 41497 16439 41531
rect 17141 41497 17175 41531
rect 9689 41429 9723 41463
rect 12357 41429 12391 41463
rect 19257 41429 19291 41463
rect 20453 41429 20487 41463
rect 10977 41225 11011 41259
rect 15945 41157 15979 41191
rect 19450 41157 19484 41191
rect 9229 41089 9263 41123
rect 9321 41089 9355 41123
rect 9413 41089 9447 41123
rect 9597 41089 9631 41123
rect 10241 41089 10275 41123
rect 10425 41089 10459 41123
rect 12613 41089 12647 41123
rect 12725 41089 12759 41123
rect 12822 41089 12856 41123
rect 13001 41089 13035 41123
rect 14749 41089 14783 41123
rect 14912 41089 14946 41123
rect 15025 41089 15059 41123
rect 15163 41089 15197 41123
rect 20361 41089 20395 41123
rect 20545 41089 20579 41123
rect 22569 41089 22603 41123
rect 22753 41089 22787 41123
rect 19717 41021 19751 41055
rect 13553 40953 13587 40987
rect 8953 40885 8987 40919
rect 10057 40885 10091 40919
rect 12357 40885 12391 40919
rect 15393 40885 15427 40919
rect 18337 40885 18371 40919
rect 20177 40885 20211 40919
rect 22937 40885 22971 40919
rect 23489 40885 23523 40919
rect 14933 40681 14967 40715
rect 18705 40681 18739 40715
rect 17877 40613 17911 40647
rect 13185 40545 13219 40579
rect 20729 40545 20763 40579
rect 4057 40477 4091 40511
rect 4166 40471 4200 40505
rect 4266 40477 4300 40511
rect 4445 40477 4479 40511
rect 6101 40477 6135 40511
rect 9965 40477 9999 40511
rect 10057 40477 10091 40511
rect 10149 40477 10183 40511
rect 10333 40477 10367 40511
rect 11161 40477 11195 40511
rect 13461 40477 13495 40511
rect 14565 40477 14599 40511
rect 15393 40477 15427 40511
rect 18521 40477 18555 40511
rect 19533 40477 19567 40511
rect 19625 40477 19659 40511
rect 19717 40477 19751 40511
rect 19901 40477 19935 40511
rect 22569 40477 22603 40511
rect 22753 40477 22787 40511
rect 22845 40477 22879 40511
rect 22937 40477 22971 40511
rect 27261 40477 27295 40511
rect 58173 40477 58207 40511
rect 4905 40409 4939 40443
rect 6346 40409 6380 40443
rect 10977 40409 11011 40443
rect 14749 40409 14783 40443
rect 15660 40409 15694 40443
rect 18337 40409 18371 40443
rect 20996 40409 21030 40443
rect 27506 40409 27540 40443
rect 3801 40341 3835 40375
rect 5641 40341 5675 40375
rect 7481 40341 7515 40375
rect 9689 40341 9723 40375
rect 10793 40341 10827 40375
rect 12081 40341 12115 40375
rect 16773 40341 16807 40375
rect 19257 40341 19291 40375
rect 22109 40341 22143 40375
rect 23213 40341 23247 40375
rect 23673 40341 23707 40375
rect 28641 40341 28675 40375
rect 3893 40137 3927 40171
rect 4353 40137 4387 40171
rect 5825 40137 5859 40171
rect 12909 40137 12943 40171
rect 14749 40137 14783 40171
rect 2780 40069 2814 40103
rect 4537 40069 4571 40103
rect 6377 40069 6411 40103
rect 6561 40069 6595 40103
rect 11796 40069 11830 40103
rect 15862 40069 15896 40103
rect 17969 40069 18003 40103
rect 20913 40069 20947 40103
rect 21097 40069 21131 40103
rect 28181 40069 28215 40103
rect 28365 40069 28399 40103
rect 4721 40001 4755 40035
rect 5205 40001 5239 40035
rect 5344 40007 5378 40041
rect 5460 40001 5494 40035
rect 5595 40001 5629 40035
rect 6745 40001 6779 40035
rect 7472 40001 7506 40035
rect 10057 40001 10091 40035
rect 10149 40001 10183 40035
rect 10241 40001 10275 40035
rect 10425 40001 10459 40035
rect 16129 40001 16163 40035
rect 22477 40001 22511 40035
rect 22661 40001 22695 40035
rect 22753 40001 22787 40035
rect 22845 40001 22879 40035
rect 24694 40001 24728 40035
rect 30573 40001 30607 40035
rect 30736 40007 30770 40041
rect 30849 40001 30883 40035
rect 30987 40001 31021 40035
rect 2513 39933 2547 39967
rect 7205 39933 7239 39967
rect 11529 39933 11563 39967
rect 23121 39933 23155 39967
rect 24961 39933 24995 39967
rect 8585 39797 8619 39831
rect 9781 39797 9815 39831
rect 10977 39797 11011 39831
rect 17417 39797 17451 39831
rect 19257 39797 19291 39831
rect 20269 39797 20303 39831
rect 21281 39797 21315 39831
rect 23581 39797 23615 39831
rect 27997 39797 28031 39831
rect 30021 39797 30055 39831
rect 31217 39797 31251 39831
rect 11253 39593 11287 39627
rect 15485 39593 15519 39627
rect 21373 39593 21407 39627
rect 6285 39457 6319 39491
rect 7573 39457 7607 39491
rect 31033 39457 31067 39491
rect 4445 39389 4479 39423
rect 6561 39389 6595 39423
rect 9137 39389 9171 39423
rect 9404 39389 9438 39423
rect 12366 39389 12400 39423
rect 12633 39389 12667 39423
rect 16865 39389 16899 39423
rect 19257 39389 19291 39423
rect 19524 39389 19558 39423
rect 21649 39389 21683 39423
rect 21741 39389 21775 39423
rect 21833 39389 21867 39423
rect 22017 39389 22051 39423
rect 23857 39389 23891 39423
rect 27169 39389 27203 39423
rect 31300 39389 31334 39423
rect 4712 39321 4746 39355
rect 16598 39321 16632 39355
rect 23590 39321 23624 39355
rect 27436 39321 27470 39355
rect 5825 39253 5859 39287
rect 10517 39253 10551 39287
rect 20637 39253 20671 39287
rect 22477 39253 22511 39287
rect 28549 39253 28583 39287
rect 29745 39253 29779 39287
rect 30389 39253 30423 39287
rect 32413 39253 32447 39287
rect 5181 39049 5215 39083
rect 12633 39049 12667 39083
rect 22845 39049 22879 39083
rect 27169 39049 27203 39083
rect 4721 38981 4755 39015
rect 9220 38981 9254 39015
rect 22477 38981 22511 39015
rect 32137 38981 32171 39015
rect 2953 38913 2987 38947
rect 3046 38913 3080 38947
rect 3162 38913 3196 38947
rect 3341 38913 3375 38947
rect 5457 38913 5491 38947
rect 5546 38913 5580 38947
rect 5641 38913 5675 38947
rect 5825 38913 5859 38947
rect 6561 38913 6595 38947
rect 6745 38913 6779 38947
rect 8953 38913 8987 38947
rect 12449 38913 12483 38947
rect 13461 38913 13495 38947
rect 22661 38913 22695 38947
rect 25237 38913 25271 38947
rect 25421 38913 25455 38947
rect 25513 38913 25547 38947
rect 25605 38913 25639 38947
rect 27445 38913 27479 38947
rect 27537 38913 27571 38947
rect 27629 38913 27663 38947
rect 27813 38913 27847 38947
rect 28273 38913 28307 38947
rect 30737 38913 30771 38947
rect 30846 38913 30880 38947
rect 30941 38916 30975 38950
rect 31125 38913 31159 38947
rect 32321 38913 32355 38947
rect 32505 38913 32539 38947
rect 6377 38845 6411 38879
rect 7481 38845 7515 38879
rect 7757 38845 7791 38879
rect 13185 38845 13219 38879
rect 26341 38845 26375 38879
rect 3893 38777 3927 38811
rect 58173 38777 58207 38811
rect 2697 38709 2731 38743
rect 10333 38709 10367 38743
rect 21925 38709 21959 38743
rect 24777 38709 24811 38743
rect 25881 38709 25915 38743
rect 29561 38709 29595 38743
rect 30481 38709 30515 38743
rect 6561 38505 6595 38539
rect 7941 38505 7975 38539
rect 9137 38505 9171 38539
rect 27537 38505 27571 38539
rect 14657 38437 14691 38471
rect 19901 38437 19935 38471
rect 30205 38369 30239 38403
rect 1869 38301 1903 38335
rect 2136 38301 2170 38335
rect 8125 38301 8159 38335
rect 9321 38301 9355 38335
rect 14105 38301 14139 38335
rect 14473 38301 14507 38335
rect 17601 38301 17635 38335
rect 17694 38301 17728 38335
rect 17969 38301 18003 38335
rect 18107 38301 18141 38335
rect 19257 38301 19291 38335
rect 19350 38301 19384 38335
rect 19722 38301 19756 38335
rect 24593 38301 24627 38335
rect 24777 38301 24811 38335
rect 24869 38301 24903 38335
rect 24961 38301 24995 38335
rect 25697 38301 25731 38335
rect 25964 38301 25998 38335
rect 27813 38301 27847 38335
rect 27902 38301 27936 38335
rect 27997 38301 28031 38335
rect 28181 38301 28215 38335
rect 29009 38301 29043 38335
rect 30472 38301 30506 38335
rect 32689 38301 32723 38335
rect 5273 38233 5307 38267
rect 9505 38233 9539 38267
rect 14289 38233 14323 38267
rect 14381 38233 14415 38267
rect 17877 38233 17911 38267
rect 19533 38233 19567 38267
rect 19625 38233 19659 38267
rect 20545 38233 20579 38267
rect 20729 38233 20763 38267
rect 28641 38233 28675 38267
rect 28825 38233 28859 38267
rect 32956 38233 32990 38267
rect 3249 38165 3283 38199
rect 18245 38165 18279 38199
rect 20361 38165 20395 38199
rect 23857 38165 23891 38199
rect 25237 38165 25271 38199
rect 27077 38165 27111 38199
rect 31585 38165 31619 38199
rect 34069 38165 34103 38199
rect 4629 37961 4663 37995
rect 14381 37961 14415 37995
rect 26065 37961 26099 37995
rect 31125 37961 31159 37995
rect 33057 37961 33091 37995
rect 4169 37893 4203 37927
rect 4997 37893 5031 37927
rect 11805 37893 11839 37927
rect 14013 37893 14047 37927
rect 14105 37893 14139 37927
rect 21097 37893 21131 37927
rect 26433 37893 26467 37927
rect 31493 37893 31527 37927
rect 2927 37825 2961 37859
rect 3046 37831 3080 37865
rect 3162 37825 3196 37859
rect 3341 37825 3375 37859
rect 3985 37825 4019 37859
rect 4813 37825 4847 37859
rect 11529 37825 11563 37859
rect 11713 37825 11747 37859
rect 11897 37825 11931 37859
rect 13829 37825 13863 37859
rect 14197 37825 14231 37859
rect 18153 37825 18187 37859
rect 18409 37825 18443 37859
rect 19993 37825 20027 37859
rect 20177 37825 20211 37859
rect 20269 37825 20303 37859
rect 20361 37825 20395 37859
rect 25338 37825 25372 37859
rect 25605 37825 25639 37859
rect 26249 37825 26283 37859
rect 29357 37825 29391 37859
rect 31309 37825 31343 37859
rect 32413 37825 32447 37859
rect 32597 37825 32631 37859
rect 32689 37825 32723 37859
rect 32781 37825 32815 37859
rect 3801 37757 3835 37791
rect 29101 37757 29135 37791
rect 2697 37621 2731 37655
rect 7205 37621 7239 37655
rect 12081 37621 12115 37655
rect 19533 37621 19567 37655
rect 20637 37621 20671 37655
rect 24225 37621 24259 37655
rect 27353 37621 27387 37655
rect 30481 37621 30515 37655
rect 33517 37621 33551 37655
rect 34161 37621 34195 37655
rect 58173 37621 58207 37655
rect 3801 37417 3835 37451
rect 18061 37417 18095 37451
rect 18521 37417 18555 37451
rect 20453 37417 20487 37451
rect 24685 37417 24719 37451
rect 30481 37417 30515 37451
rect 33057 37417 33091 37451
rect 16681 37349 16715 37383
rect 1869 37281 1903 37315
rect 14749 37281 14783 37315
rect 31493 37281 31527 37315
rect 31723 37281 31757 37315
rect 2136 37213 2170 37247
rect 6009 37213 6043 37247
rect 7849 37213 7883 37247
rect 8125 37213 8159 37247
rect 8217 37213 8251 37247
rect 15301 37213 15335 37247
rect 17417 37213 17451 37247
rect 17601 37213 17635 37247
rect 17693 37213 17727 37247
rect 17785 37213 17819 37247
rect 19257 37213 19291 37247
rect 19350 37213 19384 37247
rect 19625 37213 19659 37247
rect 19722 37213 19756 37247
rect 21566 37213 21600 37247
rect 21833 37213 21867 37247
rect 32689 37213 32723 37247
rect 33517 37213 33551 37247
rect 33701 37213 33735 37247
rect 33793 37213 33827 37247
rect 33931 37213 33965 37247
rect 36093 37213 36127 37247
rect 6276 37145 6310 37179
rect 8033 37145 8067 37179
rect 11345 37145 11379 37179
rect 11805 37145 11839 37179
rect 14381 37145 14415 37179
rect 14565 37145 14599 37179
rect 15568 37145 15602 37179
rect 19533 37145 19567 37179
rect 24869 37145 24903 37179
rect 25053 37145 25087 37179
rect 32873 37145 32907 37179
rect 34161 37145 34195 37179
rect 35826 37145 35860 37179
rect 3249 37077 3283 37111
rect 7389 37077 7423 37111
rect 8401 37077 8435 37111
rect 13277 37077 13311 37111
rect 19901 37077 19935 37111
rect 23397 37077 23431 37111
rect 34713 37077 34747 37111
rect 12909 36873 12943 36907
rect 15485 36873 15519 36907
rect 18061 36873 18095 36907
rect 19901 36873 19935 36907
rect 6653 36805 6687 36839
rect 7573 36805 7607 36839
rect 16865 36805 16899 36839
rect 17877 36805 17911 36839
rect 23029 36805 23063 36839
rect 6377 36737 6411 36771
rect 6561 36737 6595 36771
rect 6745 36737 6779 36771
rect 7389 36737 7423 36771
rect 10793 36737 10827 36771
rect 12173 36737 12207 36771
rect 13001 36737 13035 36771
rect 13820 36737 13854 36771
rect 15761 36737 15795 36771
rect 15853 36737 15887 36771
rect 15945 36737 15979 36771
rect 16129 36737 16163 36771
rect 17049 36737 17083 36771
rect 17693 36737 17727 36771
rect 22937 36737 22971 36771
rect 23121 36737 23155 36771
rect 23305 36737 23339 36771
rect 23765 36737 23799 36771
rect 25973 36737 26007 36771
rect 34253 36737 34287 36771
rect 36470 36737 36504 36771
rect 10517 36669 10551 36703
rect 13553 36669 13587 36703
rect 16681 36669 16715 36703
rect 36737 36669 36771 36703
rect 14933 36601 14967 36635
rect 6929 36533 6963 36567
rect 7757 36533 7791 36567
rect 12265 36533 12299 36567
rect 22293 36533 22327 36567
rect 22753 36533 22787 36567
rect 25053 36533 25087 36567
rect 27997 36533 28031 36567
rect 32965 36533 32999 36567
rect 34805 36533 34839 36567
rect 35357 36533 35391 36567
rect 5181 36329 5215 36363
rect 7113 36329 7147 36363
rect 14105 36329 14139 36363
rect 16313 36329 16347 36363
rect 33793 36329 33827 36363
rect 35357 36329 35391 36363
rect 27905 36261 27939 36295
rect 3801 36193 3835 36227
rect 12725 36193 12759 36227
rect 15209 36193 15243 36227
rect 29009 36193 29043 36227
rect 7389 36125 7423 36159
rect 7478 36125 7512 36159
rect 7573 36122 7607 36156
rect 7757 36125 7791 36159
rect 9413 36125 9447 36159
rect 10057 36125 10091 36159
rect 12449 36125 12483 36159
rect 14381 36125 14415 36159
rect 14473 36125 14507 36159
rect 14565 36125 14599 36159
rect 14749 36125 14783 36159
rect 22201 36125 22235 36159
rect 22293 36125 22327 36159
rect 22569 36125 22603 36159
rect 24409 36125 24443 36159
rect 28365 36125 28399 36159
rect 28549 36125 28583 36159
rect 28641 36125 28675 36159
rect 28733 36125 28767 36159
rect 29745 36125 29779 36159
rect 32413 36125 32447 36159
rect 34713 36125 34747 36159
rect 34897 36125 34931 36159
rect 34989 36125 35023 36159
rect 35081 36125 35115 36159
rect 58173 36125 58207 36159
rect 4068 36057 4102 36091
rect 8309 36057 8343 36091
rect 10324 36057 10358 36091
rect 22385 36057 22419 36091
rect 29561 36057 29595 36091
rect 29929 36057 29963 36091
rect 33425 36057 33459 36091
rect 33609 36057 33643 36091
rect 9597 35989 9631 36023
rect 11437 35989 11471 36023
rect 22017 35989 22051 36023
rect 23121 35989 23155 36023
rect 23673 35989 23707 36023
rect 27077 35989 27111 36023
rect 13369 35785 13403 35819
rect 35081 35785 35115 35819
rect 4997 35717 5031 35751
rect 11897 35717 11931 35751
rect 12357 35717 12391 35751
rect 12541 35717 12575 35751
rect 4813 35649 4847 35683
rect 8309 35649 8343 35683
rect 9873 35649 9907 35683
rect 11713 35649 11747 35683
rect 13277 35649 13311 35683
rect 14473 35649 14507 35683
rect 17233 35649 17267 35683
rect 17325 35649 17359 35683
rect 17417 35649 17451 35683
rect 17601 35649 17635 35683
rect 22661 35649 22695 35683
rect 22753 35649 22787 35683
rect 22845 35649 22879 35683
rect 23029 35649 23063 35683
rect 24225 35649 24259 35683
rect 24481 35649 24515 35683
rect 27353 35649 27387 35683
rect 27620 35649 27654 35683
rect 30113 35649 30147 35683
rect 30297 35649 30331 35683
rect 30389 35649 30423 35683
rect 30481 35649 30515 35683
rect 34713 35649 34747 35683
rect 34897 35649 34931 35683
rect 8033 35581 8067 35615
rect 9597 35581 9631 35615
rect 10977 35581 11011 35615
rect 23489 35581 23523 35615
rect 32137 35581 32171 35615
rect 32413 35581 32447 35615
rect 11529 35513 11563 35547
rect 13921 35513 13955 35547
rect 18061 35513 18095 35547
rect 29561 35513 29595 35547
rect 5181 35445 5215 35479
rect 12725 35445 12759 35479
rect 16957 35445 16991 35479
rect 22477 35445 22511 35479
rect 25605 35445 25639 35479
rect 28733 35445 28767 35479
rect 30757 35445 30791 35479
rect 31493 35445 31527 35479
rect 4721 35241 4755 35275
rect 11805 35241 11839 35275
rect 21097 35241 21131 35275
rect 25789 35241 25823 35275
rect 27445 35241 27479 35275
rect 8125 35173 8159 35207
rect 10425 35105 10459 35139
rect 22753 35105 22787 35139
rect 24409 35105 24443 35139
rect 32045 35105 32079 35139
rect 4997 35037 5031 35071
rect 5089 35037 5123 35071
rect 5181 35037 5215 35071
rect 5365 35037 5399 35071
rect 6101 35037 6135 35071
rect 8309 35037 8343 35071
rect 9321 35037 9355 35071
rect 9505 35037 9539 35071
rect 9597 35037 9631 35071
rect 9689 35037 9723 35071
rect 13001 35037 13035 35071
rect 13277 35037 13311 35071
rect 13369 35037 13403 35071
rect 17141 35037 17175 35071
rect 17397 35037 17431 35071
rect 19901 35037 19935 35071
rect 21925 35037 21959 35071
rect 22017 35037 22051 35071
rect 22109 35037 22143 35071
rect 22293 35037 22327 35071
rect 26433 35037 26467 35071
rect 27721 35037 27755 35071
rect 27810 35034 27844 35068
rect 27905 35037 27939 35071
rect 28089 35037 28123 35071
rect 28733 35037 28767 35071
rect 31778 35037 31812 35071
rect 32505 35037 32539 35071
rect 32781 35037 32815 35071
rect 58173 35037 58207 35071
rect 6368 34969 6402 35003
rect 9965 34969 9999 35003
rect 10670 34969 10704 35003
rect 13185 34969 13219 35003
rect 19717 34969 19751 35003
rect 22937 34969 22971 35003
rect 23121 34969 23155 35003
rect 24654 34969 24688 35003
rect 26617 34969 26651 35003
rect 28549 34969 28583 35003
rect 28917 34969 28951 35003
rect 7481 34901 7515 34935
rect 13553 34901 13587 34935
rect 18521 34901 18555 34935
rect 20085 34901 20119 34935
rect 21649 34901 21683 34935
rect 23857 34901 23891 34935
rect 26249 34901 26283 34935
rect 30113 34901 30147 34935
rect 30665 34901 30699 34935
rect 33885 34901 33919 34935
rect 3893 34697 3927 34731
rect 7021 34697 7055 34731
rect 10333 34697 10367 34731
rect 12817 34697 12851 34731
rect 17325 34697 17359 34731
rect 19901 34697 19935 34731
rect 23213 34697 23247 34731
rect 24501 34697 24535 34731
rect 27077 34697 27111 34731
rect 27629 34697 27663 34731
rect 29929 34697 29963 34731
rect 32321 34697 32355 34731
rect 4537 34629 4571 34663
rect 8217 34629 8251 34663
rect 12541 34629 12575 34663
rect 17509 34629 17543 34663
rect 19073 34629 19107 34663
rect 19162 34629 19196 34663
rect 22078 34629 22112 34663
rect 24041 34629 24075 34663
rect 25789 34629 25823 34663
rect 25973 34629 26007 34663
rect 29745 34629 29779 34663
rect 33333 34629 33367 34663
rect 33517 34629 33551 34663
rect 2780 34561 2814 34595
rect 4721 34561 4755 34595
rect 7297 34561 7331 34595
rect 7389 34561 7423 34595
rect 7481 34561 7515 34595
rect 7665 34561 7699 34595
rect 10609 34561 10643 34595
rect 10701 34561 10735 34595
rect 10793 34561 10827 34595
rect 10977 34561 11011 34595
rect 12265 34561 12299 34595
rect 12449 34561 12483 34595
rect 12633 34561 12667 34595
rect 17693 34561 17727 34595
rect 18797 34561 18831 34595
rect 18890 34561 18924 34595
rect 19281 34561 19315 34595
rect 21014 34561 21048 34595
rect 21281 34561 21315 34595
rect 21833 34561 21867 34595
rect 24731 34561 24765 34595
rect 24869 34561 24903 34595
rect 24961 34561 24995 34595
rect 25145 34561 25179 34595
rect 29561 34561 29595 34595
rect 30941 34561 30975 34595
rect 32137 34561 32171 34595
rect 33149 34561 33183 34595
rect 33977 34561 34011 34595
rect 34161 34561 34195 34595
rect 34256 34561 34290 34595
rect 34345 34561 34379 34595
rect 2513 34493 2547 34527
rect 5549 34493 5583 34527
rect 25605 34493 25639 34527
rect 31217 34493 31251 34527
rect 34621 34493 34655 34527
rect 19441 34425 19475 34459
rect 4353 34357 4387 34391
rect 11621 34357 11655 34391
rect 16773 34357 16807 34391
rect 2605 34153 2639 34187
rect 7389 34153 7423 34187
rect 20361 34153 20395 34187
rect 24409 34153 24443 34187
rect 33057 34153 33091 34187
rect 7849 34085 7883 34119
rect 29745 34085 29779 34119
rect 14381 34017 14415 34051
rect 16773 34017 16807 34051
rect 31769 34017 31803 34051
rect 2881 33949 2915 33983
rect 2973 33949 3007 33983
rect 3065 33949 3099 33983
rect 3249 33949 3283 33983
rect 4077 33949 4111 33983
rect 4169 33949 4203 33983
rect 4261 33949 4295 33983
rect 4445 33949 4479 33983
rect 5549 33949 5583 33983
rect 7205 33949 7239 33983
rect 8953 33949 8987 33983
rect 9046 33949 9080 33983
rect 9321 33949 9355 33983
rect 9459 33949 9493 33983
rect 14105 33949 14139 33983
rect 15945 33949 15979 33983
rect 16037 33949 16071 33983
rect 16129 33949 16163 33983
rect 16313 33949 16347 33983
rect 17141 33949 17175 33983
rect 18705 33949 18739 33983
rect 19717 33949 19751 33983
rect 19901 33949 19935 33983
rect 19993 33949 20027 33983
rect 20131 33949 20165 33983
rect 20821 33949 20855 33983
rect 23765 33949 23799 33983
rect 24639 33949 24673 33983
rect 24777 33949 24811 33983
rect 24869 33949 24903 33983
rect 25053 33949 25087 33983
rect 26709 33949 26743 33983
rect 27537 33949 27571 33983
rect 27626 33943 27660 33977
rect 27726 33949 27760 33983
rect 27905 33949 27939 33983
rect 30527 33949 30561 33983
rect 30665 33949 30699 33983
rect 30757 33949 30791 33983
rect 30941 33949 30975 33983
rect 33517 33949 33551 33983
rect 33701 33949 33735 33983
rect 33793 33949 33827 33983
rect 33885 33949 33919 33983
rect 36093 33949 36127 33983
rect 38485 33949 38519 33983
rect 2145 33881 2179 33915
rect 7021 33881 7055 33915
rect 9229 33881 9263 33915
rect 16957 33881 16991 33915
rect 17969 33881 18003 33915
rect 18521 33881 18555 33915
rect 31401 33881 31435 33915
rect 31585 33881 31619 33915
rect 34161 33881 34195 33915
rect 35826 33881 35860 33915
rect 36921 33881 36955 33915
rect 3801 33813 3835 33847
rect 4997 33813 5031 33847
rect 9597 33813 9631 33847
rect 11161 33813 11195 33847
rect 15669 33813 15703 33847
rect 27261 33813 27295 33847
rect 30297 33813 30331 33847
rect 34713 33813 34747 33847
rect 4353 33609 4387 33643
rect 6745 33609 6779 33643
rect 12633 33609 12667 33643
rect 15209 33609 15243 33643
rect 19717 33609 19751 33643
rect 30205 33609 30239 33643
rect 34069 33609 34103 33643
rect 34805 33609 34839 33643
rect 2780 33541 2814 33575
rect 17049 33541 17083 33575
rect 27414 33541 27448 33575
rect 35918 33541 35952 33575
rect 4537 33473 4571 33507
rect 4721 33473 4755 33507
rect 12725 33473 12759 33507
rect 13277 33473 13311 33507
rect 13544 33473 13578 33507
rect 15301 33473 15335 33507
rect 16681 33473 16715 33507
rect 16829 33473 16863 33507
rect 16957 33473 16991 33507
rect 17165 33473 17199 33507
rect 18521 33473 18555 33507
rect 18705 33473 18739 33507
rect 24685 33473 24719 33507
rect 24869 33473 24903 33507
rect 24961 33473 24995 33507
rect 25053 33473 25087 33507
rect 30021 33473 30055 33507
rect 33701 33473 33735 33507
rect 33885 33473 33919 33507
rect 2513 33405 2547 33439
rect 27169 33405 27203 33439
rect 32413 33405 32447 33439
rect 32689 33405 32723 33439
rect 36185 33405 36219 33439
rect 3893 33337 3927 33371
rect 58173 33337 58207 33371
rect 7941 33269 7975 33303
rect 14657 33269 14691 33303
rect 17325 33269 17359 33303
rect 18337 33269 18371 33303
rect 19257 33269 19291 33303
rect 24041 33269 24075 33303
rect 25329 33269 25363 33303
rect 25789 33269 25823 33303
rect 28549 33269 28583 33303
rect 29561 33269 29595 33303
rect 37289 33269 37323 33303
rect 3893 33065 3927 33099
rect 8309 33065 8343 33099
rect 13553 33065 13587 33099
rect 16957 33065 16991 33099
rect 27813 33065 27847 33099
rect 31217 33065 31251 33099
rect 20637 32997 20671 33031
rect 14381 32929 14415 32963
rect 24685 32929 24719 32963
rect 4905 32861 4939 32895
rect 7389 32861 7423 32895
rect 7481 32861 7515 32895
rect 7573 32861 7607 32895
rect 7757 32861 7791 32895
rect 10241 32861 10275 32895
rect 12909 32861 12943 32895
rect 13093 32861 13127 32895
rect 13185 32861 13219 32895
rect 13277 32861 13311 32895
rect 14105 32861 14139 32895
rect 15577 32861 15611 32895
rect 18067 32861 18101 32895
rect 18245 32861 18279 32895
rect 18337 32861 18371 32895
rect 18429 32861 18463 32895
rect 19257 32861 19291 32895
rect 24409 32861 24443 32895
rect 27997 32861 28031 32895
rect 29837 32861 29871 32895
rect 6653 32793 6687 32827
rect 12449 32793 12483 32827
rect 15822 32793 15856 32827
rect 18705 32793 18739 32827
rect 19502 32793 19536 32827
rect 28181 32793 28215 32827
rect 30104 32793 30138 32827
rect 32137 32793 32171 32827
rect 32321 32793 32355 32827
rect 7113 32725 7147 32759
rect 10333 32725 10367 32759
rect 21833 32725 21867 32759
rect 23857 32725 23891 32759
rect 32505 32725 32539 32759
rect 5181 32521 5215 32555
rect 5825 32521 5859 32555
rect 6469 32521 6503 32555
rect 8769 32521 8803 32555
rect 13737 32521 13771 32555
rect 18889 32521 18923 32555
rect 21189 32521 21223 32555
rect 22109 32521 22143 32555
rect 24501 32521 24535 32555
rect 24961 32521 24995 32555
rect 28733 32521 28767 32555
rect 29745 32521 29779 32555
rect 8953 32453 8987 32487
rect 12909 32453 12943 32487
rect 13921 32453 13955 32487
rect 17049 32453 17083 32487
rect 18981 32453 19015 32487
rect 19625 32453 19659 32487
rect 22753 32453 22787 32487
rect 24317 32453 24351 32487
rect 26074 32453 26108 32487
rect 27997 32453 28031 32487
rect 29009 32453 29043 32487
rect 30573 32453 30607 32487
rect 7196 32385 7230 32419
rect 9137 32385 9171 32419
rect 12725 32385 12759 32419
rect 14105 32385 14139 32419
rect 16865 32385 16899 32419
rect 17785 32385 17819 32419
rect 21925 32385 21959 32419
rect 23397 32385 23431 32419
rect 24133 32385 24167 32419
rect 27905 32385 27939 32419
rect 28089 32385 28123 32419
rect 28273 32385 28307 32419
rect 28917 32385 28951 32419
rect 29101 32385 29135 32419
rect 29285 32385 29319 32419
rect 33710 32385 33744 32419
rect 33977 32385 34011 32419
rect 37473 32385 37507 32419
rect 37729 32385 37763 32419
rect 6929 32317 6963 32351
rect 10517 32317 10551 32351
rect 10793 32317 10827 32351
rect 17509 32317 17543 32351
rect 26341 32317 26375 32351
rect 8309 32249 8343 32283
rect 23581 32249 23615 32283
rect 13093 32181 13127 32215
rect 27721 32181 27755 32215
rect 30481 32181 30515 32215
rect 32597 32181 32631 32215
rect 35909 32181 35943 32215
rect 38853 32181 38887 32215
rect 58173 32181 58207 32215
rect 22937 31977 22971 32011
rect 23673 31977 23707 32011
rect 30021 31977 30055 32011
rect 32873 31977 32907 32011
rect 36645 31977 36679 32011
rect 11897 31909 11931 31943
rect 22155 31909 22189 31943
rect 30757 31909 30791 31943
rect 8125 31841 8159 31875
rect 9597 31841 9631 31875
rect 16405 31841 16439 31875
rect 22385 31841 22419 31875
rect 27169 31841 27203 31875
rect 35541 31841 35575 31875
rect 1869 31773 1903 31807
rect 4997 31773 5031 31807
rect 5181 31773 5215 31807
rect 5273 31773 5307 31807
rect 5365 31773 5399 31807
rect 6469 31773 6503 31807
rect 6561 31773 6595 31807
rect 6653 31773 6687 31807
rect 6837 31773 6871 31807
rect 8401 31773 8435 31807
rect 9864 31773 9898 31807
rect 13277 31773 13311 31807
rect 16957 31773 16991 31807
rect 21005 31773 21039 31807
rect 23489 31773 23523 31807
rect 28825 31773 28859 31807
rect 30205 31773 30239 31807
rect 30941 31773 30975 31807
rect 31033 31773 31067 31807
rect 31309 31773 31343 31807
rect 32229 31773 32263 31807
rect 32413 31773 32447 31807
rect 32524 31773 32558 31807
rect 32617 31773 32651 31807
rect 35357 31773 35391 31807
rect 36001 31773 36035 31807
rect 36185 31773 36219 31807
rect 36277 31773 36311 31807
rect 36389 31773 36423 31807
rect 2136 31705 2170 31739
rect 13010 31705 13044 31739
rect 31125 31705 31159 31739
rect 35173 31705 35207 31739
rect 3249 31637 3283 31671
rect 5641 31637 5675 31671
rect 6193 31637 6227 31671
rect 10977 31637 11011 31671
rect 14197 31637 14231 31671
rect 18245 31637 18279 31671
rect 2145 31433 2179 31467
rect 5457 31433 5491 31467
rect 13093 31433 13127 31467
rect 17693 31433 17727 31467
rect 24225 31433 24259 31467
rect 35449 31433 35483 31467
rect 5641 31365 5675 31399
rect 6622 31365 6656 31399
rect 12357 31365 12391 31399
rect 14933 31365 14967 31399
rect 15853 31365 15887 31399
rect 16037 31365 16071 31399
rect 23029 31365 23063 31399
rect 28181 31365 28215 31399
rect 30297 31365 30331 31399
rect 31125 31365 31159 31399
rect 31217 31365 31251 31399
rect 35081 31365 35115 31399
rect 36553 31365 36587 31399
rect 38270 31365 38304 31399
rect 2401 31297 2435 31331
rect 2513 31297 2547 31331
rect 2610 31300 2644 31334
rect 2789 31297 2823 31331
rect 3433 31297 3467 31331
rect 3617 31297 3651 31331
rect 5825 31297 5859 31331
rect 10425 31297 10459 31331
rect 10609 31297 10643 31331
rect 12081 31297 12115 31331
rect 12265 31297 12299 31331
rect 12449 31297 12483 31331
rect 13369 31297 13403 31331
rect 13461 31297 13495 31331
rect 13553 31297 13587 31331
rect 13737 31297 13771 31331
rect 14565 31297 14599 31331
rect 14658 31297 14692 31331
rect 14841 31297 14875 31331
rect 15071 31297 15105 31331
rect 21097 31297 21131 31331
rect 22201 31297 22235 31331
rect 22293 31297 22327 31331
rect 22385 31297 22419 31331
rect 22569 31297 22603 31331
rect 23213 31297 23247 31331
rect 24041 31297 24075 31331
rect 27997 31297 28031 31331
rect 28641 31297 28675 31331
rect 31033 31297 31067 31331
rect 31401 31297 31435 31331
rect 35265 31297 35299 31331
rect 35909 31297 35943 31331
rect 36093 31297 36127 31331
rect 36185 31297 36219 31331
rect 36277 31297 36311 31331
rect 37289 31297 37323 31331
rect 38025 31297 38059 31331
rect 3249 31229 3283 31263
rect 6377 31229 6411 31263
rect 9689 31229 9723 31263
rect 9965 31229 9999 31263
rect 20821 31229 20855 31263
rect 23397 31229 23431 31263
rect 15209 31161 15243 31195
rect 27261 31161 27295 31195
rect 7757 31093 7791 31127
rect 8309 31093 8343 31127
rect 10793 31093 10827 31127
rect 12633 31093 12667 31127
rect 15669 31093 15703 31127
rect 19165 31093 19199 31127
rect 19809 31093 19843 31127
rect 21925 31093 21959 31127
rect 24777 31093 24811 31127
rect 27813 31093 27847 31127
rect 30849 31093 30883 31127
rect 32229 31093 32263 31127
rect 39405 31093 39439 31127
rect 7205 30889 7239 30923
rect 10885 30889 10919 30923
rect 12725 30889 12759 30923
rect 22937 30889 22971 30923
rect 23673 30889 23707 30923
rect 27813 30889 27847 30923
rect 35265 30889 35299 30923
rect 14105 30821 14139 30855
rect 16129 30821 16163 30855
rect 5365 30753 5399 30787
rect 14749 30753 14783 30787
rect 19257 30753 19291 30787
rect 24685 30753 24719 30787
rect 30665 30753 30699 30787
rect 37933 30753 37967 30787
rect 5632 30685 5666 30719
rect 7573 30685 7607 30719
rect 12173 30685 12207 30719
rect 18337 30685 18371 30719
rect 18429 30685 18463 30719
rect 18521 30685 18555 30719
rect 18705 30685 18739 30719
rect 21557 30685 21591 30719
rect 23857 30685 23891 30719
rect 24409 30685 24443 30719
rect 27077 30685 27111 30719
rect 28549 30685 28583 30719
rect 28641 30685 28675 30719
rect 28733 30685 28767 30719
rect 28917 30685 28951 30719
rect 30941 30685 30975 30719
rect 31401 30685 31435 30719
rect 31585 30685 31619 30719
rect 33149 30685 33183 30719
rect 33241 30685 33275 30719
rect 33517 30685 33551 30719
rect 35817 30685 35851 30719
rect 36001 30685 36035 30719
rect 36093 30685 36127 30719
rect 36185 30685 36219 30719
rect 58173 30685 58207 30719
rect 7389 30617 7423 30651
rect 14994 30617 15028 30651
rect 19524 30617 19558 30651
rect 21824 30617 21858 30651
rect 26810 30617 26844 30651
rect 33333 30617 33367 30651
rect 36461 30617 36495 30651
rect 38178 30617 38212 30651
rect 2881 30549 2915 30583
rect 6745 30549 6779 30583
rect 17509 30549 17543 30583
rect 18061 30549 18095 30583
rect 20637 30549 20671 30583
rect 25697 30549 25731 30583
rect 28273 30549 28307 30583
rect 31769 30549 31803 30583
rect 32965 30549 32999 30583
rect 39313 30549 39347 30583
rect 14749 30345 14783 30379
rect 19809 30345 19843 30379
rect 29469 30345 29503 30379
rect 35909 30345 35943 30379
rect 9873 30277 9907 30311
rect 11529 30277 11563 30311
rect 12081 30277 12115 30311
rect 18214 30277 18248 30311
rect 21189 30277 21223 30311
rect 22477 30277 22511 30311
rect 23857 30277 23891 30311
rect 25237 30277 25271 30311
rect 26985 30277 27019 30311
rect 30205 30277 30239 30311
rect 32597 30277 32631 30311
rect 32689 30277 32723 30311
rect 33701 30277 33735 30311
rect 35725 30277 35759 30311
rect 2421 30209 2455 30243
rect 2677 30209 2711 30243
rect 10149 30209 10183 30243
rect 10241 30209 10275 30243
rect 10333 30209 10367 30243
rect 10517 30209 10551 30243
rect 12265 30209 12299 30243
rect 15025 30209 15059 30243
rect 15117 30209 15151 30243
rect 15209 30209 15243 30243
rect 15393 30209 15427 30243
rect 16957 30209 16991 30243
rect 20085 30209 20119 30243
rect 20177 30209 20211 30243
rect 20269 30209 20303 30243
rect 20453 30209 20487 30243
rect 21005 30209 21039 30243
rect 22385 30209 22419 30243
rect 22569 30209 22603 30243
rect 22753 30209 22787 30243
rect 23673 30209 23707 30243
rect 24593 30209 24627 30243
rect 24777 30209 24811 30243
rect 24869 30209 24903 30243
rect 25007 30209 25041 30243
rect 25697 30209 25731 30243
rect 28089 30209 28123 30243
rect 28356 30209 28390 30243
rect 30113 30209 30147 30243
rect 30297 30209 30331 30243
rect 30481 30209 30515 30243
rect 32413 30209 32447 30243
rect 32781 30209 32815 30243
rect 33609 30209 33643 30243
rect 33793 30209 33827 30243
rect 33977 30209 34011 30243
rect 35541 30209 35575 30243
rect 12449 30141 12483 30175
rect 13001 30141 13035 30175
rect 16773 30141 16807 30175
rect 17969 30141 18003 30175
rect 24041 30141 24075 30175
rect 3801 30005 3835 30039
rect 9413 30005 9447 30039
rect 15945 30005 15979 30039
rect 17141 30005 17175 30039
rect 19349 30005 19383 30039
rect 22201 30005 22235 30039
rect 25881 30005 25915 30039
rect 29929 30005 29963 30039
rect 31217 30005 31251 30039
rect 32965 30005 32999 30039
rect 33425 30005 33459 30039
rect 36645 30005 36679 30039
rect 2237 29801 2271 29835
rect 8953 29801 8987 29835
rect 18705 29801 18739 29835
rect 20269 29801 20303 29835
rect 23857 29801 23891 29835
rect 29837 29801 29871 29835
rect 3801 29733 3835 29767
rect 24501 29733 24535 29767
rect 9321 29665 9355 29699
rect 26617 29665 26651 29699
rect 35817 29665 35851 29699
rect 2467 29597 2501 29631
rect 2605 29597 2639 29631
rect 2697 29597 2731 29631
rect 2881 29597 2915 29631
rect 4353 29597 4387 29631
rect 4629 29597 4663 29631
rect 4721 29597 4755 29631
rect 9137 29597 9171 29631
rect 10517 29597 10551 29631
rect 18521 29597 18555 29631
rect 21281 29597 21315 29631
rect 22385 29597 22419 29631
rect 22569 29597 22603 29631
rect 22753 29597 22787 29631
rect 24685 29597 24719 29631
rect 30849 29597 30883 29631
rect 31012 29597 31046 29631
rect 31125 29597 31159 29631
rect 31217 29597 31251 29631
rect 31953 29597 31987 29631
rect 34161 29597 34195 29631
rect 34713 29597 34747 29631
rect 35541 29597 35575 29631
rect 36829 29597 36863 29631
rect 37013 29597 37047 29631
rect 37105 29597 37139 29631
rect 37197 29597 37231 29631
rect 58173 29597 58207 29631
rect 4537 29529 4571 29563
rect 10784 29529 10818 29563
rect 17785 29529 17819 29563
rect 18337 29529 18371 29563
rect 19901 29529 19935 29563
rect 20085 29529 20119 29563
rect 22477 29529 22511 29563
rect 26350 29529 26384 29563
rect 31493 29529 31527 29563
rect 32198 29529 32232 29563
rect 33793 29529 33827 29563
rect 33977 29529 34011 29563
rect 4905 29461 4939 29495
rect 7849 29461 7883 29495
rect 10057 29461 10091 29495
rect 11897 29461 11931 29495
rect 16589 29461 16623 29495
rect 19349 29461 19383 29495
rect 20729 29461 20763 29495
rect 22201 29461 22235 29495
rect 23305 29461 23339 29495
rect 25237 29461 25271 29495
rect 30297 29461 30331 29495
rect 33333 29461 33367 29495
rect 34897 29461 34931 29495
rect 37473 29461 37507 29495
rect 10793 29257 10827 29291
rect 14381 29257 14415 29291
rect 25421 29257 25455 29291
rect 30389 29257 30423 29291
rect 30849 29257 30883 29291
rect 38117 29257 38151 29291
rect 4813 29189 4847 29223
rect 8217 29189 8251 29223
rect 8585 29189 8619 29223
rect 11713 29189 11747 29223
rect 15485 29189 15519 29223
rect 19901 29189 19935 29223
rect 19993 29189 20027 29223
rect 22569 29189 22603 29223
rect 23581 29189 23615 29223
rect 23765 29189 23799 29223
rect 35265 29189 35299 29223
rect 35633 29189 35667 29223
rect 39230 29189 39264 29223
rect 3065 29121 3099 29155
rect 3157 29121 3191 29155
rect 3254 29121 3288 29155
rect 3433 29121 3467 29155
rect 4537 29121 4571 29155
rect 4721 29121 4755 29155
rect 4905 29121 4939 29155
rect 7481 29121 7515 29155
rect 7665 29121 7699 29155
rect 8401 29121 8435 29155
rect 9275 29121 9309 29155
rect 9394 29127 9428 29161
rect 9505 29121 9539 29155
rect 9689 29121 9723 29155
rect 10149 29121 10183 29155
rect 10333 29121 10367 29155
rect 10425 29121 10459 29155
rect 10517 29121 10551 29155
rect 11897 29121 11931 29155
rect 15669 29121 15703 29155
rect 18061 29121 18095 29155
rect 18613 29121 18647 29155
rect 19717 29121 19751 29155
rect 20085 29121 20119 29155
rect 23397 29121 23431 29155
rect 24225 29121 24259 29155
rect 24388 29124 24422 29158
rect 24504 29124 24538 29158
rect 24593 29121 24627 29155
rect 25605 29121 25639 29155
rect 30205 29121 30239 29155
rect 30849 29121 30883 29155
rect 31033 29121 31067 29155
rect 33425 29121 33459 29155
rect 35449 29121 35483 29155
rect 36093 29121 36127 29155
rect 36277 29121 36311 29155
rect 36369 29121 36403 29155
rect 36507 29121 36541 29155
rect 11529 29053 11563 29087
rect 29469 29053 29503 29087
rect 30021 29053 30055 29087
rect 33701 29053 33735 29087
rect 39497 29053 39531 29087
rect 5089 28985 5123 29019
rect 7481 28985 7515 29019
rect 18797 28985 18831 29019
rect 20269 28985 20303 29019
rect 22753 28985 22787 29019
rect 24869 28985 24903 29019
rect 26157 28985 26191 29019
rect 36737 28985 36771 29019
rect 2789 28917 2823 28951
rect 3985 28917 4019 28951
rect 9045 28917 9079 28951
rect 13829 28917 13863 28951
rect 15853 28917 15887 28951
rect 16957 28917 16991 28951
rect 31493 28917 31527 28951
rect 37289 28917 37323 28951
rect 2605 28713 2639 28747
rect 3801 28713 3835 28747
rect 7573 28713 7607 28747
rect 10333 28713 10367 28747
rect 10793 28713 10827 28747
rect 15209 28713 15243 28747
rect 25053 28713 25087 28747
rect 36461 28713 36495 28747
rect 16589 28577 16623 28611
rect 30481 28577 30515 28611
rect 33517 28577 33551 28611
rect 2789 28509 2823 28543
rect 3985 28509 4019 28543
rect 4721 28509 4755 28543
rect 4997 28509 5031 28543
rect 5089 28509 5123 28543
rect 8953 28509 8987 28543
rect 13185 28509 13219 28543
rect 13277 28509 13311 28543
rect 13369 28509 13403 28543
rect 13553 28509 13587 28543
rect 14105 28509 14139 28543
rect 14198 28509 14232 28543
rect 14473 28509 14507 28543
rect 14570 28509 14604 28543
rect 17049 28509 17083 28543
rect 21281 28509 21315 28543
rect 21373 28509 21407 28543
rect 21649 28509 21683 28543
rect 29009 28509 29043 28543
rect 30757 28509 30791 28543
rect 31217 28509 31251 28543
rect 31401 28509 31435 28543
rect 31861 28509 31895 28543
rect 33793 28509 33827 28543
rect 34897 28509 34931 28543
rect 34989 28509 35023 28543
rect 35265 28509 35299 28543
rect 36093 28509 36127 28543
rect 36277 28509 36311 28543
rect 38402 28509 38436 28543
rect 38669 28509 38703 28543
rect 2973 28441 3007 28475
rect 4169 28441 4203 28475
rect 4905 28441 4939 28475
rect 7665 28441 7699 28475
rect 9198 28441 9232 28475
rect 14381 28441 14415 28475
rect 16322 28441 16356 28475
rect 21465 28441 21499 28475
rect 22661 28441 22695 28475
rect 25145 28441 25179 28475
rect 35081 28441 35115 28475
rect 5273 28373 5307 28407
rect 11989 28373 12023 28407
rect 12909 28373 12943 28407
rect 14749 28373 14783 28407
rect 17233 28373 17267 28407
rect 21097 28373 21131 28407
rect 22753 28373 22787 28407
rect 23765 28373 23799 28407
rect 31401 28373 31435 28407
rect 34713 28373 34747 28407
rect 37289 28373 37323 28407
rect 3985 28169 4019 28203
rect 9413 28169 9447 28203
rect 10057 28169 10091 28203
rect 13093 28169 13127 28203
rect 13921 28169 13955 28203
rect 16037 28169 16071 28203
rect 6745 28101 6779 28135
rect 12725 28101 12759 28135
rect 12817 28101 12851 28135
rect 13737 28101 13771 28135
rect 34253 28101 34287 28135
rect 2872 28033 2906 28067
rect 6377 28033 6411 28067
rect 6470 28033 6504 28067
rect 6653 28033 6687 28067
rect 6842 28033 6876 28067
rect 9321 28033 9355 28067
rect 9505 28033 9539 28067
rect 11713 28033 11747 28067
rect 11897 28033 11931 28067
rect 12541 28033 12575 28067
rect 12909 28033 12943 28067
rect 13553 28033 13587 28067
rect 15393 28033 15427 28067
rect 15577 28033 15611 28067
rect 15669 28033 15703 28067
rect 15761 28033 15795 28067
rect 17141 28033 17175 28067
rect 18061 28033 18095 28067
rect 19993 28033 20027 28067
rect 26433 28033 26467 28067
rect 27261 28033 27295 28067
rect 30021 28033 30055 28067
rect 31585 28033 31619 28067
rect 32137 28033 32171 28067
rect 34161 28033 34195 28067
rect 34345 28033 34379 28067
rect 34529 28033 34563 28067
rect 39701 28033 39735 28067
rect 2605 27965 2639 27999
rect 14933 27965 14967 27999
rect 17785 27965 17819 27999
rect 19717 27965 19751 27999
rect 30297 27965 30331 27999
rect 31309 27965 31343 27999
rect 39957 27965 39991 27999
rect 24685 27897 24719 27931
rect 58173 27897 58207 27931
rect 7021 27829 7055 27863
rect 8861 27829 8895 27863
rect 10609 27829 10643 27863
rect 11529 27829 11563 27863
rect 17233 27829 17267 27863
rect 19165 27829 19199 27863
rect 27077 27829 27111 27863
rect 29009 27829 29043 27863
rect 33977 27829 34011 27863
rect 38577 27829 38611 27863
rect 9045 27625 9079 27659
rect 13553 27625 13587 27659
rect 16957 27625 16991 27659
rect 29009 27557 29043 27591
rect 30481 27557 30515 27591
rect 9597 27489 9631 27523
rect 12173 27489 12207 27523
rect 31033 27489 31067 27523
rect 4905 27421 4939 27455
rect 4998 27421 5032 27455
rect 5273 27421 5307 27455
rect 5411 27421 5445 27455
rect 7297 27421 7331 27455
rect 8401 27421 8435 27455
rect 8953 27421 8987 27455
rect 9137 27421 9171 27455
rect 9873 27421 9907 27455
rect 10885 27421 10919 27455
rect 11161 27421 11195 27455
rect 12440 27421 12474 27455
rect 17785 27421 17819 27455
rect 18245 27421 18279 27455
rect 19257 27421 19291 27455
rect 22845 27421 22879 27455
rect 23397 27421 23431 27455
rect 26617 27421 26651 27455
rect 31309 27421 31343 27455
rect 32505 27421 32539 27455
rect 32597 27421 32631 27455
rect 32873 27421 32907 27455
rect 33471 27421 33505 27455
rect 33609 27421 33643 27455
rect 33885 27421 33919 27455
rect 34897 27421 34931 27455
rect 5181 27353 5215 27387
rect 7113 27353 7147 27387
rect 21097 27353 21131 27387
rect 25973 27353 26007 27387
rect 26157 27353 26191 27387
rect 26884 27353 26918 27387
rect 28825 27353 28859 27387
rect 32689 27353 32723 27387
rect 33701 27353 33735 27387
rect 34713 27353 34747 27387
rect 5549 27285 5583 27319
rect 7481 27285 7515 27319
rect 16313 27285 16347 27319
rect 18429 27285 18463 27319
rect 19441 27285 19475 27319
rect 24685 27285 24719 27319
rect 25789 27285 25823 27319
rect 27997 27285 28031 27319
rect 29561 27285 29595 27319
rect 32321 27285 32355 27319
rect 33333 27285 33367 27319
rect 35081 27285 35115 27319
rect 2697 27081 2731 27115
rect 6377 27081 6411 27115
rect 10149 27081 10183 27115
rect 11529 27081 11563 27115
rect 16037 27081 16071 27115
rect 17049 27081 17083 27115
rect 25697 27081 25731 27115
rect 3341 27013 3375 27047
rect 5089 27013 5123 27047
rect 5181 27013 5215 27047
rect 10977 27013 11011 27047
rect 15485 27013 15519 27047
rect 21189 27013 21223 27047
rect 24501 27013 24535 27047
rect 31493 27013 31527 27047
rect 3525 26945 3559 26979
rect 4813 26945 4847 26979
rect 4906 26945 4940 26979
rect 5319 26945 5353 26979
rect 7490 26945 7524 26979
rect 9321 26945 9355 26979
rect 9505 26945 9539 26979
rect 10793 26945 10827 26979
rect 12357 26945 12391 26979
rect 15945 26945 15979 26979
rect 16129 26945 16163 26979
rect 16865 26945 16899 26979
rect 17785 26945 17819 26979
rect 18429 26945 18463 26979
rect 20186 26945 20220 26979
rect 22468 26945 22502 26979
rect 25053 26945 25087 26979
rect 25216 26948 25250 26982
rect 25329 26945 25363 26979
rect 25467 26945 25501 26979
rect 29294 26945 29328 26979
rect 32413 26945 32447 26979
rect 32597 26945 32631 26979
rect 32689 26945 32723 26979
rect 32781 26945 32815 26979
rect 34253 26945 34287 26979
rect 34437 26945 34471 26979
rect 34529 26945 34563 26979
rect 34621 26945 34655 26979
rect 39701 26945 39735 26979
rect 7757 26877 7791 26911
rect 12081 26877 12115 26911
rect 16681 26877 16715 26911
rect 20453 26877 20487 26911
rect 22201 26877 22235 26911
rect 29561 26877 29595 26911
rect 39957 26877 39991 26911
rect 4077 26809 4111 26843
rect 9321 26809 9355 26843
rect 17969 26809 18003 26843
rect 33793 26809 33827 26843
rect 3157 26741 3191 26775
rect 5457 26741 5491 26775
rect 19073 26741 19107 26775
rect 23581 26741 23615 26775
rect 26157 26741 26191 26775
rect 28181 26741 28215 26775
rect 33057 26741 33091 26775
rect 34897 26741 34931 26775
rect 38577 26741 38611 26775
rect 58173 26741 58207 26775
rect 5089 26537 5123 26571
rect 7297 26537 7331 26571
rect 11713 26537 11747 26571
rect 19901 26537 19935 26571
rect 22201 26537 22235 26571
rect 28733 26537 28767 26571
rect 31493 26537 31527 26571
rect 34713 26537 34747 26571
rect 5641 26469 5675 26503
rect 12633 26469 12667 26503
rect 18061 26469 18095 26503
rect 27077 26469 27111 26503
rect 23029 26401 23063 26435
rect 32045 26401 32079 26435
rect 2881 26333 2915 26367
rect 2973 26333 3007 26367
rect 3065 26333 3099 26367
rect 3249 26333 3283 26367
rect 3985 26333 4019 26367
rect 6101 26333 6135 26367
rect 6285 26333 6319 26367
rect 6377 26333 6411 26367
rect 6469 26333 6503 26367
rect 7573 26333 7607 26367
rect 7665 26333 7699 26367
rect 7757 26333 7791 26367
rect 7941 26333 7975 26367
rect 9321 26333 9355 26367
rect 16681 26333 16715 26367
rect 19257 26333 19291 26367
rect 19441 26333 19475 26367
rect 19533 26333 19567 26367
rect 19625 26333 19659 26367
rect 20453 26333 20487 26367
rect 20637 26333 20671 26367
rect 20729 26333 20763 26367
rect 20821 26333 20855 26367
rect 21557 26333 21591 26367
rect 21741 26333 21775 26367
rect 21833 26333 21867 26367
rect 21925 26333 21959 26367
rect 22845 26333 22879 26367
rect 24593 26333 24627 26367
rect 24756 26327 24790 26361
rect 24869 26333 24903 26367
rect 25007 26333 25041 26367
rect 25697 26333 25731 26367
rect 33793 26333 33827 26367
rect 35826 26333 35860 26367
rect 36093 26333 36127 26367
rect 38945 26333 38979 26367
rect 39313 26333 39347 26367
rect 2605 26265 2639 26299
rect 4169 26265 4203 26299
rect 11805 26265 11839 26299
rect 12449 26265 12483 26299
rect 16948 26265 16982 26299
rect 21097 26265 21131 26299
rect 22661 26265 22695 26299
rect 25237 26265 25271 26299
rect 25942 26265 25976 26299
rect 27537 26265 27571 26299
rect 27721 26265 27755 26299
rect 39129 26265 39163 26299
rect 39865 26265 39899 26299
rect 40049 26265 40083 26299
rect 3801 26197 3835 26231
rect 6745 26197 6779 26231
rect 10609 26197 10643 26231
rect 13093 26197 13127 26231
rect 27905 26197 27939 26231
rect 40233 26197 40267 26231
rect 3985 25993 4019 26027
rect 5825 25993 5859 26027
rect 13553 25993 13587 26027
rect 17325 25993 17359 26027
rect 18889 25993 18923 26027
rect 20913 25993 20947 26027
rect 26249 25993 26283 26027
rect 32781 25993 32815 26027
rect 38209 25993 38243 26027
rect 2872 25925 2906 25959
rect 5457 25925 5491 25959
rect 5641 25925 5675 25959
rect 7297 25925 7331 25959
rect 9321 25925 9355 25959
rect 18521 25925 18555 25959
rect 19717 25925 19751 25959
rect 20453 25925 20487 25959
rect 21281 25925 21315 25959
rect 22078 25925 22112 25959
rect 26985 25925 27019 25959
rect 28641 25925 28675 25959
rect 29837 25925 29871 25959
rect 33894 25925 33928 25959
rect 38761 25925 38795 25959
rect 2605 25857 2639 25891
rect 6929 25857 6963 25891
rect 7022 25857 7056 25891
rect 7205 25857 7239 25891
rect 7435 25857 7469 25891
rect 9505 25857 9539 25891
rect 10333 25857 10367 25891
rect 11897 25857 11931 25891
rect 13645 25857 13679 25891
rect 15669 25857 15703 25891
rect 16865 25857 16899 25891
rect 17601 25857 17635 25891
rect 17693 25857 17727 25891
rect 17785 25857 17819 25891
rect 17969 25857 18003 25891
rect 18705 25857 18739 25891
rect 19533 25857 19567 25891
rect 21097 25857 21131 25891
rect 25605 25857 25639 25891
rect 25768 25857 25802 25891
rect 25881 25857 25915 25891
rect 26019 25857 26053 25891
rect 28825 25857 28859 25891
rect 30021 25857 30055 25891
rect 10057 25789 10091 25823
rect 12173 25789 12207 25823
rect 15393 25789 15427 25823
rect 19349 25789 19383 25823
rect 21833 25789 21867 25823
rect 34161 25789 34195 25823
rect 7573 25721 7607 25755
rect 40049 25721 40083 25755
rect 6377 25653 6411 25687
rect 8125 25653 8159 25687
rect 16681 25653 16715 25687
rect 23213 25653 23247 25687
rect 29009 25653 29043 25687
rect 30205 25653 30239 25687
rect 31125 25653 31159 25687
rect 37473 25653 37507 25687
rect 7757 25449 7791 25483
rect 25789 25449 25823 25483
rect 39221 25449 39255 25483
rect 39865 25449 39899 25483
rect 41613 25449 41647 25483
rect 10609 25381 10643 25415
rect 20085 25381 20119 25415
rect 31401 25381 31435 25415
rect 2145 25313 2179 25347
rect 15853 25313 15887 25347
rect 18061 25313 18095 25347
rect 18337 25313 18371 25347
rect 2881 25245 2915 25279
rect 2973 25245 3007 25279
rect 3065 25245 3099 25279
rect 3249 25245 3283 25279
rect 6377 25245 6411 25279
rect 10793 25245 10827 25279
rect 11529 25245 11563 25279
rect 15669 25245 15703 25279
rect 16313 25245 16347 25279
rect 21695 25245 21729 25279
rect 21833 25245 21867 25279
rect 22063 25245 22097 25279
rect 22201 25245 22235 25279
rect 26157 25245 26191 25279
rect 28549 25245 28583 25279
rect 30297 25245 30331 25279
rect 30481 25245 30515 25279
rect 30573 25245 30607 25279
rect 30711 25245 30745 25279
rect 32781 25245 32815 25279
rect 37105 25245 37139 25279
rect 37841 25245 37875 25279
rect 37933 25245 37967 25279
rect 38025 25245 38059 25279
rect 38209 25245 38243 25279
rect 40141 25245 40175 25279
rect 40233 25245 40267 25279
rect 40325 25245 40359 25279
rect 40509 25245 40543 25279
rect 40969 25245 41003 25279
rect 41153 25245 41187 25279
rect 41245 25242 41279 25276
rect 41383 25245 41417 25279
rect 58173 25245 58207 25279
rect 4169 25177 4203 25211
rect 5917 25177 5951 25211
rect 6644 25177 6678 25211
rect 14933 25177 14967 25211
rect 15117 25177 15151 25211
rect 21925 25177 21959 25211
rect 25973 25177 26007 25211
rect 26801 25177 26835 25211
rect 30941 25177 30975 25211
rect 32514 25177 32548 25211
rect 36860 25177 36894 25211
rect 37565 25177 37599 25211
rect 2605 25109 2639 25143
rect 11437 25109 11471 25143
rect 13277 25109 13311 25143
rect 14749 25109 14783 25143
rect 17049 25109 17083 25143
rect 19349 25109 19383 25143
rect 21557 25109 21591 25143
rect 29837 25109 29871 25143
rect 35725 25109 35759 25143
rect 6469 24905 6503 24939
rect 24409 24905 24443 24939
rect 37657 24905 37691 24939
rect 2872 24837 2906 24871
rect 32505 24837 32539 24871
rect 2605 24769 2639 24803
rect 9853 24769 9887 24803
rect 9962 24769 9996 24803
rect 10062 24769 10096 24803
rect 10241 24769 10275 24803
rect 14453 24769 14487 24803
rect 17969 24769 18003 24803
rect 18153 24769 18187 24803
rect 18245 24769 18279 24803
rect 18337 24769 18371 24803
rect 19073 24769 19107 24803
rect 19340 24769 19374 24803
rect 22433 24769 22467 24803
rect 22569 24769 22603 24803
rect 22661 24769 22695 24803
rect 22844 24769 22878 24803
rect 22937 24769 22971 24803
rect 24961 24769 24995 24803
rect 25145 24769 25179 24803
rect 25237 24769 25271 24803
rect 25329 24769 25363 24803
rect 28549 24769 28583 24803
rect 28816 24769 28850 24803
rect 30665 24769 30699 24803
rect 30754 24772 30788 24806
rect 30854 24769 30888 24803
rect 31033 24769 31067 24803
rect 32321 24769 32355 24803
rect 32689 24769 32723 24803
rect 37289 24769 37323 24803
rect 37473 24769 37507 24803
rect 39885 24769 39919 24803
rect 40141 24769 40175 24803
rect 14197 24701 14231 24735
rect 25605 24701 25639 24735
rect 3985 24633 4019 24667
rect 13645 24633 13679 24667
rect 9045 24565 9079 24599
rect 9597 24565 9631 24599
rect 11621 24565 11655 24599
rect 12633 24565 12667 24599
rect 13093 24565 13127 24599
rect 15577 24565 15611 24599
rect 18613 24565 18647 24599
rect 20453 24565 20487 24599
rect 22293 24565 22327 24599
rect 29929 24565 29963 24599
rect 30389 24565 30423 24599
rect 31493 24565 31527 24599
rect 38761 24565 38795 24599
rect 40877 24565 40911 24599
rect 3801 24361 3835 24395
rect 10793 24361 10827 24395
rect 14105 24361 14139 24395
rect 16129 24361 16163 24395
rect 19257 24361 19291 24395
rect 24685 24361 24719 24395
rect 29009 24361 29043 24395
rect 18705 24293 18739 24327
rect 29561 24293 29595 24327
rect 15209 24225 15243 24259
rect 30941 24225 30975 24259
rect 8953 24157 8987 24191
rect 12081 24157 12115 24191
rect 12173 24157 12207 24191
rect 12265 24157 12299 24191
rect 12449 24157 12483 24191
rect 12909 24157 12943 24191
rect 13093 24157 13127 24191
rect 13185 24157 13219 24191
rect 13323 24157 13357 24191
rect 14335 24157 14369 24191
rect 14470 24151 14504 24185
rect 14565 24154 14599 24188
rect 14749 24157 14783 24191
rect 15577 24157 15611 24191
rect 16313 24157 16347 24191
rect 17785 24157 17819 24191
rect 18061 24157 18095 24191
rect 18521 24157 18555 24191
rect 19441 24157 19475 24191
rect 21419 24157 21453 24191
rect 21777 24157 21811 24191
rect 21925 24157 21959 24191
rect 25513 24157 25547 24191
rect 28825 24157 28859 24191
rect 30674 24157 30708 24191
rect 41245 24157 41279 24191
rect 58173 24157 58207 24191
rect 9220 24089 9254 24123
rect 10977 24089 11011 24123
rect 11161 24089 11195 24123
rect 15393 24089 15427 24123
rect 19625 24089 19659 24123
rect 21557 24089 21591 24123
rect 21649 24089 21683 24123
rect 24869 24089 24903 24123
rect 25053 24089 25087 24123
rect 25758 24089 25792 24123
rect 28641 24089 28675 24123
rect 40233 24089 40267 24123
rect 40417 24089 40451 24123
rect 41061 24089 41095 24123
rect 10333 24021 10367 24055
rect 11805 24021 11839 24055
rect 13553 24021 13587 24055
rect 21281 24021 21315 24055
rect 26893 24021 26927 24055
rect 40601 24021 40635 24055
rect 41429 24021 41463 24055
rect 8953 23817 8987 23851
rect 12081 23817 12115 23851
rect 24409 23817 24443 23851
rect 24961 23817 24995 23851
rect 29101 23817 29135 23851
rect 41705 23817 41739 23851
rect 10977 23749 11011 23783
rect 11713 23749 11747 23783
rect 17049 23749 17083 23783
rect 17417 23749 17451 23783
rect 22661 23749 22695 23783
rect 22753 23749 22787 23783
rect 32965 23749 32999 23783
rect 33425 23749 33459 23783
rect 35909 23749 35943 23783
rect 39896 23749 39930 23783
rect 40601 23749 40635 23783
rect 2237 23681 2271 23715
rect 2421 23681 2455 23715
rect 9781 23681 9815 23715
rect 9873 23681 9907 23715
rect 9965 23681 9999 23715
rect 10149 23681 10183 23715
rect 10793 23681 10827 23715
rect 11897 23681 11931 23715
rect 13185 23681 13219 23715
rect 13452 23681 13486 23715
rect 17233 23681 17267 23715
rect 17877 23681 17911 23715
rect 18040 23681 18074 23715
rect 18140 23681 18174 23715
rect 18265 23681 18299 23715
rect 22385 23681 22419 23715
rect 22533 23681 22567 23715
rect 22850 23681 22884 23715
rect 25513 23681 25547 23715
rect 25697 23681 25731 23715
rect 25792 23681 25826 23715
rect 25901 23681 25935 23715
rect 29331 23681 29365 23715
rect 29469 23681 29503 23715
rect 29566 23681 29600 23715
rect 29745 23681 29779 23715
rect 32689 23681 32723 23715
rect 32781 23681 32815 23715
rect 33701 23681 33735 23715
rect 35817 23681 35851 23715
rect 36001 23681 36035 23715
rect 36185 23681 36219 23715
rect 40141 23681 40175 23715
rect 40857 23681 40891 23715
rect 40969 23681 41003 23715
rect 41066 23681 41100 23715
rect 41245 23681 41279 23715
rect 7389 23613 7423 23647
rect 7665 23613 7699 23647
rect 10609 23613 10643 23647
rect 30205 23613 30239 23647
rect 33609 23613 33643 23647
rect 37933 23613 37967 23647
rect 8217 23545 8251 23579
rect 14565 23545 14599 23579
rect 15117 23545 15151 23579
rect 35633 23545 35667 23579
rect 37473 23545 37507 23579
rect 2605 23477 2639 23511
rect 9505 23477 9539 23511
rect 12633 23477 12667 23511
rect 15853 23477 15887 23511
rect 18521 23477 18555 23511
rect 23029 23477 23063 23511
rect 26157 23477 26191 23511
rect 28641 23477 28675 23511
rect 32505 23477 32539 23511
rect 32689 23477 32723 23511
rect 33425 23477 33459 23511
rect 33885 23477 33919 23511
rect 38761 23477 38795 23511
rect 3801 23273 3835 23307
rect 18245 23273 18279 23307
rect 23213 23273 23247 23307
rect 40141 23273 40175 23307
rect 35909 23205 35943 23239
rect 25881 23137 25915 23171
rect 34161 23137 34195 23171
rect 2559 23069 2593 23103
rect 2697 23069 2731 23103
rect 2789 23069 2823 23103
rect 2973 23069 3007 23103
rect 7389 23069 7423 23103
rect 7665 23069 7699 23103
rect 8953 23069 8987 23103
rect 10977 23069 11011 23103
rect 11244 23069 11278 23103
rect 14841 23069 14875 23103
rect 15209 23069 15243 23103
rect 16037 23069 16071 23103
rect 23213 23069 23247 23103
rect 23305 23069 23339 23103
rect 24409 23069 24443 23103
rect 24685 23069 24719 23103
rect 26148 23069 26182 23103
rect 35081 23069 35115 23103
rect 35449 23069 35483 23103
rect 37289 23069 37323 23103
rect 38025 23069 38059 23103
rect 38117 23069 38151 23103
rect 38209 23069 38243 23103
rect 38393 23069 38427 23103
rect 40397 23069 40431 23103
rect 40509 23069 40543 23103
rect 40606 23069 40640 23103
rect 40785 23069 40819 23103
rect 9220 23001 9254 23035
rect 14381 23001 14415 23035
rect 15025 23001 15059 23035
rect 15117 23001 15151 23035
rect 20453 23001 20487 23035
rect 21005 23001 21039 23035
rect 33894 23001 33928 23035
rect 35173 23001 35207 23035
rect 35265 23001 35299 23035
rect 37044 23001 37078 23035
rect 37749 23001 37783 23035
rect 2329 22933 2363 22967
rect 8217 22933 8251 22967
rect 10333 22933 10367 22967
rect 12357 22933 12391 22967
rect 15393 22933 15427 22967
rect 17325 22933 17359 22967
rect 22293 22933 22327 22967
rect 23581 22933 23615 22967
rect 27261 22933 27295 22967
rect 28825 22933 28859 22967
rect 32781 22933 32815 22967
rect 34897 22933 34931 22967
rect 1593 22729 1627 22763
rect 3801 22729 3835 22763
rect 15945 22729 15979 22763
rect 19349 22729 19383 22763
rect 23765 22729 23799 22763
rect 25237 22729 25271 22763
rect 31585 22729 31619 22763
rect 33425 22729 33459 22763
rect 35633 22729 35667 22763
rect 37289 22729 37323 22763
rect 40049 22729 40083 22763
rect 1961 22661 1995 22695
rect 9505 22661 9539 22695
rect 10241 22661 10275 22695
rect 14473 22661 14507 22695
rect 15393 22661 15427 22695
rect 18236 22661 18270 22695
rect 24409 22661 24443 22695
rect 24593 22661 24627 22695
rect 27169 22661 27203 22695
rect 28457 22661 28491 22695
rect 31217 22661 31251 22695
rect 31309 22661 31343 22695
rect 33885 22661 33919 22695
rect 35909 22661 35943 22695
rect 37473 22661 37507 22695
rect 37657 22661 37691 22695
rect 1777 22593 1811 22627
rect 2421 22593 2455 22627
rect 2688 22593 2722 22627
rect 4445 22593 4479 22627
rect 4629 22593 4663 22627
rect 5457 22593 5491 22627
rect 5641 22593 5675 22627
rect 6561 22593 6595 22627
rect 6828 22593 6862 22627
rect 8585 22593 8619 22627
rect 9689 22593 9723 22627
rect 11805 22593 11839 22627
rect 11989 22593 12023 22627
rect 14381 22593 14415 22627
rect 14565 22593 14599 22627
rect 14749 22593 14783 22627
rect 17969 22593 18003 22627
rect 20177 22593 20211 22627
rect 21189 22593 21223 22627
rect 25053 22593 25087 22627
rect 27353 22593 27387 22627
rect 28641 22593 28675 22627
rect 31033 22593 31067 22627
rect 31401 22593 31435 22627
rect 32781 22593 32815 22627
rect 32944 22593 32978 22627
rect 33057 22593 33091 22627
rect 33149 22593 33183 22627
rect 34161 22593 34195 22627
rect 35817 22593 35851 22627
rect 36001 22593 36035 22627
rect 36185 22593 36219 22627
rect 38209 22593 38243 22627
rect 38393 22593 38427 22627
rect 12541 22525 12575 22559
rect 20085 22525 20119 22559
rect 21097 22525 21131 22559
rect 33977 22525 34011 22559
rect 7941 22457 7975 22491
rect 34345 22457 34379 22491
rect 58173 22457 58207 22491
rect 4261 22389 4295 22423
rect 5825 22389 5859 22423
rect 8401 22389 8435 22423
rect 11897 22389 11931 22423
rect 14197 22389 14231 22423
rect 16681 22389 16715 22423
rect 19809 22389 19843 22423
rect 19993 22389 20027 22423
rect 20821 22389 20855 22423
rect 21005 22389 21039 22423
rect 26985 22389 27019 22423
rect 28273 22389 28307 22423
rect 32229 22389 32263 22423
rect 33885 22389 33919 22423
rect 38577 22389 38611 22423
rect 3249 22185 3283 22219
rect 6837 22185 6871 22219
rect 8125 22185 8159 22219
rect 14933 22185 14967 22219
rect 21189 22185 21223 22219
rect 33333 22185 33367 22219
rect 37565 22185 37599 22219
rect 22017 22117 22051 22151
rect 15761 22049 15795 22083
rect 1869 21981 1903 22015
rect 3801 21981 3835 22015
rect 6193 21981 6227 22015
rect 6372 21981 6406 22015
rect 6469 21981 6503 22015
rect 6607 21981 6641 22015
rect 7665 21981 7699 22015
rect 9873 21981 9907 22015
rect 10241 21981 10275 22015
rect 11437 21981 11471 22015
rect 11713 21981 11747 22015
rect 11805 21981 11839 22015
rect 13553 21981 13587 22015
rect 14105 21981 14139 22015
rect 15577 21981 15611 22015
rect 16773 21981 16807 22015
rect 17049 21981 17083 22015
rect 21097 21981 21131 22015
rect 21189 21981 21223 22015
rect 22569 21981 22603 22015
rect 22753 21981 22787 22015
rect 22845 21981 22879 22015
rect 22937 21981 22971 22015
rect 27629 21981 27663 22015
rect 31769 21981 31803 22015
rect 32037 21981 32071 22015
rect 32183 21981 32217 22015
rect 32781 21981 32815 22015
rect 33057 21981 33091 22015
rect 33149 21981 33183 22015
rect 38945 21981 38979 22015
rect 2136 21913 2170 21947
rect 4046 21913 4080 21947
rect 7481 21913 7515 21947
rect 10057 21913 10091 21947
rect 10149 21913 10183 21947
rect 11621 21913 11655 21947
rect 27896 21913 27930 21947
rect 31953 21913 31987 21947
rect 32965 21913 32999 21947
rect 38678 21913 38712 21947
rect 5181 21845 5215 21879
rect 7297 21845 7331 21879
rect 9045 21845 9079 21879
rect 10425 21845 10459 21879
rect 11989 21845 12023 21879
rect 14289 21845 14323 21879
rect 15393 21845 15427 21879
rect 20821 21845 20855 21879
rect 23213 21845 23247 21879
rect 29009 21845 29043 21879
rect 32321 21845 32355 21879
rect 2145 21641 2179 21675
rect 3617 21641 3651 21675
rect 14841 21641 14875 21675
rect 15669 21641 15703 21675
rect 38485 21641 38519 21675
rect 5825 21573 5859 21607
rect 6622 21573 6656 21607
rect 10149 21573 10183 21607
rect 14289 21573 14323 21607
rect 20085 21573 20119 21607
rect 20729 21573 20763 21607
rect 23020 21573 23054 21607
rect 24961 21573 24995 21607
rect 27905 21573 27939 21607
rect 32965 21573 32999 21607
rect 2421 21505 2455 21539
rect 2513 21505 2547 21539
rect 2605 21505 2639 21539
rect 2789 21505 2823 21539
rect 3893 21505 3927 21539
rect 3985 21505 4019 21539
rect 4077 21505 4111 21539
rect 4261 21505 4295 21539
rect 5181 21505 5215 21539
rect 5344 21511 5378 21545
rect 5457 21505 5491 21539
rect 5549 21505 5583 21539
rect 9873 21505 9907 21539
rect 10057 21505 10091 21539
rect 10241 21505 10275 21539
rect 15761 21505 15795 21539
rect 17049 21505 17083 21539
rect 17141 21505 17175 21539
rect 17233 21505 17267 21539
rect 17417 21505 17451 21539
rect 20545 21505 20579 21539
rect 24593 21505 24627 21539
rect 24777 21505 24811 21539
rect 27445 21505 27479 21539
rect 28135 21505 28169 21539
rect 28273 21505 28307 21539
rect 28370 21511 28404 21545
rect 28549 21505 28583 21539
rect 29009 21505 29043 21539
rect 29745 21505 29779 21539
rect 30021 21505 30055 21539
rect 33149 21505 33183 21539
rect 38761 21505 38795 21539
rect 38853 21505 38887 21539
rect 38945 21505 38979 21539
rect 39129 21505 39163 21539
rect 6377 21437 6411 21471
rect 22753 21437 22787 21471
rect 29929 21437 29963 21471
rect 32781 21437 32815 21471
rect 7757 21369 7791 21403
rect 17877 21369 17911 21403
rect 29561 21369 29595 21403
rect 10425 21301 10459 21335
rect 16773 21301 16807 21335
rect 22201 21301 22235 21335
rect 24133 21301 24167 21335
rect 29837 21301 29871 21335
rect 37933 21301 37967 21335
rect 58173 21301 58207 21335
rect 5917 21097 5951 21131
rect 10149 21097 10183 21131
rect 14657 21097 14691 21131
rect 21189 21097 21223 21131
rect 21833 21097 21867 21131
rect 23029 21097 23063 21131
rect 10977 21029 11011 21063
rect 15945 21029 15979 21063
rect 19901 21029 19935 21063
rect 23489 21029 23523 21063
rect 12909 20893 12943 20927
rect 14565 20893 14599 20927
rect 15301 20893 15335 20927
rect 15394 20893 15428 20927
rect 15577 20893 15611 20927
rect 15807 20893 15841 20927
rect 16405 20893 16439 20927
rect 20080 20893 20114 20927
rect 20269 20893 20303 20927
rect 20452 20893 20486 20927
rect 20545 20893 20579 20927
rect 22385 20893 22419 20927
rect 22569 20893 22603 20927
rect 22661 20893 22695 20927
rect 22753 20893 22787 20927
rect 29009 20893 29043 20927
rect 30021 20893 30055 20927
rect 40601 20893 40635 20927
rect 2973 20825 3007 20859
rect 10425 20825 10459 20859
rect 11161 20825 11195 20859
rect 12725 20825 12759 20859
rect 15669 20825 15703 20859
rect 16672 20825 16706 20859
rect 20177 20825 20211 20859
rect 21097 20825 21131 20859
rect 23673 20825 23707 20859
rect 23857 20825 23891 20859
rect 25697 20825 25731 20859
rect 27445 20825 27479 20859
rect 30205 20825 30239 20859
rect 40417 20825 40451 20859
rect 41245 20825 41279 20859
rect 4445 20757 4479 20791
rect 6653 20757 6687 20791
rect 9505 20757 9539 20791
rect 11713 20757 11747 20791
rect 13093 20757 13127 20791
rect 17785 20757 17819 20791
rect 28457 20757 28491 20791
rect 37473 20757 37507 20791
rect 40785 20757 40819 20791
rect 7113 20553 7147 20587
rect 8033 20553 8067 20587
rect 13645 20553 13679 20587
rect 17141 20553 17175 20587
rect 27537 20553 27571 20587
rect 28733 20553 28767 20587
rect 29837 20553 29871 20587
rect 30297 20553 30331 20587
rect 37289 20553 37323 20587
rect 17325 20485 17359 20519
rect 19625 20485 19659 20519
rect 20729 20485 20763 20519
rect 22109 20485 22143 20519
rect 30757 20485 30791 20519
rect 33241 20485 33275 20519
rect 34814 20485 34848 20519
rect 37657 20485 37691 20519
rect 39120 20485 39154 20519
rect 40693 20485 40727 20519
rect 7205 20417 7239 20451
rect 8125 20417 8159 20451
rect 12532 20417 12566 20451
rect 14381 20417 14415 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 17509 20417 17543 20451
rect 18337 20417 18371 20451
rect 19436 20417 19470 20451
rect 19533 20417 19567 20451
rect 19808 20417 19842 20451
rect 19901 20417 19935 20451
rect 20361 20417 20395 20451
rect 20454 20417 20488 20451
rect 20637 20417 20671 20451
rect 20826 20417 20860 20451
rect 23029 20417 23063 20451
rect 23296 20417 23330 20451
rect 26166 20417 26200 20451
rect 27445 20417 27479 20451
rect 28641 20417 28675 20451
rect 29285 20417 29319 20451
rect 29469 20417 29503 20451
rect 29561 20417 29595 20451
rect 29653 20417 29687 20451
rect 30481 20417 30515 20451
rect 32597 20417 32631 20451
rect 32781 20417 32815 20451
rect 32876 20417 32910 20451
rect 32965 20417 32999 20451
rect 37473 20417 37507 20451
rect 37565 20417 37599 20451
rect 37841 20417 37875 20451
rect 40923 20417 40957 20451
rect 41058 20417 41092 20451
rect 41158 20417 41192 20451
rect 41337 20417 41371 20451
rect 4997 20349 5031 20383
rect 12265 20349 12299 20383
rect 14105 20349 14139 20383
rect 15485 20349 15519 20383
rect 18245 20349 18279 20383
rect 26433 20349 26467 20383
rect 30573 20349 30607 20383
rect 35081 20349 35115 20383
rect 38853 20349 38887 20383
rect 19257 20281 19291 20315
rect 25053 20281 25087 20315
rect 17969 20213 18003 20247
rect 18153 20213 18187 20247
rect 21005 20213 21039 20247
rect 24409 20213 24443 20247
rect 30481 20213 30515 20247
rect 33701 20213 33735 20247
rect 40233 20213 40267 20247
rect 6377 20009 6411 20043
rect 9137 20009 9171 20043
rect 11345 20009 11379 20043
rect 12449 20009 12483 20043
rect 15209 20009 15243 20043
rect 21833 20009 21867 20043
rect 25789 20009 25823 20043
rect 27721 20009 27755 20043
rect 29009 20009 29043 20043
rect 32965 20009 32999 20043
rect 41429 20009 41463 20043
rect 4629 19873 4663 19907
rect 15209 19873 15243 19907
rect 22385 19873 22419 19907
rect 26893 19873 26927 19907
rect 36277 19873 36311 19907
rect 2513 19805 2547 19839
rect 9229 19805 9263 19839
rect 9321 19805 9355 19839
rect 12679 19805 12713 19839
rect 12814 19805 12848 19839
rect 12909 19805 12943 19839
rect 13093 19805 13127 19839
rect 14473 19805 14507 19839
rect 15301 19805 15335 19839
rect 21741 19805 21775 19839
rect 21925 19805 21959 19839
rect 26065 19805 26099 19839
rect 26154 19805 26188 19839
rect 26249 19805 26283 19839
rect 26433 19805 26467 19839
rect 27077 19805 27111 19839
rect 28457 19805 28491 19839
rect 28825 19805 28859 19839
rect 29837 19805 29871 19839
rect 30113 19805 30147 19839
rect 33149 19805 33183 19839
rect 33333 19805 33367 19839
rect 36001 19805 36035 19839
rect 37565 19805 37599 19839
rect 40601 19805 40635 19839
rect 40693 19805 40727 19839
rect 40785 19805 40819 19839
rect 40969 19805 41003 19839
rect 58173 19805 58207 19839
rect 3893 19737 3927 19771
rect 4445 19737 4479 19771
rect 5825 19737 5859 19771
rect 6653 19737 6687 19771
rect 9873 19737 9907 19771
rect 27261 19737 27295 19771
rect 28641 19737 28675 19771
rect 28733 19737 28767 19771
rect 2329 19669 2363 19703
rect 5181 19669 5215 19703
rect 7573 19669 7607 19703
rect 8953 19669 8987 19703
rect 11989 19669 12023 19703
rect 14289 19669 14323 19703
rect 14933 19669 14967 19703
rect 15853 19669 15887 19703
rect 32505 19669 32539 19703
rect 38853 19669 38887 19703
rect 40325 19669 40359 19703
rect 3341 19465 3375 19499
rect 10609 19465 10643 19499
rect 14197 19465 14231 19499
rect 15301 19465 15335 19499
rect 18797 19465 18831 19499
rect 22385 19465 22419 19499
rect 26433 19465 26467 19499
rect 26985 19465 27019 19499
rect 29193 19465 29227 19499
rect 30941 19465 30975 19499
rect 35817 19465 35851 19499
rect 40141 19465 40175 19499
rect 40969 19465 41003 19499
rect 3801 19397 3835 19431
rect 25421 19397 25455 19431
rect 25513 19397 25547 19431
rect 27445 19397 27479 19431
rect 28917 19397 28951 19431
rect 31401 19397 31435 19431
rect 36093 19397 36127 19431
rect 36185 19397 36219 19431
rect 39028 19397 39062 19431
rect 1961 19329 1995 19363
rect 2228 19329 2262 19363
rect 6653 19329 6687 19363
rect 6920 19329 6954 19363
rect 9229 19329 9263 19363
rect 9496 19329 9530 19363
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 14197 19329 14231 19363
rect 14381 19329 14415 19363
rect 15669 19329 15703 19363
rect 17417 19329 17451 19363
rect 17673 19329 17707 19363
rect 21281 19329 21315 19363
rect 22201 19329 22235 19363
rect 25237 19329 25271 19363
rect 25605 19329 25639 19363
rect 27169 19329 27203 19363
rect 28641 19329 28675 19363
rect 28825 19329 28859 19363
rect 29009 19329 29043 19363
rect 31125 19329 31159 19363
rect 31217 19329 31251 19363
rect 33802 19329 33836 19363
rect 34069 19329 34103 19363
rect 36001 19329 36035 19363
rect 36369 19329 36403 19363
rect 37565 19329 37599 19363
rect 40601 19329 40635 19363
rect 40785 19329 40819 19363
rect 15577 19261 15611 19295
rect 21005 19261 21039 19295
rect 22017 19261 22051 19295
rect 22845 19261 22879 19295
rect 27261 19261 27295 19295
rect 29653 19261 29687 19295
rect 29929 19261 29963 19295
rect 37289 19261 37323 19295
rect 38761 19261 38795 19295
rect 5089 19193 5123 19227
rect 12357 19193 12391 19227
rect 25789 19193 25823 19227
rect 32689 19193 32723 19227
rect 8033 19125 8067 19159
rect 8493 19125 8527 19159
rect 11529 19125 11563 19159
rect 15485 19125 15519 19159
rect 27169 19125 27203 19159
rect 27905 19125 27939 19159
rect 31125 19125 31159 19159
rect 2513 18921 2547 18955
rect 5457 18921 5491 18955
rect 7205 18921 7239 18955
rect 8309 18921 8343 18955
rect 10425 18921 10459 18955
rect 14473 18921 14507 18955
rect 17509 18921 17543 18955
rect 22201 18921 22235 18955
rect 30205 18921 30239 18955
rect 30849 18921 30883 18955
rect 35909 18921 35943 18955
rect 37289 18921 37323 18955
rect 4077 18853 4111 18887
rect 23213 18853 23247 18887
rect 30665 18853 30699 18887
rect 32781 18853 32815 18887
rect 4721 18785 4755 18819
rect 8309 18785 8343 18819
rect 24409 18785 24443 18819
rect 24685 18785 24719 18819
rect 34161 18785 34195 18819
rect 2697 18717 2731 18751
rect 2789 18717 2823 18751
rect 4445 18717 4479 18751
rect 7021 18717 7055 18751
rect 8401 18717 8435 18751
rect 10701 18717 10735 18751
rect 10793 18717 10827 18751
rect 10885 18717 10919 18751
rect 11069 18717 11103 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 11989 18717 12023 18751
rect 12173 18717 12207 18751
rect 12817 18717 12851 18751
rect 17049 18717 17083 18751
rect 17785 18717 17819 18751
rect 17877 18717 17911 18751
rect 17969 18717 18003 18751
rect 18153 18717 18187 18751
rect 20821 18717 20855 18751
rect 25973 18717 26007 18751
rect 29653 18717 29687 18751
rect 29837 18717 29871 18751
rect 30021 18717 30055 18751
rect 30849 18717 30883 18751
rect 30941 18717 30975 18751
rect 31125 18717 31159 18751
rect 32137 18717 32171 18751
rect 36093 18717 36127 18751
rect 36277 18717 36311 18751
rect 36461 18717 36495 18751
rect 37473 18717 37507 18751
rect 37565 18717 37599 18751
rect 37841 18717 37875 18751
rect 40141 18717 40175 18751
rect 58173 18717 58207 18751
rect 4537 18649 4571 18683
rect 5365 18649 5399 18683
rect 6469 18649 6503 18683
rect 9873 18649 9907 18683
rect 12633 18649 12667 18683
rect 13001 18649 13035 18683
rect 21066 18649 21100 18683
rect 23029 18649 23063 18683
rect 26157 18649 26191 18683
rect 27445 18649 27479 18683
rect 29929 18649 29963 18683
rect 31953 18649 31987 18683
rect 33894 18649 33928 18683
rect 36185 18649 36219 18683
rect 37657 18649 37691 18683
rect 39957 18649 39991 18683
rect 6377 18581 6411 18615
rect 8033 18581 8067 18615
rect 9321 18581 9355 18615
rect 11529 18581 11563 18615
rect 25789 18581 25823 18615
rect 26617 18581 26651 18615
rect 27537 18581 27571 18615
rect 32321 18581 32355 18615
rect 40325 18581 40359 18615
rect 6837 18377 6871 18411
rect 8493 18377 8527 18411
rect 18061 18377 18095 18411
rect 20913 18377 20947 18411
rect 22661 18377 22695 18411
rect 31493 18377 31527 18411
rect 33057 18377 33091 18411
rect 33517 18377 33551 18411
rect 34713 18377 34747 18411
rect 40141 18377 40175 18411
rect 9864 18309 9898 18343
rect 18245 18309 18279 18343
rect 19809 18309 19843 18343
rect 21833 18309 21867 18343
rect 22017 18309 22051 18343
rect 22201 18309 22235 18343
rect 24777 18309 24811 18343
rect 24869 18309 24903 18343
rect 39028 18309 39062 18343
rect 41245 18309 41279 18343
rect 2237 18241 2271 18275
rect 2329 18241 2363 18275
rect 2513 18241 2547 18275
rect 3157 18241 3191 18275
rect 4169 18241 4203 18275
rect 4261 18241 4295 18275
rect 5457 18241 5491 18275
rect 7021 18241 7055 18275
rect 7389 18241 7423 18275
rect 7573 18241 7607 18275
rect 9597 18241 9631 18275
rect 11897 18241 11931 18275
rect 14289 18241 14323 18275
rect 14473 18241 14507 18275
rect 18429 18241 18463 18275
rect 20269 18241 20303 18275
rect 20453 18241 20487 18275
rect 20545 18241 20579 18275
rect 20683 18241 20717 18275
rect 22845 18241 22879 18275
rect 24593 18241 24627 18275
rect 24961 18241 24995 18275
rect 25789 18241 25823 18275
rect 26065 18241 26099 18275
rect 32413 18241 32447 18275
rect 32597 18241 32631 18275
rect 32692 18241 32726 18275
rect 32781 18241 32815 18275
rect 33793 18241 33827 18275
rect 33882 18241 33916 18275
rect 33982 18241 34016 18275
rect 34161 18241 34195 18275
rect 37565 18241 37599 18275
rect 40601 18241 40635 18275
rect 40785 18241 40819 18275
rect 40877 18241 40911 18275
rect 40969 18241 41003 18275
rect 4445 18173 4479 18207
rect 7205 18173 7239 18207
rect 7297 18173 7331 18207
rect 25881 18173 25915 18207
rect 37289 18173 37323 18207
rect 38761 18173 38795 18207
rect 3801 18105 3835 18139
rect 25145 18105 25179 18139
rect 2973 18037 3007 18071
rect 5641 18037 5675 18071
rect 10977 18037 11011 18071
rect 13185 18037 13219 18071
rect 14105 18037 14139 18071
rect 25605 18037 25639 18071
rect 25789 18037 25823 18071
rect 27169 18037 27203 18071
rect 5365 17833 5399 17867
rect 7113 17833 7147 17867
rect 15485 17833 15519 17867
rect 25881 17833 25915 17867
rect 26617 17833 26651 17867
rect 33057 17833 33091 17867
rect 39129 17833 39163 17867
rect 18337 17765 18371 17799
rect 37933 17765 37967 17799
rect 5089 17697 5123 17731
rect 14105 17697 14139 17731
rect 21373 17697 21407 17731
rect 40417 17697 40451 17731
rect 5181 17629 5215 17663
rect 12081 17629 12115 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 12449 17629 12483 17663
rect 12909 17629 12943 17663
rect 13093 17629 13127 17663
rect 13185 17629 13219 17663
rect 13277 17629 13311 17663
rect 17141 17629 17175 17663
rect 17233 17629 17267 17663
rect 17325 17629 17359 17663
rect 17509 17629 17543 17663
rect 24501 17629 24535 17663
rect 27997 17629 28031 17663
rect 31033 17629 31067 17663
rect 32873 17629 32907 17663
rect 33701 17629 33735 17663
rect 38945 17629 38979 17663
rect 7021 17561 7055 17595
rect 13553 17561 13587 17595
rect 14350 17561 14384 17595
rect 21618 17561 21652 17595
rect 24768 17561 24802 17595
rect 27730 17561 27764 17595
rect 32689 17561 32723 17595
rect 33517 17561 33551 17595
rect 36277 17561 36311 17595
rect 36461 17561 36495 17595
rect 37749 17561 37783 17595
rect 3893 17493 3927 17527
rect 4721 17493 4755 17527
rect 5917 17493 5951 17527
rect 6377 17493 6411 17527
rect 7665 17493 7699 17527
rect 11253 17493 11287 17527
rect 11805 17493 11839 17527
rect 16313 17493 16347 17527
rect 16865 17493 16899 17527
rect 22753 17493 22787 17527
rect 31217 17493 31251 17527
rect 33885 17493 33919 17527
rect 36093 17493 36127 17527
rect 11713 17289 11747 17323
rect 12357 17289 12391 17323
rect 13277 17289 13311 17323
rect 13921 17289 13955 17323
rect 25697 17289 25731 17323
rect 26985 17289 27019 17323
rect 36737 17289 36771 17323
rect 39957 17289 39991 17323
rect 2872 17221 2906 17255
rect 12541 17221 12575 17255
rect 14197 17221 14231 17255
rect 22017 17221 22051 17255
rect 22201 17221 22235 17255
rect 30205 17221 30239 17255
rect 7573 17153 7607 17187
rect 7941 17153 7975 17187
rect 8125 17153 8159 17187
rect 12725 17153 12759 17187
rect 14059 17153 14093 17187
rect 14289 17153 14323 17187
rect 14417 17153 14451 17187
rect 14565 17153 14599 17187
rect 15301 17153 15335 17187
rect 16681 17153 16715 17187
rect 16948 17153 16982 17187
rect 18797 17153 18831 17187
rect 18889 17153 18923 17187
rect 18981 17153 19015 17187
rect 19165 17153 19199 17187
rect 23029 17153 23063 17187
rect 24317 17153 24351 17187
rect 25927 17153 25961 17187
rect 26065 17153 26099 17187
rect 26157 17153 26191 17187
rect 26341 17153 26375 17187
rect 27261 17153 27295 17187
rect 27353 17156 27387 17190
rect 27445 17153 27479 17187
rect 27629 17153 27663 17187
rect 30021 17153 30055 17187
rect 32413 17153 32447 17187
rect 33425 17153 33459 17187
rect 33609 17153 33643 17187
rect 33701 17153 33735 17187
rect 33793 17153 33827 17187
rect 35624 17153 35658 17187
rect 40049 17153 40083 17187
rect 2605 17085 2639 17119
rect 7757 17085 7791 17119
rect 7849 17085 7883 17119
rect 15025 17085 15059 17119
rect 20269 17085 20303 17119
rect 22753 17085 22787 17119
rect 24041 17085 24075 17119
rect 32137 17085 32171 17119
rect 35357 17085 35391 17119
rect 58173 17017 58207 17051
rect 3985 16949 4019 16983
rect 5089 16949 5123 16983
rect 5733 16949 5767 16983
rect 7389 16949 7423 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 21833 16949 21867 16983
rect 30389 16949 30423 16983
rect 34069 16949 34103 16983
rect 10057 16745 10091 16779
rect 16313 16745 16347 16779
rect 17969 16745 18003 16779
rect 19257 16745 19291 16779
rect 21189 16745 21223 16779
rect 26709 16745 26743 16779
rect 33333 16745 33367 16779
rect 35725 16745 35759 16779
rect 20637 16677 20671 16711
rect 25605 16677 25639 16711
rect 35173 16677 35207 16711
rect 5181 16609 5215 16643
rect 5457 16609 5491 16643
rect 8401 16609 8435 16643
rect 29929 16609 29963 16643
rect 2421 16541 2455 16575
rect 5273 16541 5307 16575
rect 8134 16541 8168 16575
rect 10057 16541 10091 16575
rect 10241 16541 10275 16575
rect 17141 16541 17175 16575
rect 17233 16541 17267 16575
rect 17325 16541 17359 16575
rect 17509 16541 17543 16575
rect 18337 16541 18371 16575
rect 19625 16541 19659 16575
rect 21465 16541 21499 16575
rect 21557 16541 21591 16575
rect 21649 16541 21683 16575
rect 21833 16541 21867 16575
rect 26525 16541 26559 16575
rect 30205 16541 30239 16575
rect 36001 16541 36035 16575
rect 36093 16541 36127 16575
rect 36185 16541 36219 16575
rect 36369 16541 36403 16575
rect 37013 16541 37047 16575
rect 37381 16541 37415 16575
rect 39865 16541 39899 16575
rect 18153 16473 18187 16507
rect 19441 16473 19475 16507
rect 26341 16473 26375 16507
rect 27261 16473 27295 16507
rect 37105 16473 37139 16507
rect 37197 16473 37231 16507
rect 40049 16473 40083 16507
rect 2237 16405 2271 16439
rect 4813 16405 4847 16439
rect 7021 16405 7055 16439
rect 9505 16405 9539 16439
rect 10793 16405 10827 16439
rect 11529 16405 11563 16439
rect 16865 16405 16899 16439
rect 20085 16405 20119 16439
rect 22385 16405 22419 16439
rect 22845 16405 22879 16439
rect 28825 16405 28859 16439
rect 36829 16405 36863 16439
rect 40233 16405 40267 16439
rect 3341 16201 3375 16235
rect 4261 16201 4295 16235
rect 5641 16201 5675 16235
rect 9781 16201 9815 16235
rect 11897 16201 11931 16235
rect 17417 16201 17451 16235
rect 30021 16201 30055 16235
rect 32965 16201 32999 16235
rect 38301 16201 38335 16235
rect 40233 16201 40267 16235
rect 2228 16133 2262 16167
rect 4997 16133 5031 16167
rect 10609 16133 10643 16167
rect 12541 16133 12575 16167
rect 19993 16133 20027 16167
rect 20729 16133 20763 16167
rect 28273 16133 28307 16167
rect 28457 16133 28491 16167
rect 34078 16133 34112 16167
rect 37565 16133 37599 16167
rect 4169 16065 4203 16099
rect 5365 16065 5399 16099
rect 7113 16065 7147 16099
rect 7297 16065 7331 16099
rect 9137 16065 9171 16099
rect 9689 16065 9723 16099
rect 9873 16065 9907 16099
rect 10512 16065 10546 16099
rect 10701 16065 10735 16099
rect 10829 16065 10863 16099
rect 10977 16065 11011 16099
rect 11805 16065 11839 16099
rect 11989 16065 12023 16099
rect 14473 16065 14507 16099
rect 17601 16065 17635 16099
rect 17785 16065 17819 16099
rect 18245 16065 18279 16099
rect 20637 16065 20671 16099
rect 20821 16065 20855 16099
rect 22753 16065 22787 16099
rect 23029 16065 23063 16099
rect 23489 16065 23523 16099
rect 27169 16065 27203 16099
rect 28089 16065 28123 16099
rect 28917 16065 28951 16099
rect 29101 16065 29135 16099
rect 29193 16065 29227 16099
rect 29285 16065 29319 16099
rect 31134 16065 31168 16099
rect 35817 16065 35851 16099
rect 37473 16065 37507 16099
rect 37657 16065 37691 16099
rect 37841 16065 37875 16099
rect 38853 16065 38887 16099
rect 39120 16065 39154 16099
rect 1961 15997 1995 16031
rect 4445 15997 4479 16031
rect 5457 15997 5491 16031
rect 14749 15997 14783 16031
rect 23765 15997 23799 16031
rect 27353 15997 27387 16031
rect 31401 15997 31435 16031
rect 34345 15997 34379 16031
rect 35541 15997 35575 16031
rect 40693 15997 40727 16031
rect 40969 15997 41003 16031
rect 10333 15929 10367 15963
rect 26985 15929 27019 15963
rect 37289 15929 37323 15963
rect 3801 15861 3835 15895
rect 7113 15861 7147 15895
rect 7481 15861 7515 15895
rect 8033 15861 8067 15895
rect 8677 15861 8711 15895
rect 16957 15861 16991 15895
rect 26341 15861 26375 15895
rect 29561 15861 29595 15895
rect 58173 15861 58207 15895
rect 2513 15657 2547 15691
rect 9965 15657 9999 15691
rect 14473 15657 14507 15691
rect 18521 15657 18555 15691
rect 19349 15657 19383 15691
rect 19901 15657 19935 15691
rect 20361 15657 20395 15691
rect 22753 15657 22787 15691
rect 23397 15657 23431 15691
rect 26341 15657 26375 15691
rect 29561 15657 29595 15691
rect 36737 15657 36771 15691
rect 39865 15657 39899 15691
rect 13093 15589 13127 15623
rect 17233 15589 17267 15623
rect 22109 15589 22143 15623
rect 29009 15589 29043 15623
rect 2145 15521 2179 15555
rect 10057 15521 10091 15555
rect 11713 15521 11747 15555
rect 35633 15521 35667 15555
rect 37749 15521 37783 15555
rect 41061 15521 41095 15555
rect 2329 15453 2363 15487
rect 8309 15453 8343 15487
rect 10149 15453 10183 15487
rect 10788 15453 10822 15487
rect 11160 15453 11194 15487
rect 11253 15453 11287 15487
rect 11969 15453 12003 15487
rect 14289 15453 14323 15487
rect 14473 15453 14507 15487
rect 18337 15453 18371 15487
rect 18521 15453 18555 15487
rect 20361 15453 20395 15487
rect 20545 15453 20579 15487
rect 21925 15453 21959 15487
rect 22109 15453 22143 15487
rect 22569 15453 22603 15487
rect 22753 15453 22787 15487
rect 23213 15453 23247 15487
rect 23397 15453 23431 15487
rect 25789 15453 25823 15487
rect 26249 15453 26283 15487
rect 26433 15453 26467 15487
rect 28825 15453 28859 15487
rect 30674 15453 30708 15487
rect 30941 15453 30975 15487
rect 33333 15453 33367 15487
rect 33609 15453 33643 15487
rect 35357 15453 35391 15487
rect 38209 15453 38243 15487
rect 38393 15453 38427 15487
rect 38485 15453 38519 15487
rect 38577 15453 38611 15487
rect 40141 15453 40175 15487
rect 40230 15450 40264 15484
rect 40325 15447 40359 15481
rect 40509 15453 40543 15487
rect 8042 15385 8076 15419
rect 10885 15385 10919 15419
rect 10977 15385 11011 15419
rect 14933 15385 14967 15419
rect 24409 15385 24443 15419
rect 27077 15385 27111 15419
rect 27261 15385 27295 15419
rect 37381 15385 37415 15419
rect 37565 15385 37599 15419
rect 4721 15317 4755 15351
rect 6929 15317 6963 15351
rect 9781 15317 9815 15351
rect 10609 15317 10643 15351
rect 16313 15317 16347 15351
rect 17785 15317 17819 15351
rect 21373 15317 21407 15351
rect 26893 15317 26927 15351
rect 32873 15317 32907 15351
rect 38853 15317 38887 15351
rect 7297 15113 7331 15147
rect 14013 15113 14047 15147
rect 21097 15113 21131 15147
rect 30021 15113 30055 15147
rect 36093 15113 36127 15147
rect 40233 15113 40267 15147
rect 16037 15045 16071 15079
rect 23121 15045 23155 15079
rect 23213 15045 23247 15079
rect 27353 15045 27387 15079
rect 37841 15045 37875 15079
rect 39098 15045 39132 15079
rect 3433 14977 3467 15011
rect 3700 14977 3734 15011
rect 6561 14977 6595 15011
rect 6745 14977 6779 15011
rect 6837 14977 6871 15011
rect 7113 14977 7147 15011
rect 8125 14977 8159 15011
rect 10241 14977 10275 15011
rect 10425 14977 10459 15011
rect 12449 14977 12483 15011
rect 12597 14977 12631 15011
rect 12725 14977 12759 15011
rect 12817 14977 12851 15011
rect 12955 14977 12989 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 18061 14977 18095 15011
rect 18328 14977 18362 15011
rect 20269 14977 20303 15011
rect 20453 14977 20487 15011
rect 20913 14977 20947 15011
rect 21097 14977 21131 15011
rect 22293 14977 22327 15011
rect 22477 14977 22511 15011
rect 22937 14977 22971 15011
rect 23305 14977 23339 15011
rect 24225 14977 24259 15011
rect 24501 14977 24535 15011
rect 27537 14977 27571 15011
rect 30297 14977 30331 15011
rect 30389 14977 30423 15011
rect 30481 14977 30515 15011
rect 30665 14977 30699 15011
rect 33333 14977 33367 15011
rect 35449 14977 35483 15011
rect 35909 14977 35943 15011
rect 36093 14977 36127 15011
rect 36553 14977 36587 15011
rect 6929 14909 6963 14943
rect 8033 14909 8067 14943
rect 10333 14909 10367 14943
rect 24317 14909 24351 14943
rect 25053 14909 25087 14943
rect 33609 14909 33643 14943
rect 35173 14909 35207 14943
rect 38853 14909 38887 14943
rect 7757 14841 7791 14875
rect 13093 14841 13127 14875
rect 16865 14841 16899 14875
rect 19441 14841 19475 14875
rect 22477 14841 22511 14875
rect 37657 14841 37691 14875
rect 4813 14773 4847 14807
rect 7941 14773 7975 14807
rect 9689 14773 9723 14807
rect 10885 14773 10919 14807
rect 17509 14773 17543 14807
rect 23489 14773 23523 14807
rect 24041 14773 24075 14807
rect 24225 14773 24259 14807
rect 25513 14773 25547 14807
rect 27721 14773 27755 14807
rect 29561 14773 29595 14807
rect 3065 14569 3099 14603
rect 3801 14569 3835 14603
rect 14105 14569 14139 14603
rect 17969 14569 18003 14603
rect 23581 14569 23615 14603
rect 24501 14569 24535 14603
rect 25145 14569 25179 14603
rect 30573 14569 30607 14603
rect 40417 14569 40451 14603
rect 28365 14501 28399 14535
rect 18613 14433 18647 14467
rect 20177 14433 20211 14467
rect 21465 14433 21499 14467
rect 26525 14433 26559 14467
rect 26985 14433 27019 14467
rect 35633 14433 35667 14467
rect 38393 14433 38427 14467
rect 3249 14365 3283 14399
rect 3985 14365 4019 14399
rect 9873 14365 9907 14399
rect 12437 14365 12471 14399
rect 15485 14365 15519 14399
rect 16589 14365 16623 14399
rect 16856 14365 16890 14399
rect 19533 14365 19567 14399
rect 19717 14365 19751 14399
rect 20453 14365 20487 14399
rect 22017 14365 22051 14399
rect 22201 14365 22235 14399
rect 22385 14365 22419 14399
rect 23029 14365 23063 14399
rect 23213 14365 23247 14399
rect 23305 14365 23339 14399
rect 23397 14365 23431 14399
rect 29561 14365 29595 14399
rect 35357 14365 35391 14399
rect 36185 14365 36219 14399
rect 40325 14365 40359 14399
rect 58173 14365 58207 14399
rect 15218 14297 15252 14331
rect 22293 14297 22327 14331
rect 26280 14297 26314 14331
rect 27252 14297 27286 14331
rect 32873 14297 32907 14331
rect 7481 14229 7515 14263
rect 9965 14229 9999 14263
rect 12633 14229 12667 14263
rect 19625 14229 19659 14263
rect 22569 14229 22603 14263
rect 31585 14229 31619 14263
rect 37473 14229 37507 14263
rect 3157 14025 3191 14059
rect 8493 14025 8527 14059
rect 23029 14025 23063 14059
rect 23949 14025 23983 14059
rect 24961 14025 24995 14059
rect 27261 14025 27295 14059
rect 31401 14025 31435 14059
rect 39773 14025 39807 14059
rect 14473 13957 14507 13991
rect 19349 13957 19383 13991
rect 22293 13957 22327 13991
rect 24409 13957 24443 13991
rect 28641 13957 28675 13991
rect 28825 13957 28859 13991
rect 29009 13957 29043 13991
rect 30665 13957 30699 13991
rect 35541 13957 35575 13991
rect 39865 13957 39899 13991
rect 2789 13889 2823 13923
rect 2973 13889 3007 13923
rect 6745 13889 6779 13923
rect 14289 13889 14323 13923
rect 18797 13889 18831 13923
rect 19901 13889 19935 13923
rect 20085 13889 20119 13923
rect 20913 13889 20947 13923
rect 23213 13889 23247 13923
rect 23489 13889 23523 13923
rect 24133 13889 24167 13923
rect 26433 13889 26467 13923
rect 27491 13889 27525 13923
rect 27610 13889 27644 13923
rect 27721 13895 27755 13929
rect 27905 13889 27939 13923
rect 29469 13889 29503 13923
rect 29632 13895 29666 13929
rect 29745 13889 29779 13923
rect 29837 13889 29871 13923
rect 30849 13889 30883 13923
rect 34446 13889 34480 13923
rect 34713 13889 34747 13923
rect 35173 13889 35207 13923
rect 35357 13889 35391 13923
rect 36277 13889 36311 13923
rect 38577 13889 38611 13923
rect 38761 13889 38795 13923
rect 38853 13889 38887 13923
rect 38945 13889 38979 13923
rect 6377 13821 6411 13855
rect 6837 13821 6871 13855
rect 7021 13821 7055 13855
rect 20269 13821 20303 13855
rect 23305 13821 23339 13855
rect 24225 13821 24259 13855
rect 30113 13821 30147 13855
rect 36093 13821 36127 13855
rect 37289 13821 37323 13855
rect 37565 13821 37599 13855
rect 20729 13753 20763 13787
rect 14657 13685 14691 13719
rect 23213 13685 23247 13719
rect 24133 13685 24167 13719
rect 33333 13685 33367 13719
rect 36461 13685 36495 13719
rect 39221 13685 39255 13719
rect 5181 13481 5215 13515
rect 11989 13481 12023 13515
rect 14473 13481 14507 13515
rect 21281 13481 21315 13515
rect 22201 13481 22235 13515
rect 27077 13481 27111 13515
rect 28181 13481 28215 13515
rect 29561 13481 29595 13515
rect 33149 13481 33183 13515
rect 37289 13481 37323 13515
rect 38209 13481 38243 13515
rect 18613 13413 18647 13447
rect 20821 13413 20855 13447
rect 2513 13345 2547 13379
rect 5641 13345 5675 13379
rect 5825 13345 5859 13379
rect 8309 13345 8343 13379
rect 8953 13345 8987 13379
rect 23857 13345 23891 13379
rect 26525 13345 26559 13379
rect 30941 13345 30975 13379
rect 32045 13345 32079 13379
rect 2329 13277 2363 13311
rect 6653 13277 6687 13311
rect 9229 13277 9263 13311
rect 11805 13277 11839 13311
rect 14749 13277 14783 13311
rect 14838 13277 14872 13311
rect 14933 13271 14967 13305
rect 15117 13277 15151 13311
rect 17693 13277 17727 13311
rect 19349 13277 19383 13311
rect 20637 13277 20671 13311
rect 23581 13277 23615 13311
rect 24777 13277 24811 13311
rect 27307 13277 27341 13311
rect 27445 13277 27479 13311
rect 27537 13277 27571 13311
rect 27721 13277 27755 13311
rect 32505 13277 32539 13311
rect 32689 13277 32723 13311
rect 32781 13277 32815 13311
rect 32873 13277 32907 13311
rect 35725 13277 35759 13311
rect 36001 13277 36035 13311
rect 36553 13277 36587 13311
rect 36737 13277 36771 13311
rect 38025 13277 38059 13311
rect 58173 13277 58207 13311
rect 15577 13209 15611 13243
rect 17509 13209 17543 13243
rect 19901 13209 19935 13243
rect 20085 13209 20119 13243
rect 30674 13209 30708 13243
rect 37841 13209 37875 13243
rect 2145 13141 2179 13175
rect 4629 13141 4663 13175
rect 5549 13141 5583 13175
rect 17877 13141 17911 13175
rect 33609 13141 33643 13175
rect 36737 13141 36771 13175
rect 4813 12937 4847 12971
rect 6469 12937 6503 12971
rect 10609 12937 10643 12971
rect 21833 12937 21867 12971
rect 23581 12937 23615 12971
rect 24133 12937 24167 12971
rect 32689 12937 32723 12971
rect 35081 12937 35115 12971
rect 40049 12937 40083 12971
rect 13921 12869 13955 12903
rect 14105 12869 14139 12903
rect 14289 12869 14323 12903
rect 24685 12869 24719 12903
rect 32505 12869 32539 12903
rect 35633 12869 35667 12903
rect 37473 12869 37507 12903
rect 37657 12869 37691 12903
rect 38936 12869 38970 12903
rect 2053 12801 2087 12835
rect 2697 12801 2731 12835
rect 2953 12801 2987 12835
rect 5181 12801 5215 12835
rect 5273 12801 5307 12835
rect 8134 12801 8168 12835
rect 8401 12801 8435 12835
rect 9505 12801 9539 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 11713 12801 11747 12835
rect 12081 12801 12115 12835
rect 12265 12801 12299 12835
rect 15025 12801 15059 12835
rect 15117 12801 15151 12835
rect 15209 12801 15243 12835
rect 15393 12801 15427 12835
rect 17897 12801 17931 12835
rect 18153 12801 18187 12835
rect 18889 12801 18923 12835
rect 18978 12801 19012 12835
rect 19073 12801 19107 12835
rect 19257 12801 19291 12835
rect 21005 12801 21039 12835
rect 22937 12801 22971 12835
rect 23489 12801 23523 12835
rect 32321 12801 32355 12835
rect 36093 12801 36127 12835
rect 36256 12801 36290 12835
rect 36369 12801 36403 12835
rect 36507 12801 36541 12835
rect 38669 12801 38703 12835
rect 5365 12733 5399 12767
rect 9321 12733 9355 12767
rect 9689 12733 9723 12767
rect 9781 12733 9815 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 18613 12733 18647 12767
rect 20729 12733 20763 12767
rect 33149 12733 33183 12767
rect 33425 12733 33459 12767
rect 2237 12665 2271 12699
rect 4077 12665 4111 12699
rect 15853 12665 15887 12699
rect 37289 12665 37323 12699
rect 7021 12597 7055 12631
rect 11529 12597 11563 12631
rect 14749 12597 14783 12631
rect 16773 12597 16807 12631
rect 27077 12597 27111 12631
rect 36737 12597 36771 12631
rect 7573 12393 7607 12427
rect 9045 12393 9079 12427
rect 14105 12393 14139 12427
rect 21925 12393 21959 12427
rect 22569 12393 22603 12427
rect 35909 12393 35943 12427
rect 38209 12393 38243 12427
rect 17509 12325 17543 12359
rect 19349 12325 19383 12359
rect 28457 12325 28491 12359
rect 30665 12325 30699 12359
rect 3801 12257 3835 12291
rect 6101 12257 6135 12291
rect 6193 12257 6227 12291
rect 8033 12257 8067 12291
rect 9505 12257 9539 12291
rect 19809 12257 19843 12291
rect 24501 12257 24535 12291
rect 2605 12189 2639 12223
rect 2697 12189 2731 12223
rect 7757 12189 7791 12223
rect 7941 12189 7975 12223
rect 8125 12189 8159 12223
rect 8309 12189 8343 12223
rect 9772 12189 9806 12223
rect 11345 12189 11379 12223
rect 11612 12189 11646 12223
rect 13553 12189 13587 12223
rect 15218 12189 15252 12223
rect 15485 12189 15519 12223
rect 16221 12189 16255 12223
rect 16313 12189 16347 12223
rect 16405 12189 16439 12223
rect 16589 12189 16623 12223
rect 17141 12189 17175 12223
rect 18245 12189 18279 12223
rect 18337 12189 18371 12223
rect 18434 12183 18468 12217
rect 18613 12189 18647 12223
rect 20177 12189 20211 12223
rect 20867 12189 20901 12223
rect 21005 12189 21039 12223
rect 21097 12189 21131 12223
rect 21281 12189 21315 12223
rect 25191 12189 25225 12223
rect 25329 12189 25363 12223
rect 25421 12189 25455 12223
rect 25605 12189 25639 12223
rect 27445 12189 27479 12223
rect 31125 12189 31159 12223
rect 31309 12189 31343 12223
rect 31401 12189 31435 12223
rect 31493 12189 31527 12223
rect 33609 12189 33643 12223
rect 36829 12189 36863 12223
rect 4046 12121 4080 12155
rect 13369 12121 13403 12155
rect 17325 12121 17359 12155
rect 19993 12121 20027 12155
rect 21833 12121 21867 12155
rect 27629 12121 27663 12155
rect 28273 12121 28307 12155
rect 31769 12121 31803 12155
rect 33342 12121 33376 12155
rect 37074 12121 37108 12155
rect 2881 12053 2915 12087
rect 5181 12053 5215 12087
rect 5641 12053 5675 12087
rect 6009 12053 6043 12087
rect 6929 12053 6963 12087
rect 10885 12053 10919 12087
rect 12725 12053 12759 12087
rect 13185 12053 13219 12087
rect 15945 12053 15979 12087
rect 17969 12053 18003 12087
rect 20637 12053 20671 12087
rect 23121 12053 23155 12087
rect 24961 12053 24995 12087
rect 32229 12053 32263 12087
rect 3065 11849 3099 11883
rect 5825 11849 5859 11883
rect 13737 11849 13771 11883
rect 17049 11849 17083 11883
rect 19901 11849 19935 11883
rect 23305 11849 23339 11883
rect 29653 11849 29687 11883
rect 32137 11849 32171 11883
rect 35173 11849 35207 11883
rect 14850 11781 14884 11815
rect 21014 11781 21048 11815
rect 25114 11781 25148 11815
rect 32505 11781 32539 11815
rect 35449 11781 35483 11815
rect 39497 11781 39531 11815
rect 2881 11713 2915 11747
rect 4721 11713 4755 11747
rect 5549 11713 5583 11747
rect 6929 11713 6963 11747
rect 8870 11713 8904 11747
rect 9137 11713 9171 11747
rect 11805 11713 11839 11747
rect 15117 11713 15151 11747
rect 18162 11713 18196 11747
rect 18429 11713 18463 11747
rect 18981 11713 19015 11747
rect 22385 11713 22419 11747
rect 22477 11713 22511 11747
rect 22569 11713 22603 11747
rect 22753 11713 22787 11747
rect 23213 11713 23247 11747
rect 23397 11713 23431 11747
rect 28365 11713 28399 11747
rect 30389 11713 30423 11747
rect 30481 11713 30515 11747
rect 30573 11713 30607 11747
rect 30757 11713 30791 11747
rect 32321 11713 32355 11747
rect 34529 11713 34563 11747
rect 35357 11713 35391 11747
rect 35541 11713 35575 11747
rect 35725 11713 35759 11747
rect 38577 11713 38611 11747
rect 4445 11645 4479 11679
rect 5181 11645 5215 11679
rect 5641 11645 5675 11679
rect 6469 11645 6503 11679
rect 6837 11645 6871 11679
rect 11529 11645 11563 11679
rect 21281 11645 21315 11679
rect 24869 11645 24903 11679
rect 38301 11645 38335 11679
rect 19165 11577 19199 11611
rect 28549 11577 28583 11611
rect 39313 11577 39347 11611
rect 58173 11577 58207 11611
rect 7113 11509 7147 11543
rect 7757 11509 7791 11543
rect 15853 11509 15887 11543
rect 22109 11509 22143 11543
rect 23857 11509 23891 11543
rect 26249 11509 26283 11543
rect 30113 11509 30147 11543
rect 34621 11509 34655 11543
rect 8033 11305 8067 11339
rect 18705 11305 18739 11339
rect 20545 11305 20579 11339
rect 36277 11305 36311 11339
rect 38117 11305 38151 11339
rect 11529 11237 11563 11271
rect 7573 11169 7607 11203
rect 7665 11169 7699 11203
rect 21557 11169 21591 11203
rect 25973 11169 26007 11203
rect 32597 11169 32631 11203
rect 32873 11169 32907 11203
rect 34897 11169 34931 11203
rect 40233 11169 40267 11203
rect 7297 11101 7331 11135
rect 7481 11101 7515 11135
rect 7849 11101 7883 11135
rect 11345 11101 11379 11135
rect 21824 11101 21858 11135
rect 23581 11101 23615 11135
rect 23765 11101 23799 11135
rect 25053 11101 25087 11135
rect 25329 11101 25363 11135
rect 30205 11101 30239 11135
rect 30461 11101 30495 11135
rect 37657 11101 37691 11135
rect 38945 11101 38979 11135
rect 39037 11101 39071 11135
rect 39129 11101 39163 11135
rect 39313 11101 39347 11135
rect 40049 11101 40083 11135
rect 8953 11033 8987 11067
rect 18153 11033 18187 11067
rect 19441 11033 19475 11067
rect 26240 11033 26274 11067
rect 35164 11033 35198 11067
rect 39865 11033 39899 11067
rect 22937 10965 22971 10999
rect 23397 10965 23431 10999
rect 27353 10965 27387 10999
rect 28457 10965 28491 10999
rect 31585 10965 31619 10999
rect 38669 10965 38703 10999
rect 23305 10761 23339 10795
rect 24777 10761 24811 10795
rect 25881 10761 25915 10795
rect 30849 10761 30883 10795
rect 34529 10761 34563 10795
rect 35081 10761 35115 10795
rect 40141 10761 40175 10795
rect 17049 10693 17083 10727
rect 28641 10693 28675 10727
rect 31033 10693 31067 10727
rect 31217 10693 31251 10727
rect 36369 10693 36403 10727
rect 39006 10693 39040 10727
rect 6653 10625 6687 10659
rect 10609 10625 10643 10659
rect 11529 10625 11563 10659
rect 15945 10625 15979 10659
rect 22477 10625 22511 10659
rect 22661 10625 22695 10659
rect 24409 10625 24443 10659
rect 24593 10625 24627 10659
rect 25237 10625 25271 10659
rect 25421 10625 25455 10659
rect 25513 10625 25547 10659
rect 25605 10625 25639 10659
rect 27169 10625 27203 10659
rect 27629 10625 27663 10659
rect 27813 10625 27847 10659
rect 27905 10625 27939 10659
rect 27997 10625 28031 10659
rect 33977 10625 34011 10659
rect 35357 10625 35391 10659
rect 35446 10625 35480 10659
rect 35541 10625 35575 10659
rect 35725 10625 35759 10659
rect 36553 10625 36587 10659
rect 6377 10557 6411 10591
rect 10701 10557 10735 10591
rect 10793 10557 10827 10591
rect 16129 10557 16163 10591
rect 22293 10557 22327 10591
rect 30297 10557 30331 10591
rect 36185 10557 36219 10591
rect 38761 10557 38795 10591
rect 28181 10489 28215 10523
rect 10241 10421 10275 10455
rect 18337 10421 18371 10455
rect 19349 10421 19383 10455
rect 26985 10421 27019 10455
rect 58173 10421 58207 10455
rect 4537 10217 4571 10251
rect 10885 10217 10919 10251
rect 16313 10217 16347 10251
rect 16957 10217 16991 10251
rect 25697 10217 25731 10251
rect 32781 10217 32815 10251
rect 12633 10149 12667 10183
rect 14289 10149 14323 10183
rect 25145 10149 25179 10183
rect 12909 10081 12943 10115
rect 29561 10081 29595 10115
rect 2329 10013 2363 10047
rect 2513 10013 2547 10047
rect 9597 10013 9631 10047
rect 9781 10013 9815 10047
rect 12817 10013 12851 10047
rect 14933 10013 14967 10047
rect 25881 10013 25915 10047
rect 28549 10013 28583 10047
rect 29837 10013 29871 10047
rect 30849 10013 30883 10047
rect 31033 10013 31067 10047
rect 31125 10013 31159 10047
rect 31217 10013 31251 10047
rect 32229 10013 32263 10047
rect 32597 10013 32631 10047
rect 35541 10013 35575 10047
rect 35725 10013 35759 10047
rect 38577 10013 38611 10047
rect 4629 9945 4663 9979
rect 12173 9945 12207 9979
rect 16221 9945 16255 9979
rect 26065 9945 26099 9979
rect 32413 9945 32447 9979
rect 32505 9945 32539 9979
rect 38393 9945 38427 9979
rect 2145 9877 2179 9911
rect 6837 9877 6871 9911
rect 9137 9877 9171 9911
rect 9965 9877 9999 9911
rect 13277 9877 13311 9911
rect 15393 9877 15427 9911
rect 28733 9877 28767 9911
rect 31493 9877 31527 9911
rect 35357 9877 35391 9911
rect 38761 9877 38795 9911
rect 10977 9673 11011 9707
rect 12265 9673 12299 9707
rect 39773 9673 39807 9707
rect 8375 9605 8409 9639
rect 20729 9605 20763 9639
rect 23397 9605 23431 9639
rect 25513 9605 25547 9639
rect 29745 9605 29779 9639
rect 29929 9605 29963 9639
rect 31309 9605 31343 9639
rect 33241 9605 33275 9639
rect 35256 9605 35290 9639
rect 1409 9537 1443 9571
rect 2309 9537 2343 9571
rect 4353 9537 4387 9571
rect 5549 9537 5583 9571
rect 6837 9537 6871 9571
rect 8585 9537 8619 9571
rect 9597 9537 9631 9571
rect 9864 9537 9898 9571
rect 11713 9537 11747 9571
rect 13185 9537 13219 9571
rect 13369 9537 13403 9571
rect 14473 9537 14507 9571
rect 15577 9537 15611 9571
rect 18613 9537 18647 9571
rect 23121 9537 23155 9571
rect 23305 9537 23339 9571
rect 23489 9537 23523 9571
rect 25237 9537 25271 9571
rect 25421 9537 25455 9571
rect 25605 9537 25639 9571
rect 28549 9537 28583 9571
rect 29561 9537 29595 9571
rect 31033 9537 31067 9571
rect 31217 9537 31251 9571
rect 31401 9537 31435 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 32413 9537 32447 9571
rect 32505 9537 32539 9571
rect 38660 9537 38694 9571
rect 2053 9469 2087 9503
rect 5825 9469 5859 9503
rect 8217 9469 8251 9503
rect 21833 9469 21867 9503
rect 22109 9469 22143 9503
rect 28273 9469 28307 9503
rect 30573 9469 30607 9503
rect 34989 9469 35023 9503
rect 38393 9469 38427 9503
rect 1593 9401 1627 9435
rect 7573 9401 7607 9435
rect 11529 9401 11563 9435
rect 15761 9401 15795 9435
rect 23673 9401 23707 9435
rect 25789 9401 25823 9435
rect 31585 9401 31619 9435
rect 3433 9333 3467 9367
rect 4445 9333 4479 9367
rect 6929 9333 6963 9367
rect 8769 9333 8803 9367
rect 13553 9333 13587 9367
rect 14657 9333 14691 9367
rect 18153 9333 18187 9367
rect 18797 9333 18831 9367
rect 32781 9333 32815 9367
rect 36369 9333 36403 9367
rect 37473 9333 37507 9367
rect 2421 9129 2455 9163
rect 13553 9129 13587 9163
rect 18705 9129 18739 9163
rect 20637 9129 20671 9163
rect 27721 9129 27755 9163
rect 30113 9129 30147 9163
rect 31677 9129 31711 9163
rect 32689 9129 32723 9163
rect 34989 9129 35023 9163
rect 6561 9061 6595 9095
rect 11437 9061 11471 9095
rect 14105 9061 14139 9095
rect 3065 8993 3099 9027
rect 5365 8993 5399 9027
rect 6929 8993 6963 9027
rect 8033 8993 8067 9027
rect 12541 8993 12575 9027
rect 12633 8993 12667 9027
rect 15485 8993 15519 9027
rect 21189 8993 21223 9027
rect 21925 8993 21959 9027
rect 28457 8993 28491 9027
rect 4077 8925 4111 8959
rect 4261 8925 4295 8959
rect 5917 8925 5951 8959
rect 6745 8925 6779 8959
rect 7021 8925 7055 8959
rect 7113 8925 7147 8959
rect 7297 8925 7331 8959
rect 10149 8925 10183 8959
rect 13001 8925 13035 8959
rect 16129 8925 16163 8959
rect 17325 8925 17359 8959
rect 19257 8925 19291 8959
rect 21097 8925 21131 8959
rect 21281 8925 21315 8959
rect 22201 8925 22235 8959
rect 27169 8925 27203 8959
rect 27353 8925 27387 8959
rect 27537 8925 27571 8959
rect 28181 8925 28215 8959
rect 29561 8925 29595 8959
rect 29929 8925 29963 8959
rect 31309 8925 31343 8959
rect 32137 8925 32171 8959
rect 32413 8925 32447 8959
rect 32505 8925 32539 8959
rect 35219 8925 35253 8959
rect 35370 8922 35404 8956
rect 35470 8922 35504 8956
rect 35633 8925 35667 8959
rect 36921 8925 36955 8959
rect 37565 8925 37599 8959
rect 58173 8925 58207 8959
rect 2881 8857 2915 8891
rect 5089 8857 5123 8891
rect 8217 8857 8251 8891
rect 9413 8857 9447 8891
rect 9597 8857 9631 8891
rect 15240 8857 15274 8891
rect 17570 8857 17604 8891
rect 19502 8857 19536 8891
rect 27445 8857 27479 8891
rect 29745 8857 29779 8891
rect 29837 8857 29871 8891
rect 31493 8857 31527 8891
rect 32321 8857 32355 8891
rect 36737 8857 36771 8891
rect 1961 8789 1995 8823
rect 2789 8789 2823 8823
rect 3893 8789 3927 8823
rect 4721 8789 4755 8823
rect 5181 8789 5215 8823
rect 6101 8789 6135 8823
rect 12357 8789 12391 8823
rect 15945 8789 15979 8823
rect 16589 8789 16623 8823
rect 24501 8789 24535 8823
rect 37105 8789 37139 8823
rect 38853 8789 38887 8823
rect 4629 8585 4663 8619
rect 5825 8585 5859 8619
rect 6745 8585 6779 8619
rect 7941 8585 7975 8619
rect 9413 8585 9447 8619
rect 10333 8585 10367 8619
rect 13553 8585 13587 8619
rect 14013 8585 14047 8619
rect 15117 8585 15151 8619
rect 17325 8585 17359 8619
rect 19073 8585 19107 8619
rect 21005 8585 21039 8619
rect 28917 8585 28951 8619
rect 29837 8585 29871 8619
rect 32229 8585 32263 8619
rect 38577 8585 38611 8619
rect 16773 8517 16807 8551
rect 19533 8517 19567 8551
rect 19717 8517 19751 8551
rect 23704 8517 23738 8551
rect 24409 8517 24443 8551
rect 26065 8517 26099 8551
rect 28549 8517 28583 8551
rect 28641 8517 28675 8551
rect 34805 8517 34839 8551
rect 2513 8449 2547 8483
rect 2780 8449 2814 8483
rect 5181 8449 5215 8483
rect 6929 8449 6963 8483
rect 7113 8449 7147 8483
rect 8953 8449 8987 8483
rect 10701 8449 10735 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 12081 8449 12115 8483
rect 12265 8449 12299 8483
rect 13921 8449 13955 8483
rect 14933 8449 14967 8483
rect 17601 8449 17635 8483
rect 17693 8449 17727 8483
rect 17785 8449 17819 8483
rect 17969 8449 18003 8483
rect 18429 8449 18463 8483
rect 18613 8449 18647 8483
rect 18705 8449 18739 8483
rect 18843 8449 18877 8483
rect 19901 8449 19935 8483
rect 24685 8449 24719 8483
rect 24777 8449 24811 8483
rect 24869 8449 24903 8483
rect 25053 8449 25087 8483
rect 26249 8449 26283 8483
rect 28365 8449 28399 8483
rect 28733 8449 28767 8483
rect 31125 8449 31159 8483
rect 36645 8449 36679 8483
rect 37473 8449 37507 8483
rect 37636 8452 37670 8486
rect 37749 8449 37783 8483
rect 37887 8449 37921 8483
rect 38853 8449 38887 8483
rect 38945 8449 38979 8483
rect 39037 8449 39071 8483
rect 39221 8449 39255 8483
rect 39681 8449 39715 8483
rect 5549 8381 5583 8415
rect 5641 8381 5675 8415
rect 8033 8381 8067 8415
rect 8217 8381 8251 8415
rect 10793 8381 10827 8415
rect 11989 8381 12023 8415
rect 14105 8381 14139 8415
rect 23949 8381 23983 8415
rect 1501 8313 1535 8347
rect 2053 8313 2087 8347
rect 3893 8313 3927 8347
rect 7573 8313 7607 8347
rect 10977 8313 11011 8347
rect 13001 8313 13035 8347
rect 11529 8245 11563 8279
rect 16037 8245 16071 8279
rect 22569 8245 22603 8279
rect 25881 8245 25915 8279
rect 38117 8245 38151 8279
rect 1593 8041 1627 8075
rect 3801 8041 3835 8075
rect 4905 8041 4939 8075
rect 7849 8041 7883 8075
rect 17693 8041 17727 8075
rect 18245 8041 18279 8075
rect 19257 8041 19291 8075
rect 23213 8041 23247 8075
rect 24777 8041 24811 8075
rect 27077 8041 27111 8075
rect 30205 8041 30239 8075
rect 34989 8041 35023 8075
rect 36093 8041 36127 8075
rect 37289 8041 37323 8075
rect 39313 8041 39347 8075
rect 16957 7973 16991 8007
rect 6469 7905 6503 7939
rect 12449 7905 12483 7939
rect 25697 7905 25731 7939
rect 37933 7905 37967 7939
rect 3985 7837 4019 7871
rect 6725 7837 6759 7871
rect 10241 7837 10275 7871
rect 12265 7837 12299 7871
rect 12532 7837 12566 7871
rect 12629 7837 12663 7871
rect 12817 7837 12851 7871
rect 14565 7837 14599 7871
rect 15577 7837 15611 7871
rect 19441 7837 19475 7871
rect 21005 7837 21039 7871
rect 21189 7837 21223 7871
rect 22661 7837 22695 7871
rect 22937 7837 22971 7871
rect 23029 7837 23063 7871
rect 24593 7837 24627 7871
rect 31329 7837 31363 7871
rect 31585 7837 31619 7871
rect 35173 7837 35207 7871
rect 35265 7837 35299 7871
rect 35541 7837 35575 7871
rect 38200 7837 38234 7871
rect 58173 7837 58207 7871
rect 2145 7769 2179 7803
rect 5457 7769 5491 7803
rect 9505 7769 9539 7803
rect 10508 7769 10542 7803
rect 15822 7769 15856 7803
rect 19625 7769 19659 7803
rect 21097 7769 21131 7803
rect 22845 7769 22879 7803
rect 24409 7769 24443 7803
rect 25964 7769 25998 7803
rect 35357 7769 35391 7803
rect 2697 7701 2731 7735
rect 3249 7701 3283 7735
rect 6009 7701 6043 7735
rect 8401 7701 8435 7735
rect 8953 7701 8987 7735
rect 11621 7701 11655 7735
rect 12081 7701 12115 7735
rect 13461 7701 13495 7735
rect 14657 7701 14691 7735
rect 21649 7701 21683 7735
rect 3893 7497 3927 7531
rect 7757 7497 7791 7531
rect 9873 7497 9907 7531
rect 11713 7497 11747 7531
rect 12449 7497 12483 7531
rect 15209 7497 15243 7531
rect 20361 7497 20395 7531
rect 22937 7497 22971 7531
rect 26065 7497 26099 7531
rect 27169 7497 27203 7531
rect 36001 7497 36035 7531
rect 10885 7429 10919 7463
rect 15117 7429 15151 7463
rect 16865 7429 16899 7463
rect 22661 7429 22695 7463
rect 24133 7429 24167 7463
rect 28457 7429 28491 7463
rect 30573 7429 30607 7463
rect 33618 7429 33652 7463
rect 36369 7429 36403 7463
rect 38853 7429 38887 7463
rect 5549 7361 5583 7395
rect 8125 7361 8159 7395
rect 8217 7361 8251 7395
rect 11529 7361 11563 7395
rect 17049 7361 17083 7395
rect 18061 7361 18095 7395
rect 19533 7361 19567 7395
rect 20913 7361 20947 7395
rect 21097 7361 21131 7395
rect 22385 7361 22419 7395
rect 22569 7361 22603 7395
rect 22753 7361 22787 7395
rect 24317 7361 24351 7395
rect 25421 7361 25455 7395
rect 25605 7361 25639 7395
rect 25697 7361 25731 7395
rect 25789 7361 25823 7395
rect 26985 7361 27019 7395
rect 28273 7361 28307 7395
rect 30757 7361 30791 7395
rect 33885 7361 33919 7395
rect 35127 7361 35161 7395
rect 35265 7361 35299 7395
rect 35357 7361 35391 7395
rect 35541 7361 35575 7395
rect 36185 7361 36219 7395
rect 36277 7361 36311 7395
rect 36553 7361 36587 7395
rect 38669 7361 38703 7395
rect 2329 7293 2363 7327
rect 5825 7293 5859 7327
rect 6469 7293 6503 7327
rect 6745 7293 6779 7327
rect 18337 7293 18371 7327
rect 8861 7225 8895 7259
rect 13277 7225 13311 7259
rect 16129 7225 16163 7259
rect 21281 7225 21315 7259
rect 32505 7225 32539 7259
rect 1777 7157 1811 7191
rect 2881 7157 2915 7191
rect 3433 7157 3467 7191
rect 4537 7157 4571 7191
rect 8401 7157 8435 7191
rect 10333 7157 10367 7191
rect 13829 7157 13863 7191
rect 14381 7157 14415 7191
rect 16681 7157 16715 7191
rect 17601 7157 17635 7191
rect 19349 7157 19383 7191
rect 23489 7157 23523 7191
rect 23949 7157 23983 7191
rect 24961 7157 24995 7191
rect 28089 7157 28123 7191
rect 30389 7157 30423 7191
rect 34345 7157 34379 7191
rect 34897 7157 34931 7191
rect 39037 7157 39071 7191
rect 15393 6953 15427 6987
rect 27629 6953 27663 6987
rect 31401 6953 31435 6987
rect 36921 6953 36955 6987
rect 2513 6817 2547 6851
rect 9229 6817 9263 6851
rect 14933 6817 14967 6851
rect 16957 6817 16991 6851
rect 22201 6817 22235 6851
rect 25789 6817 25823 6851
rect 29009 6817 29043 6851
rect 30021 6817 30055 6851
rect 36461 6817 36495 6851
rect 2329 6749 2363 6783
rect 3985 6749 4019 6783
rect 4169 6749 4203 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 6469 6749 6503 6783
rect 7297 6749 7331 6783
rect 8125 6749 8159 6783
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 9321 6749 9355 6783
rect 9505 6749 9539 6783
rect 12826 6749 12860 6783
rect 13093 6749 13127 6783
rect 15669 6749 15703 6783
rect 15761 6749 15795 6783
rect 15853 6749 15887 6783
rect 16037 6749 16071 6783
rect 17969 6749 18003 6783
rect 21925 6749 21959 6783
rect 23469 6749 23503 6783
rect 23581 6749 23615 6783
rect 23673 6749 23707 6783
rect 23857 6749 23891 6783
rect 24409 6749 24443 6783
rect 24593 6749 24627 6783
rect 24685 6749 24719 6783
rect 24777 6749 24811 6783
rect 26065 6749 26099 6783
rect 34069 6749 34103 6783
rect 34943 6749 34977 6783
rect 35081 6749 35115 6783
rect 35194 6749 35228 6783
rect 35357 6749 35391 6783
rect 35817 6749 35851 6783
rect 36001 6749 36035 6783
rect 36093 6749 36127 6783
rect 36185 6749 36219 6783
rect 38761 6749 38795 6783
rect 38853 6749 38887 6783
rect 38945 6749 38979 6783
rect 39129 6749 39163 6783
rect 1685 6681 1719 6715
rect 5457 6681 5491 6715
rect 10701 6681 10735 6715
rect 19441 6681 19475 6715
rect 28742 6681 28776 6715
rect 30288 6681 30322 6715
rect 37105 6681 37139 6715
rect 37289 6681 37323 6715
rect 38025 6681 38059 6715
rect 39865 6681 39899 6715
rect 2145 6613 2179 6647
rect 3249 6613 3283 6647
rect 3801 6613 3835 6647
rect 5549 6613 5583 6647
rect 6653 6613 6687 6647
rect 7481 6613 7515 6647
rect 7941 6613 7975 6647
rect 9689 6613 9723 6647
rect 11253 6613 11287 6647
rect 11713 6613 11747 6647
rect 14381 6613 14415 6647
rect 18429 6613 18463 6647
rect 19993 6613 20027 6647
rect 20729 6613 20763 6647
rect 21189 6613 21223 6647
rect 23213 6613 23247 6647
rect 25053 6613 25087 6647
rect 27077 6613 27111 6647
rect 34713 6613 34747 6647
rect 38485 6613 38519 6647
rect 6469 6409 6503 6443
rect 15301 6409 15335 6443
rect 23673 6409 23707 6443
rect 24225 6409 24259 6443
rect 25145 6409 25179 6443
rect 27537 6409 27571 6443
rect 29193 6409 29227 6443
rect 30389 6409 30423 6443
rect 36093 6409 36127 6443
rect 39681 6409 39715 6443
rect 3249 6341 3283 6375
rect 4997 6341 5031 6375
rect 12357 6341 12391 6375
rect 15945 6341 15979 6375
rect 17049 6341 17083 6375
rect 23305 6341 23339 6375
rect 23397 6341 23431 6375
rect 26433 6341 26467 6375
rect 31033 6341 31067 6375
rect 34958 6341 34992 6375
rect 36553 6341 36587 6375
rect 1501 6273 1535 6307
rect 2789 6273 2823 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 7113 6273 7147 6307
rect 7941 6273 7975 6307
rect 8401 6273 8435 6307
rect 9137 6273 9171 6307
rect 9404 6273 9438 6307
rect 13921 6273 13955 6307
rect 14188 6273 14222 6307
rect 16129 6273 16163 6307
rect 19441 6273 19475 6307
rect 19625 6273 19659 6307
rect 22109 6273 22143 6307
rect 23121 6273 23155 6307
rect 23489 6273 23523 6307
rect 26985 6273 27019 6307
rect 27813 6273 27847 6307
rect 27905 6273 27939 6307
rect 27997 6273 28031 6307
rect 28181 6273 28215 6307
rect 29745 6273 29779 6307
rect 29929 6276 29963 6310
rect 30024 6276 30058 6310
rect 30133 6273 30167 6307
rect 31217 6273 31251 6307
rect 34713 6273 34747 6307
rect 38301 6273 38335 6307
rect 38568 6273 38602 6307
rect 18797 6205 18831 6239
rect 21833 6205 21867 6239
rect 7297 6137 7331 6171
rect 11805 6137 11839 6171
rect 58173 6137 58207 6171
rect 1685 6069 1719 6103
rect 2237 6069 2271 6103
rect 5641 6069 5675 6103
rect 7757 6069 7791 6103
rect 8585 6069 8619 6103
rect 10517 6069 10551 6103
rect 12909 6069 12943 6103
rect 13461 6069 13495 6103
rect 15761 6069 15795 6103
rect 19257 6069 19291 6103
rect 20269 6069 20303 6103
rect 20821 6069 20855 6103
rect 30849 6069 30883 6103
rect 3985 5865 4019 5899
rect 14473 5865 14507 5899
rect 20637 5865 20671 5899
rect 24409 5865 24443 5899
rect 33885 5865 33919 5899
rect 34989 5865 35023 5899
rect 36001 5865 36035 5899
rect 3249 5797 3283 5831
rect 6929 5797 6963 5831
rect 31585 5797 31619 5831
rect 4261 5729 4295 5763
rect 4629 5729 4663 5763
rect 1869 5661 1903 5695
rect 4169 5661 4203 5695
rect 5457 5661 5491 5695
rect 5641 5661 5675 5695
rect 6101 5661 6135 5695
rect 6193 5661 6227 5695
rect 7389 5661 7423 5695
rect 8125 5661 8159 5695
rect 9137 5661 9171 5695
rect 9781 5661 9815 5695
rect 10425 5661 10459 5695
rect 11069 5661 11103 5695
rect 11713 5661 11747 5695
rect 12541 5661 12575 5695
rect 13369 5661 13403 5695
rect 14749 5661 14783 5695
rect 14841 5661 14875 5695
rect 14933 5661 14967 5695
rect 15117 5661 15151 5695
rect 16681 5661 16715 5695
rect 16957 5661 16991 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 18337 5661 18371 5695
rect 18429 5661 18463 5695
rect 19257 5661 19291 5695
rect 25605 5661 25639 5695
rect 25881 5661 25915 5695
rect 27721 5661 27755 5695
rect 30113 5661 30147 5695
rect 30297 5661 30331 5695
rect 30392 5661 30426 5695
rect 30481 5661 30515 5695
rect 32413 5661 32447 5695
rect 35173 5661 35207 5695
rect 36185 5661 36219 5695
rect 36369 5661 36403 5695
rect 2114 5593 2148 5627
rect 6377 5593 6411 5627
rect 16037 5593 16071 5627
rect 16221 5593 16255 5627
rect 18705 5593 18739 5627
rect 19502 5593 19536 5627
rect 24593 5593 24627 5627
rect 24777 5593 24811 5627
rect 27537 5593 27571 5627
rect 31217 5593 31251 5627
rect 31401 5593 31435 5627
rect 35357 5593 35391 5627
rect 5549 5525 5583 5559
rect 6101 5525 6135 5559
rect 7573 5525 7607 5559
rect 8309 5525 8343 5559
rect 8953 5525 8987 5559
rect 9597 5525 9631 5559
rect 15853 5525 15887 5559
rect 21649 5525 21683 5559
rect 22201 5525 22235 5559
rect 22661 5525 22695 5559
rect 23213 5525 23247 5559
rect 27353 5525 27387 5559
rect 29561 5525 29595 5559
rect 30757 5525 30791 5559
rect 2421 5321 2455 5355
rect 2881 5321 2915 5355
rect 4537 5321 4571 5355
rect 4997 5321 5031 5355
rect 5181 5321 5215 5355
rect 12725 5321 12759 5355
rect 25421 5321 25455 5355
rect 29745 5321 29779 5355
rect 32229 5321 32263 5355
rect 37289 5321 37323 5355
rect 5733 5253 5767 5287
rect 6377 5253 6411 5287
rect 8401 5253 8435 5287
rect 19349 5253 19383 5287
rect 19717 5253 19751 5287
rect 26433 5253 26467 5287
rect 2789 5185 2823 5219
rect 3709 5185 3743 5219
rect 4353 5185 4387 5219
rect 6561 5185 6595 5219
rect 6745 5185 6779 5219
rect 7573 5185 7607 5219
rect 9045 5185 9079 5219
rect 12633 5185 12667 5219
rect 12817 5185 12851 5219
rect 14565 5185 14599 5219
rect 15301 5185 15335 5219
rect 15485 5185 15519 5219
rect 15577 5185 15611 5219
rect 15669 5185 15703 5219
rect 18245 5185 18279 5219
rect 18429 5185 18463 5219
rect 18521 5185 18555 5219
rect 18613 5185 18647 5219
rect 19533 5185 19567 5219
rect 27261 5185 27295 5219
rect 27353 5185 27387 5219
rect 27445 5185 27479 5219
rect 27629 5185 27663 5219
rect 30205 5185 30239 5219
rect 30389 5185 30423 5219
rect 30481 5185 30515 5219
rect 30593 5185 30627 5219
rect 38402 5185 38436 5219
rect 38669 5185 38703 5219
rect 3065 5117 3099 5151
rect 5273 5117 5307 5151
rect 7481 5117 7515 5151
rect 8033 5117 8067 5151
rect 54401 5117 54435 5151
rect 5733 5049 5767 5083
rect 8861 5049 8895 5083
rect 15945 5049 15979 5083
rect 18889 5049 18923 5083
rect 23305 5049 23339 5083
rect 55045 5049 55079 5083
rect 1961 4981 1995 5015
rect 3893 4981 3927 5015
rect 7941 4981 7975 5015
rect 9689 4981 9723 5015
rect 10333 4981 10367 5015
rect 10977 4981 11011 5015
rect 11989 4981 12023 5015
rect 13461 4981 13495 5015
rect 14105 4981 14139 5015
rect 14749 4981 14783 5015
rect 16865 4981 16899 5015
rect 17785 4981 17819 5015
rect 20177 4981 20211 5015
rect 21005 4981 21039 5015
rect 21833 4981 21867 5015
rect 22661 4981 22695 5015
rect 23857 4981 23891 5015
rect 26985 4981 27019 5015
rect 30849 4981 30883 5015
rect 53757 4981 53791 5015
rect 58173 4981 58207 5015
rect 6101 4777 6135 4811
rect 7481 4777 7515 4811
rect 7757 4777 7791 4811
rect 8953 4777 8987 4811
rect 9413 4777 9447 4811
rect 10241 4777 10275 4811
rect 22477 4777 22511 4811
rect 24409 4777 24443 4811
rect 2329 4709 2363 4743
rect 4997 4709 5031 4743
rect 8401 4709 8435 4743
rect 10609 4709 10643 4743
rect 16773 4709 16807 4743
rect 21373 4709 21407 4743
rect 32413 4709 32447 4743
rect 52837 4709 52871 4743
rect 55321 4709 55355 4743
rect 4353 4641 4387 4675
rect 7481 4641 7515 4675
rect 9045 4641 9079 4675
rect 10517 4641 10551 4675
rect 12909 4641 12943 4675
rect 18061 4641 18095 4675
rect 54125 4641 54159 4675
rect 55965 4641 55999 4675
rect 2973 4573 3007 4607
rect 3985 4573 4019 4607
rect 4169 4573 4203 4607
rect 5181 4573 5215 4607
rect 5641 4573 5675 4607
rect 6009 4573 6043 4607
rect 6193 4573 6227 4607
rect 7113 4573 7147 4607
rect 7573 4573 7607 4607
rect 9229 4573 9263 4607
rect 10738 4573 10772 4607
rect 11621 4573 11655 4607
rect 12265 4573 12299 4607
rect 13369 4573 13403 4607
rect 14841 4573 14875 4607
rect 15485 4573 15519 4607
rect 16129 4573 16163 4607
rect 17417 4573 17451 4607
rect 18705 4573 18739 4607
rect 19441 4573 19475 4607
rect 20085 4573 20119 4607
rect 20729 4573 20763 4607
rect 22017 4573 22051 4607
rect 23590 4573 23624 4607
rect 23857 4573 23891 4607
rect 25789 4573 25823 4607
rect 31033 4573 31067 4607
rect 31289 4573 31323 4607
rect 52193 4573 52227 4607
rect 53481 4573 53515 4607
rect 1777 4505 1811 4539
rect 8953 4505 8987 4539
rect 10885 4505 10919 4539
rect 25522 4505 25556 4539
rect 2789 4437 2823 4471
rect 5825 4437 5859 4471
rect 13553 4437 13587 4471
rect 14197 4437 14231 4471
rect 6745 4233 6779 4267
rect 6377 4165 6411 4199
rect 6561 4165 6595 4199
rect 27252 4165 27286 4199
rect 2605 4097 2639 4131
rect 3525 4097 3559 4131
rect 4077 4097 4111 4131
rect 4261 4097 4295 4131
rect 4997 4097 5031 4131
rect 5825 4097 5859 4131
rect 7849 4097 7883 4131
rect 9505 4097 9539 4131
rect 10057 4097 10091 4131
rect 11713 4097 11747 4131
rect 12081 4097 12115 4131
rect 13369 4097 13403 4131
rect 16681 4097 16715 4131
rect 16948 4097 16982 4131
rect 19533 4097 19567 4131
rect 19789 4097 19823 4131
rect 26985 4097 27019 4131
rect 34621 4097 34655 4131
rect 34877 4097 34911 4131
rect 54677 4097 54711 4131
rect 5733 4029 5767 4063
rect 8401 4029 8435 4063
rect 8585 4029 8619 4063
rect 10425 4029 10459 4063
rect 10977 4029 11011 4063
rect 11621 4029 11655 4063
rect 14841 4029 14875 4063
rect 52745 4029 52779 4063
rect 55965 4029 55999 4063
rect 8309 3961 8343 3995
rect 10609 3961 10643 3995
rect 12909 3961 12943 3995
rect 14197 3961 14231 3995
rect 15485 3961 15519 3995
rect 18061 3961 18095 3995
rect 20913 3961 20947 3995
rect 24961 3961 24995 3995
rect 28365 3961 28399 3995
rect 36001 3961 36035 3995
rect 1593 3893 1627 3927
rect 2145 3893 2179 3927
rect 2789 3893 2823 3927
rect 3341 3893 3375 3927
rect 4813 3893 4847 3927
rect 5457 3893 5491 3927
rect 5825 3893 5859 3927
rect 6561 3893 6595 3927
rect 7389 3893 7423 3927
rect 8217 3893 8251 3927
rect 9321 3893 9355 3927
rect 10517 3893 10551 3927
rect 12081 3893 12115 3927
rect 12265 3893 12299 3927
rect 13553 3893 13587 3927
rect 16129 3893 16163 3927
rect 19073 3893 19107 3927
rect 22385 3893 22419 3927
rect 23029 3893 23063 3927
rect 23489 3893 23523 3927
rect 24317 3893 24351 3927
rect 25513 3893 25547 3927
rect 51181 3893 51215 3927
rect 51825 3893 51859 3927
rect 53389 3893 53423 3927
rect 54033 3893 54067 3927
rect 55321 3893 55355 3927
rect 58173 3893 58207 3927
rect 7941 3689 7975 3723
rect 9045 3689 9079 3723
rect 9781 3689 9815 3723
rect 10701 3689 10735 3723
rect 12909 3689 12943 3723
rect 17049 3689 17083 3723
rect 18613 3689 18647 3723
rect 20269 3689 20303 3723
rect 21097 3689 21131 3723
rect 21925 3689 21959 3723
rect 32321 3689 32355 3723
rect 3801 3621 3835 3655
rect 7481 3621 7515 3655
rect 7849 3621 7883 3655
rect 10885 3621 10919 3655
rect 10977 3621 11011 3655
rect 13553 3621 13587 3655
rect 14197 3621 14231 3655
rect 16221 3621 16255 3655
rect 17877 3621 17911 3655
rect 46949 3621 46983 3655
rect 52837 3621 52871 3655
rect 55321 3621 55355 3655
rect 6193 3553 6227 3587
rect 8033 3553 8067 3587
rect 8401 3553 8435 3587
rect 10793 3553 10827 3587
rect 12265 3553 12299 3587
rect 14749 3553 14783 3587
rect 19625 3553 19659 3587
rect 30941 3553 30975 3587
rect 51549 3553 51583 3587
rect 53481 3553 53515 3587
rect 56609 3553 56643 3587
rect 1869 3485 1903 3519
rect 5181 3485 5215 3519
rect 6469 3485 6503 3519
rect 9229 3485 9263 3519
rect 9965 3485 9999 3519
rect 11345 3485 11379 3519
rect 13369 3485 13403 3519
rect 14657 3485 14691 3519
rect 16037 3485 16071 3519
rect 16865 3485 16899 3519
rect 17693 3485 17727 3519
rect 18429 3485 18463 3519
rect 20085 3485 20119 3519
rect 20913 3485 20947 3519
rect 21741 3485 21775 3519
rect 23213 3485 23247 3519
rect 23857 3485 23891 3519
rect 24869 3485 24903 3519
rect 25697 3485 25731 3519
rect 26801 3485 26835 3519
rect 27629 3485 27663 3519
rect 28733 3485 28767 3519
rect 31197 3485 31231 3519
rect 34805 3485 34839 3519
rect 35449 3485 35483 3519
rect 36093 3485 36127 3519
rect 36737 3485 36771 3519
rect 37565 3485 37599 3519
rect 38669 3485 38703 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 41337 3485 41371 3519
rect 42533 3485 42567 3519
rect 43177 3485 43211 3519
rect 45017 3485 45051 3519
rect 45661 3485 45695 3519
rect 46305 3485 46339 3519
rect 47777 3485 47811 3519
rect 48421 3485 48455 3519
rect 50261 3485 50295 3519
rect 50905 3485 50939 3519
rect 52193 3485 52227 3519
rect 54125 3485 54159 3519
rect 55965 3485 55999 3519
rect 57529 3485 57563 3519
rect 58173 3485 58207 3519
rect 2136 3417 2170 3451
rect 4936 3417 4970 3451
rect 5733 3417 5767 3451
rect 14197 3417 14231 3451
rect 3249 3349 3283 3383
rect 14933 3349 14967 3383
rect 15485 3349 15519 3383
rect 22569 3349 22603 3383
rect 3801 3145 3835 3179
rect 5667 3145 5701 3179
rect 8309 3145 8343 3179
rect 11621 3145 11655 3179
rect 14473 3145 14507 3179
rect 18245 3145 18279 3179
rect 18889 3145 18923 3179
rect 20361 3145 20395 3179
rect 21097 3145 21131 3179
rect 23029 3145 23063 3179
rect 1961 3077 1995 3111
rect 2688 3077 2722 3111
rect 5457 3077 5491 3111
rect 15117 3077 15151 3111
rect 16129 3077 16163 3111
rect 17601 3077 17635 3111
rect 20453 3077 20487 3111
rect 1777 3009 1811 3043
rect 2421 3009 2455 3043
rect 4997 3009 5031 3043
rect 6561 3009 6595 3043
rect 6837 3009 6871 3043
rect 8033 3009 8067 3043
rect 8953 3009 8987 3043
rect 9873 3009 9907 3043
rect 10701 3009 10735 3043
rect 11805 3009 11839 3043
rect 13921 3009 13955 3043
rect 14565 3009 14599 3043
rect 15301 3009 15335 3043
rect 15945 3009 15979 3043
rect 17417 3009 17451 3043
rect 18061 3009 18095 3043
rect 19073 3009 19107 3043
rect 19809 3009 19843 3043
rect 21281 3009 21315 3043
rect 22109 3009 22143 3043
rect 22845 3009 22879 3043
rect 54033 3009 54067 3043
rect 54677 3009 54711 3043
rect 55321 3009 55355 3043
rect 13277 2941 13311 2975
rect 23857 2941 23891 2975
rect 33425 2941 33459 2975
rect 39221 2941 39255 2975
rect 43085 2941 43119 2975
rect 55965 2941 55999 2975
rect 56609 2941 56643 2975
rect 10885 2873 10919 2907
rect 12633 2873 12667 2907
rect 19625 2873 19659 2907
rect 34713 2873 34747 2907
rect 37933 2873 37967 2907
rect 39865 2873 39899 2907
rect 41153 2873 41187 2907
rect 43729 2873 43763 2907
rect 45017 2873 45051 2907
rect 45661 2873 45695 2907
rect 48237 2873 48271 2907
rect 49525 2873 49559 2907
rect 50813 2873 50847 2907
rect 52745 2873 52779 2907
rect 57897 2873 57931 2907
rect 4813 2805 4847 2839
rect 5641 2805 5675 2839
rect 5825 2805 5859 2839
rect 9229 2805 9263 2839
rect 9965 2805 9999 2839
rect 16865 2805 16899 2839
rect 22293 2805 22327 2839
rect 24501 2805 24535 2839
rect 25145 2805 25179 2839
rect 25789 2805 25823 2839
rect 26433 2805 26467 2839
rect 27629 2805 27663 2839
rect 28089 2805 28123 2839
rect 28917 2805 28951 2839
rect 29561 2805 29595 2839
rect 30021 2805 30055 2839
rect 30665 2805 30699 2839
rect 32137 2805 32171 2839
rect 32781 2805 32815 2839
rect 34069 2805 34103 2839
rect 35357 2805 35391 2839
rect 36001 2805 36035 2839
rect 37289 2805 37323 2839
rect 38577 2805 38611 2839
rect 40509 2805 40543 2839
rect 42441 2805 42475 2839
rect 44373 2805 44407 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48881 2805 48915 2839
rect 50169 2805 50203 2839
rect 51457 2805 51491 2839
rect 53389 2805 53423 2839
rect 1593 2601 1627 2635
rect 12357 2601 12391 2635
rect 13553 2601 13587 2635
rect 17141 2601 17175 2635
rect 17785 2601 17819 2635
rect 21097 2601 21131 2635
rect 37289 2601 37323 2635
rect 55321 2601 55355 2635
rect 2421 2533 2455 2567
rect 3157 2533 3191 2567
rect 11713 2533 11747 2567
rect 14381 2533 14415 2567
rect 15393 2533 15427 2567
rect 18521 2533 18555 2567
rect 19809 2533 19843 2567
rect 22017 2533 22051 2567
rect 22753 2533 22787 2567
rect 23581 2533 23615 2567
rect 25789 2533 25823 2567
rect 27721 2533 27755 2567
rect 39865 2533 39899 2567
rect 43729 2533 43763 2567
rect 47593 2533 47627 2567
rect 51457 2533 51491 2567
rect 54033 2533 54067 2567
rect 56609 2533 56643 2567
rect 7205 2465 7239 2499
rect 8401 2465 8435 2499
rect 32781 2465 32815 2499
rect 34713 2465 34747 2499
rect 38577 2465 38611 2499
rect 40509 2465 40543 2499
rect 42441 2465 42475 2499
rect 45017 2465 45051 2499
rect 48237 2465 48271 2499
rect 50169 2465 50203 2499
rect 53389 2465 53423 2499
rect 57897 2465 57931 2499
rect 1777 2397 1811 2431
rect 2237 2397 2271 2431
rect 2973 2397 3007 2431
rect 4077 2397 4111 2431
rect 5089 2397 5123 2431
rect 5825 2397 5859 2431
rect 6929 2397 6963 2431
rect 11529 2397 11563 2431
rect 12541 2397 12575 2431
rect 14197 2397 14231 2431
rect 15853 2397 15887 2431
rect 16957 2397 16991 2431
rect 17969 2397 18003 2431
rect 18705 2397 18739 2431
rect 20545 2397 20579 2431
rect 21281 2397 21315 2431
rect 22201 2397 22235 2431
rect 22937 2397 22971 2431
rect 23397 2397 23431 2431
rect 24409 2397 24443 2431
rect 25145 2397 25179 2431
rect 26433 2397 26467 2431
rect 28365 2397 28399 2431
rect 29009 2397 29043 2431
rect 30113 2397 30147 2431
rect 30757 2397 30791 2431
rect 31217 2397 31251 2431
rect 32137 2397 32171 2431
rect 33425 2397 33459 2431
rect 35357 2397 35391 2431
rect 36001 2397 36035 2431
rect 37933 2397 37967 2431
rect 41153 2397 41187 2431
rect 43085 2397 43119 2431
rect 45661 2397 45695 2431
rect 46305 2397 46339 2431
rect 48881 2397 48915 2431
rect 50813 2397 50847 2431
rect 52745 2397 52779 2431
rect 55965 2397 55999 2431
rect 6469 2329 6503 2363
rect 9045 2329 9079 2363
rect 10149 2329 10183 2363
rect 15209 2329 15243 2363
rect 19625 2329 19659 2363
rect 4261 2261 4295 2295
rect 4905 2261 4939 2295
rect 5641 2261 5675 2295
rect 9321 2261 9355 2295
rect 10425 2261 10459 2295
rect 16037 2261 16071 2295
rect 20361 2261 20395 2295
rect 26985 2261 27019 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 12710 57536 12716 57588
rect 12768 57576 12774 57588
rect 12897 57579 12955 57585
rect 12897 57576 12909 57579
rect 12768 57548 12909 57576
rect 12768 57536 12774 57548
rect 12897 57545 12909 57548
rect 12943 57545 12955 57579
rect 12897 57539 12955 57545
rect 14274 57536 14280 57588
rect 14332 57576 14338 57588
rect 14461 57579 14519 57585
rect 14461 57576 14473 57579
rect 14332 57548 14473 57576
rect 14332 57536 14338 57548
rect 14461 57545 14473 57548
rect 14507 57545 14519 57579
rect 14461 57539 14519 57545
rect 15838 57536 15844 57588
rect 15896 57576 15902 57588
rect 16853 57579 16911 57585
rect 16853 57576 16865 57579
rect 15896 57548 16865 57576
rect 15896 57536 15902 57548
rect 16853 57545 16865 57548
rect 16899 57545 16911 57579
rect 16853 57539 16911 57545
rect 17402 57536 17408 57588
rect 17460 57576 17466 57588
rect 17681 57579 17739 57585
rect 17681 57576 17693 57579
rect 17460 57548 17693 57576
rect 17460 57536 17466 57548
rect 17681 57545 17693 57548
rect 17727 57545 17739 57579
rect 17681 57539 17739 57545
rect 19334 57536 19340 57588
rect 19392 57576 19398 57588
rect 19429 57579 19487 57585
rect 19429 57576 19441 57579
rect 19392 57548 19441 57576
rect 19392 57536 19398 57548
rect 19429 57545 19441 57548
rect 19475 57545 19487 57579
rect 19429 57539 19487 57545
rect 20714 57536 20720 57588
rect 20772 57576 20778 57588
rect 20809 57579 20867 57585
rect 20809 57576 20821 57579
rect 20772 57548 20821 57576
rect 20772 57536 20778 57548
rect 20809 57545 20821 57548
rect 20855 57545 20867 57579
rect 20809 57539 20867 57545
rect 22094 57536 22100 57588
rect 22152 57576 22158 57588
rect 22373 57579 22431 57585
rect 22373 57576 22385 57579
rect 22152 57548 22385 57576
rect 22152 57536 22158 57548
rect 22373 57545 22385 57548
rect 22419 57545 22431 57579
rect 22373 57539 22431 57545
rect 23658 57536 23664 57588
rect 23716 57576 23722 57588
rect 24581 57579 24639 57585
rect 24581 57576 24593 57579
rect 23716 57548 24593 57576
rect 23716 57536 23722 57548
rect 24581 57545 24593 57548
rect 24627 57545 24639 57579
rect 24581 57539 24639 57545
rect 25222 57536 25228 57588
rect 25280 57576 25286 57588
rect 25501 57579 25559 57585
rect 25501 57576 25513 57579
rect 25280 57548 25513 57576
rect 25280 57536 25286 57548
rect 25501 57545 25513 57548
rect 25547 57545 25559 57579
rect 25501 57539 25559 57545
rect 26786 57536 26792 57588
rect 26844 57576 26850 57588
rect 27157 57579 27215 57585
rect 27157 57576 27169 57579
rect 26844 57548 27169 57576
rect 26844 57536 26850 57548
rect 27157 57545 27169 57548
rect 27203 57545 27215 57579
rect 27157 57539 27215 57545
rect 28350 57536 28356 57588
rect 28408 57576 28414 57588
rect 28629 57579 28687 57585
rect 28629 57576 28641 57579
rect 28408 57548 28641 57576
rect 28408 57536 28414 57548
rect 28629 57545 28641 57548
rect 28675 57545 28687 57579
rect 28629 57539 28687 57545
rect 29914 57536 29920 57588
rect 29972 57576 29978 57588
rect 30193 57579 30251 57585
rect 30193 57576 30205 57579
rect 29972 57548 30205 57576
rect 29972 57536 29978 57548
rect 30193 57545 30205 57548
rect 30239 57545 30251 57579
rect 30193 57539 30251 57545
rect 31478 57536 31484 57588
rect 31536 57576 31542 57588
rect 32309 57579 32367 57585
rect 32309 57576 32321 57579
rect 31536 57548 32321 57576
rect 31536 57536 31542 57548
rect 32309 57545 32321 57548
rect 32355 57545 32367 57579
rect 32309 57539 32367 57545
rect 33134 57536 33140 57588
rect 33192 57576 33198 57588
rect 33321 57579 33379 57585
rect 33321 57576 33333 57579
rect 33192 57548 33333 57576
rect 33192 57536 33198 57548
rect 33321 57545 33333 57548
rect 33367 57545 33379 57579
rect 33321 57539 33379 57545
rect 34606 57536 34612 57588
rect 34664 57576 34670 57588
rect 34885 57579 34943 57585
rect 34885 57576 34897 57579
rect 34664 57548 34897 57576
rect 34664 57536 34670 57548
rect 34885 57545 34897 57548
rect 34931 57545 34943 57579
rect 34885 57539 34943 57545
rect 36170 57536 36176 57588
rect 36228 57576 36234 57588
rect 36449 57579 36507 57585
rect 36449 57576 36461 57579
rect 36228 57548 36461 57576
rect 36228 57536 36234 57548
rect 36449 57545 36461 57548
rect 36495 57545 36507 57579
rect 36449 57539 36507 57545
rect 37734 57536 37740 57588
rect 37792 57576 37798 57588
rect 38013 57579 38071 57585
rect 38013 57576 38025 57579
rect 37792 57548 38025 57576
rect 37792 57536 37798 57548
rect 38013 57545 38025 57548
rect 38059 57545 38071 57579
rect 38013 57539 38071 57545
rect 39298 57536 39304 57588
rect 39356 57576 39362 57588
rect 40037 57579 40095 57585
rect 40037 57576 40049 57579
rect 39356 57548 40049 57576
rect 39356 57536 39362 57548
rect 40037 57545 40049 57548
rect 40083 57545 40095 57579
rect 40037 57539 40095 57545
rect 40862 57536 40868 57588
rect 40920 57576 40926 57588
rect 41141 57579 41199 57585
rect 41141 57576 41153 57579
rect 40920 57548 41153 57576
rect 40920 57536 40926 57548
rect 41141 57545 41153 57548
rect 41187 57545 41199 57579
rect 41141 57539 41199 57545
rect 42426 57536 42432 57588
rect 42484 57576 42490 57588
rect 42705 57579 42763 57585
rect 42705 57576 42717 57579
rect 42484 57548 42717 57576
rect 42484 57536 42490 57548
rect 42705 57545 42717 57548
rect 42751 57545 42763 57579
rect 42705 57539 42763 57545
rect 44174 57536 44180 57588
rect 44232 57576 44238 57588
rect 44269 57579 44327 57585
rect 44269 57576 44281 57579
rect 44232 57548 44281 57576
rect 44232 57536 44238 57548
rect 44269 57545 44281 57548
rect 44315 57545 44327 57579
rect 44269 57539 44327 57545
rect 45554 57536 45560 57588
rect 45612 57576 45618 57588
rect 45833 57579 45891 57585
rect 45833 57576 45845 57579
rect 45612 57548 45845 57576
rect 45612 57536 45618 57548
rect 45833 57545 45845 57548
rect 45879 57545 45891 57579
rect 45833 57539 45891 57545
rect 47118 57536 47124 57588
rect 47176 57576 47182 57588
rect 47765 57579 47823 57585
rect 47765 57576 47777 57579
rect 47176 57548 47777 57576
rect 47176 57536 47182 57548
rect 47765 57545 47777 57548
rect 47811 57545 47823 57579
rect 47765 57539 47823 57545
rect 48682 57536 48688 57588
rect 48740 57576 48746 57588
rect 48961 57579 49019 57585
rect 48961 57576 48973 57579
rect 48740 57548 48973 57576
rect 48740 57536 48746 57548
rect 48961 57545 48973 57548
rect 49007 57545 49019 57579
rect 48961 57539 49019 57545
rect 50154 57536 50160 57588
rect 50212 57576 50218 57588
rect 50525 57579 50583 57585
rect 50525 57576 50537 57579
rect 50212 57548 50537 57576
rect 50212 57536 50218 57548
rect 50525 57545 50537 57548
rect 50571 57545 50583 57579
rect 50525 57539 50583 57545
rect 51810 57536 51816 57588
rect 51868 57576 51874 57588
rect 52089 57579 52147 57585
rect 52089 57576 52101 57579
rect 51868 57548 52101 57576
rect 51868 57536 51874 57548
rect 52089 57545 52101 57548
rect 52135 57545 52147 57579
rect 52089 57539 52147 57545
rect 53374 57536 53380 57588
rect 53432 57576 53438 57588
rect 53653 57579 53711 57585
rect 53653 57576 53665 57579
rect 53432 57548 53665 57576
rect 53432 57536 53438 57548
rect 53653 57545 53665 57548
rect 53699 57545 53711 57579
rect 53653 57539 53711 57545
rect 54938 57536 54944 57588
rect 54996 57576 55002 57588
rect 55493 57579 55551 57585
rect 55493 57576 55505 57579
rect 54996 57548 55505 57576
rect 54996 57536 55002 57548
rect 55493 57545 55505 57548
rect 55539 57545 55551 57579
rect 55493 57539 55551 57545
rect 56594 57536 56600 57588
rect 56652 57576 56658 57588
rect 56781 57579 56839 57585
rect 56781 57576 56793 57579
rect 56652 57548 56793 57576
rect 56652 57536 56658 57548
rect 56781 57545 56793 57548
rect 56827 57545 56839 57579
rect 58066 57576 58072 57588
rect 58027 57548 58072 57576
rect 56781 57539 56839 57545
rect 58066 57536 58072 57548
rect 58124 57536 58130 57588
rect 20898 57468 20904 57520
rect 20956 57508 20962 57520
rect 20956 57480 26234 57508
rect 20956 57468 20962 57480
rect 1762 57400 1768 57452
rect 1820 57440 1826 57452
rect 1857 57443 1915 57449
rect 1857 57440 1869 57443
rect 1820 57412 1869 57440
rect 1820 57400 1826 57412
rect 1857 57409 1869 57412
rect 1903 57409 1915 57443
rect 1857 57403 1915 57409
rect 3326 57400 3332 57452
rect 3384 57440 3390 57452
rect 3789 57443 3847 57449
rect 3789 57440 3801 57443
rect 3384 57412 3801 57440
rect 3384 57400 3390 57412
rect 3789 57409 3801 57412
rect 3835 57409 3847 57443
rect 3789 57403 3847 57409
rect 4890 57400 4896 57452
rect 4948 57440 4954 57452
rect 4985 57443 5043 57449
rect 4985 57440 4997 57443
rect 4948 57412 4997 57440
rect 4948 57400 4954 57412
rect 4985 57409 4997 57412
rect 5031 57409 5043 57443
rect 4985 57403 5043 57409
rect 6454 57400 6460 57452
rect 6512 57440 6518 57452
rect 6549 57443 6607 57449
rect 6549 57440 6561 57443
rect 6512 57412 6561 57440
rect 6512 57400 6518 57412
rect 6549 57409 6561 57412
rect 6595 57409 6607 57443
rect 6549 57403 6607 57409
rect 8018 57400 8024 57452
rect 8076 57440 8082 57452
rect 8113 57443 8171 57449
rect 8113 57440 8125 57443
rect 8076 57412 8125 57440
rect 8076 57400 8082 57412
rect 8113 57409 8125 57412
rect 8159 57409 8171 57443
rect 9674 57440 9680 57452
rect 9635 57412 9680 57440
rect 8113 57403 8171 57409
rect 9674 57400 9680 57412
rect 9732 57400 9738 57452
rect 11146 57400 11152 57452
rect 11204 57440 11210 57452
rect 11517 57443 11575 57449
rect 11517 57440 11529 57443
rect 11204 57412 11529 57440
rect 11204 57400 11210 57412
rect 11517 57409 11529 57412
rect 11563 57409 11575 57443
rect 13078 57440 13084 57452
rect 13039 57412 13084 57440
rect 11517 57403 11575 57409
rect 13078 57400 13084 57412
rect 13136 57400 13142 57452
rect 14642 57440 14648 57452
rect 14603 57412 14648 57440
rect 14642 57400 14648 57412
rect 14700 57400 14706 57452
rect 16666 57440 16672 57452
rect 16627 57412 16672 57440
rect 16666 57400 16672 57412
rect 16724 57400 16730 57452
rect 17494 57440 17500 57452
rect 17455 57412 17500 57440
rect 17494 57400 17500 57412
rect 17552 57400 17558 57452
rect 19242 57440 19248 57452
rect 19203 57412 19248 57440
rect 19242 57400 19248 57412
rect 19300 57400 19306 57452
rect 20622 57440 20628 57452
rect 20583 57412 20628 57440
rect 20622 57400 20628 57412
rect 20680 57400 20686 57452
rect 22186 57440 22192 57452
rect 22147 57412 22192 57440
rect 22186 57400 22192 57412
rect 22244 57400 22250 57452
rect 24394 57440 24400 57452
rect 24355 57412 24400 57440
rect 24394 57400 24400 57412
rect 24452 57400 24458 57452
rect 25317 57443 25375 57449
rect 25317 57409 25329 57443
rect 25363 57409 25375 57443
rect 26206 57440 26234 57480
rect 31754 57468 31760 57520
rect 31812 57508 31818 57520
rect 31812 57480 35894 57508
rect 31812 57468 31818 57480
rect 26973 57443 27031 57449
rect 26973 57440 26985 57443
rect 26206 57412 26985 57440
rect 25317 57403 25375 57409
rect 26973 57409 26985 57412
rect 27019 57409 27031 57443
rect 28442 57440 28448 57452
rect 28403 57412 28448 57440
rect 26973 57403 27031 57409
rect 19334 57332 19340 57384
rect 19392 57372 19398 57384
rect 25332 57372 25360 57403
rect 28442 57400 28448 57412
rect 28500 57400 28506 57452
rect 28994 57400 29000 57452
rect 29052 57440 29058 57452
rect 30009 57443 30067 57449
rect 30009 57440 30021 57443
rect 29052 57412 30021 57440
rect 29052 57400 29058 57412
rect 30009 57409 30021 57412
rect 30055 57409 30067 57443
rect 32122 57440 32128 57452
rect 32083 57412 32128 57440
rect 30009 57403 30067 57409
rect 32122 57400 32128 57412
rect 32180 57400 32186 57452
rect 33134 57440 33140 57452
rect 33095 57412 33140 57440
rect 33134 57400 33140 57412
rect 33192 57400 33198 57452
rect 34698 57440 34704 57452
rect 34659 57412 34704 57440
rect 34698 57400 34704 57412
rect 34756 57400 34762 57452
rect 35866 57440 35894 57480
rect 46198 57468 46204 57520
rect 46256 57508 46262 57520
rect 46256 57480 50384 57508
rect 46256 57468 46262 57480
rect 36265 57443 36323 57449
rect 36265 57440 36277 57443
rect 35866 57412 36277 57440
rect 36265 57409 36277 57412
rect 36311 57409 36323 57443
rect 37826 57440 37832 57452
rect 37787 57412 37832 57440
rect 36265 57403 36323 57409
rect 37826 57400 37832 57412
rect 37884 57400 37890 57452
rect 39850 57440 39856 57452
rect 39811 57412 39856 57440
rect 39850 57400 39856 57412
rect 39908 57400 39914 57452
rect 40957 57443 41015 57449
rect 40957 57409 40969 57443
rect 41003 57409 41015 57443
rect 42518 57440 42524 57452
rect 42479 57412 42524 57440
rect 40957 57403 41015 57409
rect 40770 57372 40776 57384
rect 19392 57344 25360 57372
rect 26206 57344 40776 57372
rect 19392 57332 19398 57344
rect 22278 57196 22284 57248
rect 22336 57236 22342 57248
rect 26206 57236 26234 57344
rect 40770 57332 40776 57344
rect 40828 57372 40834 57384
rect 40972 57372 41000 57403
rect 42518 57400 42524 57412
rect 42576 57400 42582 57452
rect 44082 57440 44088 57452
rect 44043 57412 44088 57440
rect 44082 57400 44088 57412
rect 44140 57400 44146 57452
rect 44174 57400 44180 57452
rect 44232 57440 44238 57452
rect 45649 57443 45707 57449
rect 45649 57440 45661 57443
rect 44232 57412 45661 57440
rect 44232 57400 44238 57412
rect 45649 57409 45661 57412
rect 45695 57409 45707 57443
rect 47578 57440 47584 57452
rect 47539 57412 47584 57440
rect 45649 57403 45707 57409
rect 47578 57400 47584 57412
rect 47636 57400 47642 57452
rect 47670 57400 47676 57452
rect 47728 57440 47734 57452
rect 50356 57449 50384 57480
rect 48777 57443 48835 57449
rect 48777 57440 48789 57443
rect 47728 57412 48789 57440
rect 47728 57400 47734 57412
rect 48777 57409 48789 57412
rect 48823 57409 48835 57443
rect 48777 57403 48835 57409
rect 50341 57443 50399 57449
rect 50341 57409 50353 57443
rect 50387 57409 50399 57443
rect 50341 57403 50399 57409
rect 51905 57443 51963 57449
rect 51905 57409 51917 57443
rect 51951 57409 51963 57443
rect 53466 57440 53472 57452
rect 53427 57412 53472 57440
rect 51905 57403 51963 57409
rect 40828 57344 41000 57372
rect 40828 57332 40834 57344
rect 48314 57332 48320 57384
rect 48372 57372 48378 57384
rect 51920 57372 51948 57403
rect 53466 57400 53472 57412
rect 53524 57400 53530 57452
rect 55306 57440 55312 57452
rect 55267 57412 55312 57440
rect 55306 57400 55312 57412
rect 55364 57400 55370 57452
rect 56042 57400 56048 57452
rect 56100 57440 56106 57452
rect 56597 57443 56655 57449
rect 56597 57440 56609 57443
rect 56100 57412 56609 57440
rect 56100 57400 56106 57412
rect 56597 57409 56609 57412
rect 56643 57409 56655 57443
rect 56597 57403 56655 57409
rect 57790 57400 57796 57452
rect 57848 57440 57854 57452
rect 57885 57443 57943 57449
rect 57885 57440 57897 57443
rect 57848 57412 57897 57440
rect 57848 57400 57854 57412
rect 57885 57409 57897 57412
rect 57931 57409 57943 57443
rect 57885 57403 57943 57409
rect 48372 57344 51948 57372
rect 48372 57332 48378 57344
rect 56042 57236 56048 57248
rect 22336 57208 26234 57236
rect 56003 57208 56048 57236
rect 22336 57196 22342 57208
rect 56042 57196 56048 57208
rect 56100 57196 56106 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 21082 56992 21088 57044
rect 21140 57032 21146 57044
rect 40770 57032 40776 57044
rect 21140 57004 26234 57032
rect 40731 57004 40776 57032
rect 21140 56992 21146 57004
rect 26206 56964 26234 57004
rect 40770 56992 40776 57004
rect 40828 56992 40834 57044
rect 57514 57032 57520 57044
rect 57475 57004 57520 57032
rect 57514 56992 57520 57004
rect 57572 56992 57578 57044
rect 42337 56967 42395 56973
rect 42337 56964 42349 56967
rect 26206 56936 42349 56964
rect 42337 56933 42349 56936
rect 42383 56964 42395 56967
rect 42518 56964 42524 56976
rect 42383 56936 42524 56964
rect 42383 56933 42395 56936
rect 42337 56927 42395 56933
rect 42518 56924 42524 56936
rect 42576 56924 42582 56976
rect 57882 56788 57888 56840
rect 57940 56828 57946 56840
rect 58161 56831 58219 56837
rect 58161 56828 58173 56831
rect 57940 56800 58173 56828
rect 57940 56788 57946 56800
rect 58161 56797 58173 56800
rect 58207 56797 58219 56831
rect 58161 56791 58219 56797
rect 16117 56695 16175 56701
rect 16117 56661 16129 56695
rect 16163 56692 16175 56695
rect 16482 56692 16488 56704
rect 16163 56664 16488 56692
rect 16163 56661 16175 56664
rect 16117 56655 16175 56661
rect 16482 56652 16488 56664
rect 16540 56652 16546 56704
rect 28074 56692 28080 56704
rect 28035 56664 28080 56692
rect 28074 56652 28080 56664
rect 28132 56652 28138 56704
rect 29178 56652 29184 56704
rect 29236 56692 29242 56704
rect 29549 56695 29607 56701
rect 29549 56692 29561 56695
rect 29236 56664 29561 56692
rect 29236 56652 29242 56664
rect 29549 56661 29561 56664
rect 29595 56661 29607 56695
rect 29549 56655 29607 56661
rect 45373 56695 45431 56701
rect 45373 56661 45385 56695
rect 45419 56692 45431 56695
rect 45462 56692 45468 56704
rect 45419 56664 45468 56692
rect 45419 56661 45431 56664
rect 45373 56655 45431 56661
rect 45462 56652 45468 56664
rect 45520 56652 45526 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 13078 56448 13084 56500
rect 13136 56488 13142 56500
rect 13725 56491 13783 56497
rect 13725 56488 13737 56491
rect 13136 56460 13737 56488
rect 13136 56448 13142 56460
rect 13725 56457 13737 56460
rect 13771 56457 13783 56491
rect 13725 56451 13783 56457
rect 14642 56448 14648 56500
rect 14700 56488 14706 56500
rect 14829 56491 14887 56497
rect 14829 56488 14841 56491
rect 14700 56460 14841 56488
rect 14700 56448 14706 56460
rect 14829 56457 14841 56460
rect 14875 56457 14887 56491
rect 14829 56451 14887 56457
rect 15933 56491 15991 56497
rect 15933 56457 15945 56491
rect 15979 56488 15991 56491
rect 16666 56488 16672 56500
rect 15979 56460 16672 56488
rect 15979 56457 15991 56460
rect 15933 56451 15991 56457
rect 16666 56448 16672 56460
rect 16724 56448 16730 56500
rect 16853 56491 16911 56497
rect 16853 56457 16865 56491
rect 16899 56488 16911 56491
rect 17494 56488 17500 56500
rect 16899 56460 17500 56488
rect 16899 56457 16911 56460
rect 16853 56451 16911 56457
rect 17494 56448 17500 56460
rect 17552 56448 17558 56500
rect 18141 56491 18199 56497
rect 18141 56457 18153 56491
rect 18187 56457 18199 56491
rect 18141 56451 18199 56457
rect 18785 56491 18843 56497
rect 18785 56457 18797 56491
rect 18831 56488 18843 56491
rect 20622 56488 20628 56500
rect 18831 56460 20628 56488
rect 18831 56457 18843 56460
rect 18785 56451 18843 56457
rect 18156 56420 18184 56451
rect 20622 56448 20628 56460
rect 20680 56448 20686 56500
rect 22278 56488 22284 56500
rect 22239 56460 22284 56488
rect 22278 56448 22284 56460
rect 22336 56448 22342 56500
rect 23293 56491 23351 56497
rect 23293 56457 23305 56491
rect 23339 56488 23351 56491
rect 24394 56488 24400 56500
rect 23339 56460 24400 56488
rect 23339 56457 23351 56460
rect 23293 56451 23351 56457
rect 24394 56448 24400 56460
rect 24452 56448 24458 56500
rect 27801 56491 27859 56497
rect 27801 56457 27813 56491
rect 27847 56488 27859 56491
rect 28442 56488 28448 56500
rect 27847 56460 28448 56488
rect 27847 56457 27859 56460
rect 27801 56451 27859 56457
rect 28442 56448 28448 56460
rect 28500 56448 28506 56500
rect 30377 56491 30435 56497
rect 30377 56457 30389 56491
rect 30423 56488 30435 56491
rect 32122 56488 32128 56500
rect 30423 56460 32128 56488
rect 30423 56457 30435 56460
rect 30377 56451 30435 56457
rect 32122 56448 32128 56460
rect 32180 56448 32186 56500
rect 32309 56491 32367 56497
rect 32309 56457 32321 56491
rect 32355 56488 32367 56491
rect 33134 56488 33140 56500
rect 32355 56460 33140 56488
rect 32355 56457 32367 56460
rect 32309 56451 32367 56457
rect 33134 56448 33140 56460
rect 33192 56448 33198 56500
rect 33781 56491 33839 56497
rect 33781 56457 33793 56491
rect 33827 56488 33839 56491
rect 34698 56488 34704 56500
rect 33827 56460 34704 56488
rect 33827 56457 33839 56460
rect 33781 56451 33839 56457
rect 34698 56448 34704 56460
rect 34756 56448 34762 56500
rect 35989 56491 36047 56497
rect 35989 56457 36001 56491
rect 36035 56488 36047 56491
rect 37826 56488 37832 56500
rect 36035 56460 37832 56488
rect 36035 56457 36047 56460
rect 35989 56451 36047 56457
rect 37826 56448 37832 56460
rect 37884 56448 37890 56500
rect 43073 56491 43131 56497
rect 43073 56457 43085 56491
rect 43119 56457 43131 56491
rect 43073 56451 43131 56457
rect 43717 56491 43775 56497
rect 43717 56457 43729 56491
rect 43763 56488 43775 56491
rect 44174 56488 44180 56500
rect 43763 56460 44180 56488
rect 43763 56457 43775 56460
rect 43717 56451 43775 56457
rect 19334 56420 19340 56432
rect 18156 56392 19340 56420
rect 19334 56380 19340 56392
rect 19392 56380 19398 56432
rect 21082 56420 21088 56432
rect 21043 56392 21088 56420
rect 21082 56380 21088 56392
rect 21140 56380 21146 56432
rect 28074 56420 28080 56432
rect 26206 56392 28080 56420
rect 13909 56355 13967 56361
rect 13909 56321 13921 56355
rect 13955 56352 13967 56355
rect 14182 56352 14188 56364
rect 13955 56324 14188 56352
rect 13955 56321 13967 56324
rect 13909 56315 13967 56321
rect 14182 56312 14188 56324
rect 14240 56312 14246 56364
rect 15013 56355 15071 56361
rect 15013 56321 15025 56355
rect 15059 56352 15071 56355
rect 15102 56352 15108 56364
rect 15059 56324 15108 56352
rect 15059 56321 15071 56324
rect 15013 56315 15071 56321
rect 15102 56312 15108 56324
rect 15160 56312 15166 56364
rect 15749 56355 15807 56361
rect 15749 56321 15761 56355
rect 15795 56352 15807 56355
rect 16482 56352 16488 56364
rect 15795 56324 16488 56352
rect 15795 56321 15807 56324
rect 15749 56315 15807 56321
rect 16482 56312 16488 56324
rect 16540 56312 16546 56364
rect 16574 56312 16580 56364
rect 16632 56352 16638 56364
rect 16669 56355 16727 56361
rect 16669 56352 16681 56355
rect 16632 56324 16681 56352
rect 16632 56312 16638 56324
rect 16669 56321 16681 56324
rect 16715 56321 16727 56355
rect 16669 56315 16727 56321
rect 17218 56312 17224 56364
rect 17276 56352 17282 56364
rect 17313 56355 17371 56361
rect 17313 56352 17325 56355
rect 17276 56324 17325 56352
rect 17276 56312 17282 56324
rect 17313 56321 17325 56324
rect 17359 56321 17371 56355
rect 17313 56315 17371 56321
rect 17862 56312 17868 56364
rect 17920 56352 17926 56364
rect 17957 56355 18015 56361
rect 17957 56352 17969 56355
rect 17920 56324 17969 56352
rect 17920 56312 17926 56324
rect 17957 56321 17969 56324
rect 18003 56321 18015 56355
rect 18598 56352 18604 56364
rect 18559 56324 18604 56352
rect 17957 56315 18015 56321
rect 18598 56312 18604 56324
rect 18656 56312 18662 56364
rect 19058 56312 19064 56364
rect 19116 56352 19122 56364
rect 19245 56355 19303 56361
rect 19245 56352 19257 56355
rect 19116 56324 19257 56352
rect 19116 56312 19122 56324
rect 19245 56321 19257 56324
rect 19291 56321 19303 56355
rect 19245 56315 19303 56321
rect 20346 56312 20352 56364
rect 20404 56352 20410 56364
rect 20901 56355 20959 56361
rect 20901 56352 20913 56355
rect 20404 56324 20913 56352
rect 20404 56312 20410 56324
rect 20901 56321 20913 56324
rect 20947 56321 20959 56355
rect 20901 56315 20959 56321
rect 21910 56312 21916 56364
rect 21968 56352 21974 56364
rect 22097 56355 22155 56361
rect 22097 56352 22109 56355
rect 21968 56324 22109 56352
rect 21968 56312 21974 56324
rect 22097 56321 22109 56324
rect 22143 56321 22155 56355
rect 23106 56352 23112 56364
rect 23067 56324 23112 56352
rect 22097 56315 22155 56321
rect 23106 56312 23112 56324
rect 23164 56352 23170 56364
rect 23753 56355 23811 56361
rect 23753 56352 23765 56355
rect 23164 56324 23765 56352
rect 23164 56312 23170 56324
rect 23753 56321 23765 56324
rect 23799 56321 23811 56355
rect 23753 56315 23811 56321
rect 20162 56244 20168 56296
rect 20220 56284 20226 56296
rect 26206 56284 26234 56392
rect 28074 56380 28080 56392
rect 28132 56420 28138 56432
rect 43088 56420 43116 56451
rect 44174 56448 44180 56460
rect 44232 56448 44238 56500
rect 45005 56491 45063 56497
rect 45005 56457 45017 56491
rect 45051 56488 45063 56491
rect 46198 56488 46204 56500
rect 45051 56460 46204 56488
rect 45051 56457 45063 56460
rect 45005 56451 45063 56457
rect 46198 56448 46204 56460
rect 46256 56448 46262 56500
rect 46293 56491 46351 56497
rect 46293 56457 46305 56491
rect 46339 56488 46351 56491
rect 47578 56488 47584 56500
rect 46339 56460 47584 56488
rect 46339 56457 46351 56460
rect 46293 56451 46351 56457
rect 47578 56448 47584 56460
rect 47636 56448 47642 56500
rect 53466 56420 53472 56432
rect 28132 56392 28304 56420
rect 43088 56392 53472 56420
rect 28132 56380 28138 56392
rect 28276 56361 28304 56392
rect 53466 56380 53472 56392
rect 53524 56380 53530 56432
rect 27617 56355 27675 56361
rect 27617 56352 27629 56355
rect 20220 56256 26234 56284
rect 27080 56324 27629 56352
rect 20220 56244 20226 56256
rect 17497 56219 17555 56225
rect 17497 56185 17509 56219
rect 17543 56216 17555 56219
rect 19242 56216 19248 56228
rect 17543 56188 19248 56216
rect 17543 56185 17555 56188
rect 17497 56179 17555 56185
rect 19242 56176 19248 56188
rect 19300 56176 19306 56228
rect 19429 56219 19487 56225
rect 19429 56185 19441 56219
rect 19475 56216 19487 56219
rect 20898 56216 20904 56228
rect 19475 56188 20904 56216
rect 19475 56185 19487 56188
rect 19429 56179 19487 56185
rect 20898 56176 20904 56188
rect 20956 56176 20962 56228
rect 20346 56148 20352 56160
rect 20307 56120 20352 56148
rect 20346 56108 20352 56120
rect 20404 56108 20410 56160
rect 23566 56108 23572 56160
rect 23624 56148 23630 56160
rect 27080 56157 27108 56324
rect 27617 56321 27629 56324
rect 27663 56321 27675 56355
rect 27617 56315 27675 56321
rect 28261 56355 28319 56361
rect 28261 56321 28273 56355
rect 28307 56321 28319 56355
rect 29178 56352 29184 56364
rect 29139 56324 29184 56352
rect 28261 56315 28319 56321
rect 29178 56312 29184 56324
rect 29236 56312 29242 56364
rect 30006 56312 30012 56364
rect 30064 56352 30070 56364
rect 30193 56355 30251 56361
rect 30193 56352 30205 56355
rect 30064 56324 30205 56352
rect 30064 56312 30070 56324
rect 30193 56321 30205 56324
rect 30239 56321 30251 56355
rect 30193 56315 30251 56321
rect 30834 56312 30840 56364
rect 30892 56352 30898 56364
rect 31389 56355 31447 56361
rect 31389 56352 31401 56355
rect 30892 56324 31401 56352
rect 30892 56312 30898 56324
rect 31389 56321 31401 56324
rect 31435 56321 31447 56355
rect 32122 56352 32128 56364
rect 32083 56324 32128 56352
rect 31389 56315 31447 56321
rect 32122 56312 32128 56324
rect 32180 56352 32186 56364
rect 32769 56355 32827 56361
rect 32769 56352 32781 56355
rect 32180 56324 32781 56352
rect 32180 56312 32186 56324
rect 32769 56321 32781 56324
rect 32815 56321 32827 56355
rect 33594 56352 33600 56364
rect 33555 56324 33600 56352
rect 32769 56315 32827 56321
rect 33594 56312 33600 56324
rect 33652 56352 33658 56364
rect 34241 56355 34299 56361
rect 34241 56352 34253 56355
rect 33652 56324 34253 56352
rect 33652 56312 33658 56324
rect 34241 56321 34253 56324
rect 34287 56321 34299 56355
rect 35802 56352 35808 56364
rect 35715 56324 35808 56352
rect 34241 56315 34299 56321
rect 35802 56312 35808 56324
rect 35860 56352 35866 56364
rect 36449 56355 36507 56361
rect 36449 56352 36461 56355
rect 35860 56324 36461 56352
rect 35860 56312 35866 56324
rect 36449 56321 36461 56324
rect 36495 56321 36507 56355
rect 42886 56352 42892 56364
rect 42847 56324 42892 56352
rect 36449 56315 36507 56321
rect 42886 56312 42892 56324
rect 42944 56312 42950 56364
rect 43530 56352 43536 56364
rect 43491 56324 43536 56352
rect 43530 56312 43536 56324
rect 43588 56312 43594 56364
rect 43990 56312 43996 56364
rect 44048 56352 44054 56364
rect 44177 56355 44235 56361
rect 44177 56352 44189 56355
rect 44048 56324 44189 56352
rect 44048 56312 44054 56324
rect 44177 56321 44189 56324
rect 44223 56321 44235 56355
rect 44177 56315 44235 56321
rect 44726 56312 44732 56364
rect 44784 56352 44790 56364
rect 44821 56355 44879 56361
rect 44821 56352 44833 56355
rect 44784 56324 44833 56352
rect 44784 56312 44790 56324
rect 44821 56321 44833 56324
rect 44867 56321 44879 56355
rect 45462 56352 45468 56364
rect 45423 56324 45468 56352
rect 44821 56315 44879 56321
rect 45462 56312 45468 56324
rect 45520 56312 45526 56364
rect 46106 56352 46112 56364
rect 46067 56324 46112 56352
rect 46106 56312 46112 56324
rect 46164 56312 46170 56364
rect 46750 56352 46756 56364
rect 46711 56324 46756 56352
rect 46750 56312 46756 56324
rect 46808 56312 46814 56364
rect 58161 56355 58219 56361
rect 58161 56321 58173 56355
rect 58207 56352 58219 56355
rect 58434 56352 58440 56364
rect 58207 56324 58440 56352
rect 58207 56321 58219 56324
rect 58161 56315 58219 56321
rect 58434 56312 58440 56324
rect 58492 56312 58498 56364
rect 55306 56284 55312 56296
rect 45526 56256 55312 56284
rect 28445 56219 28503 56225
rect 28445 56185 28457 56219
rect 28491 56216 28503 56219
rect 28994 56216 29000 56228
rect 28491 56188 29000 56216
rect 28491 56185 28503 56188
rect 28445 56179 28503 56185
rect 28994 56176 29000 56188
rect 29052 56176 29058 56228
rect 29365 56219 29423 56225
rect 29365 56185 29377 56219
rect 29411 56216 29423 56219
rect 44082 56216 44088 56228
rect 29411 56188 44088 56216
rect 29411 56185 29423 56188
rect 29365 56179 29423 56185
rect 44082 56176 44088 56188
rect 44140 56176 44146 56228
rect 44361 56219 44419 56225
rect 44361 56185 44373 56219
rect 44407 56216 44419 56219
rect 45526 56216 45554 56256
rect 55306 56244 55312 56256
rect 55364 56244 55370 56296
rect 44407 56188 45554 56216
rect 46937 56219 46995 56225
rect 44407 56185 44419 56188
rect 44361 56179 44419 56185
rect 46937 56185 46949 56219
rect 46983 56216 46995 56219
rect 48314 56216 48320 56228
rect 46983 56188 48320 56216
rect 46983 56185 46995 56188
rect 46937 56179 46995 56185
rect 48314 56176 48320 56188
rect 48372 56176 48378 56228
rect 27065 56151 27123 56157
rect 27065 56148 27077 56151
rect 23624 56120 27077 56148
rect 23624 56108 23630 56120
rect 27065 56117 27077 56120
rect 27111 56117 27123 56151
rect 30834 56148 30840 56160
rect 30795 56120 30840 56148
rect 27065 56111 27123 56117
rect 30834 56108 30840 56120
rect 30892 56108 30898 56160
rect 31573 56151 31631 56157
rect 31573 56117 31585 56151
rect 31619 56148 31631 56151
rect 31754 56148 31760 56160
rect 31619 56120 31760 56148
rect 31619 56117 31631 56120
rect 31573 56111 31631 56117
rect 31754 56108 31760 56120
rect 31812 56108 31818 56160
rect 45649 56151 45707 56157
rect 45649 56117 45661 56151
rect 45695 56148 45707 56151
rect 47670 56148 47676 56160
rect 45695 56120 47676 56148
rect 45695 56117 45707 56120
rect 45649 56111 45707 56117
rect 47670 56108 47676 56120
rect 47728 56108 47734 56160
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 17862 55944 17868 55956
rect 17823 55916 17868 55944
rect 17862 55904 17868 55916
rect 17920 55904 17926 55956
rect 21177 55947 21235 55953
rect 21177 55913 21189 55947
rect 21223 55944 21235 55947
rect 22186 55944 22192 55956
rect 21223 55916 22192 55944
rect 21223 55913 21235 55916
rect 21177 55907 21235 55913
rect 22186 55904 22192 55916
rect 22244 55904 22250 55956
rect 20993 55743 21051 55749
rect 20993 55740 21005 55743
rect 20456 55712 21005 55740
rect 16390 55632 16396 55684
rect 16448 55672 16454 55684
rect 18417 55675 18475 55681
rect 18417 55672 18429 55675
rect 16448 55644 18429 55672
rect 16448 55632 16454 55644
rect 18417 55641 18429 55644
rect 18463 55672 18475 55675
rect 18598 55672 18604 55684
rect 18463 55644 18604 55672
rect 18463 55641 18475 55644
rect 18417 55635 18475 55641
rect 18598 55632 18604 55644
rect 18656 55632 18662 55684
rect 20456 55616 20484 55712
rect 20993 55709 21005 55712
rect 21039 55709 21051 55743
rect 27614 55740 27620 55752
rect 27575 55712 27620 55740
rect 20993 55703 21051 55709
rect 27614 55700 27620 55712
rect 27672 55740 27678 55752
rect 28261 55743 28319 55749
rect 28261 55740 28273 55743
rect 27672 55712 28273 55740
rect 27672 55700 27678 55712
rect 28261 55709 28273 55712
rect 28307 55709 28319 55743
rect 28261 55703 28319 55709
rect 39850 55672 39856 55684
rect 27816 55644 39856 55672
rect 14182 55604 14188 55616
rect 14143 55576 14188 55604
rect 14182 55564 14188 55576
rect 14240 55564 14246 55616
rect 15102 55604 15108 55616
rect 15063 55576 15108 55604
rect 15102 55564 15108 55576
rect 15160 55564 15166 55616
rect 16574 55564 16580 55616
rect 16632 55604 16638 55616
rect 17218 55604 17224 55616
rect 16632 55576 16677 55604
rect 17179 55576 17224 55604
rect 16632 55564 16638 55576
rect 17218 55564 17224 55576
rect 17276 55564 17282 55616
rect 19058 55564 19064 55616
rect 19116 55604 19122 55616
rect 19245 55607 19303 55613
rect 19245 55604 19257 55607
rect 19116 55576 19257 55604
rect 19116 55564 19122 55576
rect 19245 55573 19257 55576
rect 19291 55573 19303 55607
rect 20438 55604 20444 55616
rect 20399 55576 20444 55604
rect 19245 55567 19303 55573
rect 20438 55564 20444 55576
rect 20496 55564 20502 55616
rect 21910 55604 21916 55616
rect 21871 55576 21916 55604
rect 21910 55564 21916 55576
rect 21968 55564 21974 55616
rect 27816 55613 27844 55644
rect 39850 55632 39856 55644
rect 39908 55632 39914 55684
rect 27801 55607 27859 55613
rect 27801 55573 27813 55607
rect 27847 55573 27859 55607
rect 30006 55604 30012 55616
rect 29967 55576 30012 55604
rect 27801 55567 27859 55573
rect 30006 55564 30012 55576
rect 30064 55564 30070 55616
rect 42797 55607 42855 55613
rect 42797 55573 42809 55607
rect 42843 55604 42855 55607
rect 42886 55604 42892 55616
rect 42843 55576 42892 55604
rect 42843 55573 42855 55576
rect 42797 55567 42855 55573
rect 42886 55564 42892 55576
rect 42944 55564 42950 55616
rect 43441 55607 43499 55613
rect 43441 55573 43453 55607
rect 43487 55604 43499 55607
rect 43530 55604 43536 55616
rect 43487 55576 43536 55604
rect 43487 55573 43499 55576
rect 43441 55567 43499 55573
rect 43530 55564 43536 55576
rect 43588 55564 43594 55616
rect 43990 55604 43996 55616
rect 43951 55576 43996 55604
rect 43990 55564 43996 55576
rect 44048 55564 44054 55616
rect 44726 55564 44732 55616
rect 44784 55604 44790 55616
rect 45005 55607 45063 55613
rect 45005 55604 45017 55607
rect 44784 55576 45017 55604
rect 44784 55564 44790 55576
rect 45005 55573 45017 55576
rect 45051 55573 45063 55607
rect 45005 55567 45063 55573
rect 46017 55607 46075 55613
rect 46017 55573 46029 55607
rect 46063 55604 46075 55607
rect 46106 55604 46112 55616
rect 46063 55576 46112 55604
rect 46063 55573 46075 55576
rect 46017 55567 46075 55573
rect 46106 55564 46112 55576
rect 46164 55564 46170 55616
rect 46661 55607 46719 55613
rect 46661 55573 46673 55607
rect 46707 55604 46719 55607
rect 46750 55604 46756 55616
rect 46707 55576 46756 55604
rect 46707 55573 46719 55576
rect 46661 55567 46719 55573
rect 46750 55564 46756 55576
rect 46808 55564 46814 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 23934 55360 23940 55412
rect 23992 55400 23998 55412
rect 43990 55400 43996 55412
rect 23992 55372 43996 55400
rect 23992 55360 23998 55372
rect 43990 55360 43996 55372
rect 44048 55360 44054 55412
rect 58158 55128 58164 55140
rect 58119 55100 58164 55128
rect 58158 55088 58164 55100
rect 58216 55088 58222 55140
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 57882 53932 57888 53984
rect 57940 53972 57946 53984
rect 58161 53975 58219 53981
rect 58161 53972 58173 53975
rect 57940 53944 58173 53972
rect 57940 53932 57946 53944
rect 58161 53941 58173 53944
rect 58207 53941 58219 53975
rect 58161 53935 58219 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 57882 52436 57888 52488
rect 57940 52476 57946 52488
rect 58161 52479 58219 52485
rect 58161 52476 58173 52479
rect 57940 52448 58173 52476
rect 57940 52436 57946 52448
rect 58161 52445 58173 52448
rect 58207 52445 58219 52479
rect 58161 52439 58219 52445
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 43162 51388 43168 51400
rect 43123 51360 43168 51388
rect 43162 51348 43168 51360
rect 43220 51388 43226 51400
rect 43809 51391 43867 51397
rect 43809 51388 43821 51391
rect 43220 51360 43821 51388
rect 43220 51348 43226 51360
rect 43809 51357 43821 51360
rect 43855 51357 43867 51391
rect 58158 51388 58164 51400
rect 58119 51360 58164 51388
rect 43809 51351 43867 51357
rect 58158 51348 58164 51360
rect 58216 51348 58222 51400
rect 43364 51292 45554 51320
rect 43364 51261 43392 51292
rect 43349 51255 43407 51261
rect 43349 51221 43361 51255
rect 43395 51221 43407 51255
rect 45526 51252 45554 51292
rect 56042 51252 56048 51264
rect 45526 51224 56048 51252
rect 43349 51215 43407 51221
rect 56042 51212 56048 51224
rect 56100 51212 56106 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 58158 49756 58164 49768
rect 58119 49728 58164 49756
rect 58158 49716 58164 49728
rect 58216 49716 58222 49768
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 58158 48532 58164 48544
rect 58119 48504 58164 48532
rect 58158 48492 58164 48504
rect 58216 48492 58222 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58158 47036 58164 47048
rect 58119 47008 58164 47036
rect 58158 46996 58164 47008
rect 58216 46996 58222 47048
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 58158 45948 58164 45960
rect 58119 45920 58164 45948
rect 58158 45908 58164 45920
rect 58216 45908 58222 45960
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 56318 45472 56324 45484
rect 56279 45444 56324 45472
rect 56318 45432 56324 45444
rect 56376 45472 56382 45484
rect 56965 45475 57023 45481
rect 56965 45472 56977 45475
rect 56376 45444 56977 45472
rect 56376 45432 56382 45444
rect 56965 45441 56977 45444
rect 57011 45441 57023 45475
rect 56965 45435 57023 45441
rect 56505 45339 56563 45345
rect 56505 45305 56517 45339
rect 56551 45336 56563 45339
rect 57790 45336 57796 45348
rect 56551 45308 57796 45336
rect 56551 45305 56563 45308
rect 56505 45299 56563 45305
rect 57790 45296 57796 45308
rect 57848 45296 57854 45348
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 58158 44248 58164 44260
rect 58119 44220 58164 44248
rect 58158 44208 58164 44220
rect 58216 44208 58222 44260
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 58158 43092 58164 43104
rect 58119 43064 58164 43092
rect 58158 43052 58164 43064
rect 58216 43052 58222 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 16942 42712 16948 42764
rect 17000 42752 17006 42764
rect 20438 42752 20444 42764
rect 17000 42724 20444 42752
rect 17000 42712 17006 42724
rect 20438 42712 20444 42724
rect 20496 42712 20502 42764
rect 15841 42551 15899 42557
rect 15841 42517 15853 42551
rect 15887 42548 15899 42551
rect 17218 42548 17224 42560
rect 15887 42520 17224 42548
rect 15887 42517 15899 42520
rect 15841 42511 15899 42517
rect 17218 42508 17224 42520
rect 17276 42508 17282 42560
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 12253 42211 12311 42217
rect 12253 42177 12265 42211
rect 12299 42177 12311 42211
rect 12253 42171 12311 42177
rect 12437 42211 12495 42217
rect 12437 42177 12449 42211
rect 12483 42208 12495 42211
rect 12526 42208 12532 42220
rect 12483 42180 12532 42208
rect 12483 42177 12495 42180
rect 12437 42171 12495 42177
rect 12268 42140 12296 42171
rect 12526 42168 12532 42180
rect 12584 42168 12590 42220
rect 15010 42208 15016 42220
rect 14971 42180 15016 42208
rect 15010 42168 15016 42180
rect 15068 42168 15074 42220
rect 15194 42208 15200 42220
rect 15155 42180 15200 42208
rect 15194 42168 15200 42180
rect 15252 42168 15258 42220
rect 15289 42211 15347 42217
rect 15289 42177 15301 42211
rect 15335 42177 15347 42211
rect 15289 42171 15347 42177
rect 15427 42211 15485 42217
rect 15427 42177 15439 42211
rect 15473 42208 15485 42211
rect 17218 42208 17224 42220
rect 15473 42180 17224 42208
rect 15473 42177 15485 42180
rect 15427 42171 15485 42177
rect 12268 42112 12434 42140
rect 12406 42084 12434 42112
rect 12710 42100 12716 42152
rect 12768 42140 12774 42152
rect 15304 42140 15332 42171
rect 17218 42168 17224 42180
rect 17276 42168 17282 42220
rect 15562 42140 15568 42152
rect 12768 42112 15568 42140
rect 12768 42100 12774 42112
rect 15562 42100 15568 42112
rect 15620 42100 15626 42152
rect 12406 42044 12440 42084
rect 12434 42032 12440 42044
rect 12492 42032 12498 42084
rect 12621 42007 12679 42013
rect 12621 41973 12633 42007
rect 12667 42004 12679 42007
rect 12802 42004 12808 42016
rect 12667 41976 12808 42004
rect 12667 41973 12679 41976
rect 12621 41967 12679 41973
rect 12802 41964 12808 41976
rect 12860 41964 12866 42016
rect 15654 42004 15660 42016
rect 15615 41976 15660 42004
rect 15654 41964 15660 41976
rect 15712 41964 15718 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 15194 41760 15200 41812
rect 15252 41800 15258 41812
rect 16577 41803 16635 41809
rect 16577 41800 16589 41803
rect 15252 41772 16589 41800
rect 15252 41760 15258 41772
rect 16577 41769 16589 41772
rect 16623 41769 16635 41803
rect 16577 41763 16635 41769
rect 11514 41732 11520 41744
rect 11475 41704 11520 41732
rect 11514 41692 11520 41704
rect 11572 41692 11578 41744
rect 12710 41692 12716 41744
rect 12768 41692 12774 41744
rect 18693 41735 18751 41741
rect 15488 41704 17172 41732
rect 12725 41605 12753 41692
rect 12894 41664 12900 41676
rect 12820 41636 12900 41664
rect 12820 41605 12848 41636
rect 12894 41624 12900 41636
rect 12952 41624 12958 41676
rect 14645 41667 14703 41673
rect 14645 41633 14657 41667
rect 14691 41664 14703 41667
rect 14691 41636 15332 41664
rect 14691 41633 14703 41636
rect 14645 41627 14703 41633
rect 12621 41599 12679 41605
rect 12621 41593 12633 41599
rect 12544 41565 12633 41593
rect 12667 41565 12679 41599
rect 11698 41528 11704 41540
rect 11659 41500 11704 41528
rect 11698 41488 11704 41500
rect 11756 41488 11762 41540
rect 11885 41531 11943 41537
rect 11885 41497 11897 41531
rect 11931 41528 11943 41531
rect 12544 41528 12572 41565
rect 12621 41559 12679 41565
rect 12713 41599 12771 41605
rect 12713 41565 12725 41599
rect 12759 41565 12771 41599
rect 12713 41559 12771 41565
rect 12805 41599 12863 41605
rect 12805 41565 12817 41599
rect 12851 41565 12863 41599
rect 12986 41596 12992 41608
rect 12947 41568 12992 41596
rect 12805 41559 12863 41565
rect 12986 41556 12992 41568
rect 13044 41556 13050 41608
rect 14734 41556 14740 41608
rect 14792 41596 14798 41608
rect 15010 41596 15016 41608
rect 14792 41568 15016 41596
rect 14792 41556 14798 41568
rect 15010 41556 15016 41568
rect 15068 41596 15074 41608
rect 15304 41605 15332 41636
rect 15488 41605 15516 41704
rect 15749 41667 15807 41673
rect 15749 41633 15761 41667
rect 15795 41664 15807 41667
rect 16574 41664 16580 41676
rect 15795 41636 16580 41664
rect 15795 41633 15807 41636
rect 15749 41627 15807 41633
rect 16574 41624 16580 41636
rect 16632 41624 16638 41676
rect 15105 41599 15163 41605
rect 15105 41596 15117 41599
rect 15068 41568 15117 41596
rect 15068 41556 15074 41568
rect 15105 41565 15117 41568
rect 15151 41565 15163 41599
rect 15105 41559 15163 41565
rect 15289 41599 15347 41605
rect 15289 41565 15301 41599
rect 15335 41565 15347 41599
rect 15289 41559 15347 41565
rect 15381 41599 15439 41605
rect 15381 41565 15393 41599
rect 15427 41565 15439 41599
rect 15381 41559 15439 41565
rect 15473 41599 15531 41605
rect 15473 41565 15485 41599
rect 15519 41565 15531 41599
rect 15473 41559 15531 41565
rect 13541 41531 13599 41537
rect 13541 41528 13553 41531
rect 11931 41500 12480 41528
rect 12544 41500 13553 41528
rect 11931 41497 11943 41500
rect 11885 41491 11943 41497
rect 12452 41472 12480 41500
rect 13541 41497 13553 41500
rect 13587 41528 13599 41531
rect 13814 41528 13820 41540
rect 13587 41500 13820 41528
rect 13587 41497 13599 41500
rect 13541 41491 13599 41497
rect 13814 41488 13820 41500
rect 13872 41488 13878 41540
rect 14277 41531 14335 41537
rect 14277 41497 14289 41531
rect 14323 41497 14335 41531
rect 14277 41491 14335 41497
rect 14461 41531 14519 41537
rect 14461 41497 14473 41531
rect 14507 41528 14519 41531
rect 15194 41528 15200 41540
rect 14507 41500 15200 41528
rect 14507 41497 14519 41500
rect 14461 41491 14519 41497
rect 9674 41460 9680 41472
rect 9635 41432 9680 41460
rect 9674 41420 9680 41432
rect 9732 41420 9738 41472
rect 12342 41460 12348 41472
rect 12303 41432 12348 41460
rect 12342 41420 12348 41432
rect 12400 41420 12406 41472
rect 12434 41420 12440 41472
rect 12492 41460 12498 41472
rect 14292 41460 14320 41491
rect 15194 41488 15200 41500
rect 15252 41488 15258 41540
rect 15396 41528 15424 41559
rect 15562 41528 15568 41540
rect 15396 41500 15568 41528
rect 15562 41488 15568 41500
rect 15620 41488 15626 41540
rect 16209 41531 16267 41537
rect 16209 41528 16221 41531
rect 15672 41500 16221 41528
rect 14550 41460 14556 41472
rect 12492 41432 14556 41460
rect 12492 41420 12498 41432
rect 14550 41420 14556 41432
rect 14608 41460 14614 41472
rect 15672 41460 15700 41500
rect 16209 41497 16221 41500
rect 16255 41497 16267 41531
rect 16209 41491 16267 41497
rect 16393 41531 16451 41537
rect 16393 41497 16405 41531
rect 16439 41528 16451 41531
rect 16758 41528 16764 41540
rect 16439 41500 16764 41528
rect 16439 41497 16451 41500
rect 16393 41491 16451 41497
rect 16758 41488 16764 41500
rect 16816 41488 16822 41540
rect 17144 41537 17172 41704
rect 18693 41701 18705 41735
rect 18739 41732 18751 41735
rect 19886 41732 19892 41744
rect 18739 41704 19892 41732
rect 18739 41701 18751 41704
rect 18693 41695 18751 41701
rect 19886 41692 19892 41704
rect 19944 41692 19950 41744
rect 20346 41664 20352 41676
rect 19628 41636 20352 41664
rect 17218 41556 17224 41608
rect 17276 41596 17282 41608
rect 19628 41605 19656 41636
rect 20346 41624 20352 41636
rect 20404 41624 20410 41676
rect 19521 41599 19579 41605
rect 19521 41596 19533 41599
rect 17276 41568 19533 41596
rect 17276 41556 17282 41568
rect 19521 41565 19533 41568
rect 19567 41565 19579 41599
rect 19521 41559 19579 41565
rect 19613 41599 19671 41605
rect 19613 41565 19625 41599
rect 19659 41565 19671 41599
rect 19613 41559 19671 41565
rect 19705 41599 19763 41605
rect 19705 41565 19717 41599
rect 19751 41565 19763 41599
rect 19886 41596 19892 41608
rect 19847 41568 19892 41596
rect 19705 41559 19763 41565
rect 17129 41531 17187 41537
rect 17129 41497 17141 41531
rect 17175 41528 17187 41531
rect 19334 41528 19340 41540
rect 17175 41500 19340 41528
rect 17175 41497 17187 41500
rect 17129 41491 17187 41497
rect 19334 41488 19340 41500
rect 19392 41488 19398 41540
rect 19536 41528 19564 41559
rect 19720 41528 19748 41559
rect 19886 41556 19892 41568
rect 19944 41556 19950 41608
rect 58158 41596 58164 41608
rect 58119 41568 58164 41596
rect 58158 41556 58164 41568
rect 58216 41556 58222 41608
rect 20162 41528 20168 41540
rect 19536 41500 19656 41528
rect 19720 41500 20168 41528
rect 14608 41432 15700 41460
rect 19245 41463 19303 41469
rect 14608 41420 14614 41432
rect 19245 41429 19257 41463
rect 19291 41460 19303 41463
rect 19426 41460 19432 41472
rect 19291 41432 19432 41460
rect 19291 41429 19303 41432
rect 19245 41423 19303 41429
rect 19426 41420 19432 41432
rect 19484 41420 19490 41472
rect 19628 41460 19656 41500
rect 20162 41488 20168 41500
rect 20220 41488 20226 41540
rect 20441 41463 20499 41469
rect 20441 41460 20453 41463
rect 19628 41432 20453 41460
rect 20441 41429 20453 41432
rect 20487 41460 20499 41463
rect 24394 41460 24400 41472
rect 20487 41432 24400 41460
rect 20487 41429 20499 41432
rect 20441 41423 20499 41429
rect 24394 41420 24400 41432
rect 24452 41420 24458 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 9950 41216 9956 41268
rect 10008 41256 10014 41268
rect 10965 41259 11023 41265
rect 10965 41256 10977 41259
rect 10008 41228 10977 41256
rect 10008 41216 10014 41228
rect 10965 41225 10977 41228
rect 11011 41256 11023 41259
rect 18506 41256 18512 41268
rect 11011 41228 18512 41256
rect 11011 41225 11023 41228
rect 10965 41219 11023 41225
rect 18506 41216 18512 41228
rect 18564 41256 18570 41268
rect 23014 41256 23020 41268
rect 18564 41228 23020 41256
rect 18564 41216 18570 41228
rect 23014 41216 23020 41228
rect 23072 41216 23078 41268
rect 9858 41188 9864 41200
rect 9324 41160 9864 41188
rect 9324 41129 9352 41160
rect 9858 41148 9864 41160
rect 9916 41148 9922 41200
rect 14642 41148 14648 41200
rect 14700 41188 14706 41200
rect 15933 41191 15991 41197
rect 14700 41160 14872 41188
rect 14700 41148 14706 41160
rect 9217 41123 9275 41129
rect 9217 41089 9229 41123
rect 9263 41089 9275 41123
rect 9217 41083 9275 41089
rect 9309 41123 9367 41129
rect 9309 41089 9321 41123
rect 9355 41089 9367 41123
rect 9309 41083 9367 41089
rect 9232 41052 9260 41083
rect 9398 41080 9404 41132
rect 9456 41120 9462 41132
rect 9585 41123 9643 41129
rect 9456 41092 9501 41120
rect 9456 41080 9462 41092
rect 9585 41089 9597 41123
rect 9631 41120 9643 41123
rect 10229 41123 10287 41129
rect 9631 41092 9812 41120
rect 9631 41089 9643 41092
rect 9585 41083 9643 41089
rect 9674 41052 9680 41064
rect 9232 41024 9680 41052
rect 9674 41012 9680 41024
rect 9732 41012 9738 41064
rect 9784 40984 9812 41092
rect 10229 41089 10241 41123
rect 10275 41120 10287 41123
rect 10318 41120 10324 41132
rect 10275 41092 10324 41120
rect 10275 41089 10287 41092
rect 10229 41083 10287 41089
rect 10318 41080 10324 41092
rect 10376 41080 10382 41132
rect 10413 41123 10471 41129
rect 10413 41089 10425 41123
rect 10459 41120 10471 41123
rect 10870 41120 10876 41132
rect 10459 41092 10876 41120
rect 10459 41089 10471 41092
rect 10413 41083 10471 41089
rect 10870 41080 10876 41092
rect 10928 41080 10934 41132
rect 12601 41123 12659 41129
rect 12452 41120 12572 41123
rect 12601 41120 12613 41123
rect 12452 41095 12613 41120
rect 10410 40984 10416 40996
rect 9784 40956 10416 40984
rect 10410 40944 10416 40956
rect 10468 40944 10474 40996
rect 12452 40984 12480 41095
rect 12544 41092 12613 41095
rect 12601 41089 12613 41092
rect 12647 41089 12659 41123
rect 12601 41083 12659 41089
rect 12713 41123 12771 41129
rect 12713 41089 12725 41123
rect 12759 41089 12771 41123
rect 12713 41083 12771 41089
rect 12728 41052 12756 41083
rect 12802 41080 12808 41132
rect 12860 41129 12866 41132
rect 12860 41120 12868 41129
rect 12860 41092 12905 41120
rect 12860 41083 12868 41092
rect 12860 41080 12866 41083
rect 12986 41080 12992 41132
rect 13044 41120 13050 41132
rect 14734 41120 14740 41132
rect 13044 41092 14740 41120
rect 13044 41080 13050 41092
rect 14734 41080 14740 41092
rect 14792 41080 14798 41132
rect 14844 41120 14872 41160
rect 15933 41157 15945 41191
rect 15979 41188 15991 41191
rect 17770 41188 17776 41200
rect 15979 41160 17776 41188
rect 15979 41157 15991 41160
rect 15933 41151 15991 41157
rect 14900 41123 14958 41129
rect 14900 41120 14912 41123
rect 14844 41092 14912 41120
rect 14900 41089 14912 41092
rect 14946 41089 14958 41123
rect 14900 41083 14958 41089
rect 15013 41123 15071 41129
rect 15013 41089 15025 41123
rect 15059 41089 15071 41123
rect 15013 41083 15071 41089
rect 15151 41123 15209 41129
rect 15151 41089 15163 41123
rect 15197 41120 15209 41123
rect 15948 41120 15976 41151
rect 17770 41148 17776 41160
rect 17828 41148 17834 41200
rect 19426 41148 19432 41200
rect 19484 41197 19490 41200
rect 19484 41188 19496 41197
rect 24762 41188 24768 41200
rect 19484 41160 19529 41188
rect 19628 41160 24768 41188
rect 19484 41151 19496 41160
rect 19484 41148 19490 41151
rect 19628 41120 19656 41160
rect 24762 41148 24768 41160
rect 24820 41148 24826 41200
rect 15197 41092 15976 41120
rect 16546 41092 19656 41120
rect 15197 41089 15209 41092
rect 15151 41083 15209 41089
rect 12894 41052 12900 41064
rect 12728 41024 12900 41052
rect 12894 41012 12900 41024
rect 12952 41012 12958 41064
rect 15028 41052 15056 41083
rect 15562 41052 15568 41064
rect 15028 41024 15568 41052
rect 15562 41012 15568 41024
rect 15620 41012 15626 41064
rect 13541 40987 13599 40993
rect 13541 40984 13553 40987
rect 12452 40956 13553 40984
rect 13541 40953 13553 40956
rect 13587 40984 13599 40987
rect 14734 40984 14740 40996
rect 13587 40956 14740 40984
rect 13587 40953 13599 40956
rect 13541 40947 13599 40953
rect 14734 40944 14740 40956
rect 14792 40944 14798 40996
rect 15010 40944 15016 40996
rect 15068 40984 15074 40996
rect 16546 40984 16574 41092
rect 20070 41080 20076 41132
rect 20128 41120 20134 41132
rect 20349 41123 20407 41129
rect 20349 41120 20361 41123
rect 20128 41092 20361 41120
rect 20128 41080 20134 41092
rect 20349 41089 20361 41092
rect 20395 41089 20407 41123
rect 20349 41083 20407 41089
rect 20533 41123 20591 41129
rect 20533 41089 20545 41123
rect 20579 41120 20591 41123
rect 20714 41120 20720 41132
rect 20579 41092 20720 41120
rect 20579 41089 20591 41092
rect 20533 41083 20591 41089
rect 20714 41080 20720 41092
rect 20772 41080 20778 41132
rect 22094 41080 22100 41132
rect 22152 41120 22158 41132
rect 22557 41123 22615 41129
rect 22557 41120 22569 41123
rect 22152 41092 22569 41120
rect 22152 41080 22158 41092
rect 22557 41089 22569 41092
rect 22603 41089 22615 41123
rect 22557 41083 22615 41089
rect 22741 41123 22799 41129
rect 22741 41089 22753 41123
rect 22787 41120 22799 41123
rect 23382 41120 23388 41132
rect 22787 41092 23388 41120
rect 22787 41089 22799 41092
rect 22741 41083 22799 41089
rect 23382 41080 23388 41092
rect 23440 41080 23446 41132
rect 19705 41055 19763 41061
rect 19705 41021 19717 41055
rect 19751 41021 19763 41055
rect 19705 41015 19763 41021
rect 15068 40956 16574 40984
rect 19720 40984 19748 41015
rect 20622 40984 20628 40996
rect 19720 40956 20628 40984
rect 15068 40944 15074 40956
rect 8938 40916 8944 40928
rect 8899 40888 8944 40916
rect 8938 40876 8944 40888
rect 8996 40876 9002 40928
rect 10045 40919 10103 40925
rect 10045 40885 10057 40919
rect 10091 40916 10103 40919
rect 10134 40916 10140 40928
rect 10091 40888 10140 40916
rect 10091 40885 10103 40888
rect 10045 40879 10103 40885
rect 10134 40876 10140 40888
rect 10192 40876 10198 40928
rect 11790 40876 11796 40928
rect 11848 40916 11854 40928
rect 12345 40919 12403 40925
rect 12345 40916 12357 40919
rect 11848 40888 12357 40916
rect 11848 40876 11854 40888
rect 12345 40885 12357 40888
rect 12391 40885 12403 40919
rect 15378 40916 15384 40928
rect 15339 40888 15384 40916
rect 12345 40879 12403 40885
rect 15378 40876 15384 40888
rect 15436 40876 15442 40928
rect 17954 40876 17960 40928
rect 18012 40916 18018 40928
rect 18325 40919 18383 40925
rect 18325 40916 18337 40919
rect 18012 40888 18337 40916
rect 18012 40876 18018 40888
rect 18325 40885 18337 40888
rect 18371 40885 18383 40919
rect 18325 40879 18383 40885
rect 19334 40876 19340 40928
rect 19392 40916 19398 40928
rect 19720 40916 19748 40956
rect 20622 40944 20628 40956
rect 20680 40944 20686 40996
rect 19392 40888 19748 40916
rect 19392 40876 19398 40888
rect 19794 40876 19800 40928
rect 19852 40916 19858 40928
rect 20165 40919 20223 40925
rect 20165 40916 20177 40919
rect 19852 40888 20177 40916
rect 19852 40876 19858 40888
rect 20165 40885 20177 40888
rect 20211 40885 20223 40919
rect 20165 40879 20223 40885
rect 22646 40876 22652 40928
rect 22704 40916 22710 40928
rect 22925 40919 22983 40925
rect 22925 40916 22937 40919
rect 22704 40888 22937 40916
rect 22704 40876 22710 40888
rect 22925 40885 22937 40888
rect 22971 40885 22983 40919
rect 22925 40879 22983 40885
rect 23014 40876 23020 40928
rect 23072 40916 23078 40928
rect 23477 40919 23535 40925
rect 23477 40916 23489 40919
rect 23072 40888 23489 40916
rect 23072 40876 23078 40888
rect 23477 40885 23489 40888
rect 23523 40916 23535 40919
rect 26602 40916 26608 40928
rect 23523 40888 26608 40916
rect 23523 40885 23535 40888
rect 23477 40879 23535 40885
rect 26602 40876 26608 40888
rect 26660 40876 26666 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 14642 40672 14648 40724
rect 14700 40712 14706 40724
rect 14921 40715 14979 40721
rect 14921 40712 14933 40715
rect 14700 40684 14933 40712
rect 14700 40672 14706 40684
rect 14921 40681 14933 40684
rect 14967 40681 14979 40715
rect 14921 40675 14979 40681
rect 18693 40715 18751 40721
rect 18693 40681 18705 40715
rect 18739 40712 18751 40715
rect 20162 40712 20168 40724
rect 18739 40684 20168 40712
rect 18739 40681 18751 40684
rect 18693 40675 18751 40681
rect 20162 40672 20168 40684
rect 20220 40672 20226 40724
rect 4890 40644 4896 40656
rect 3988 40616 4896 40644
rect 3988 40505 4016 40616
rect 4890 40604 4896 40616
rect 4948 40604 4954 40656
rect 9674 40604 9680 40656
rect 9732 40644 9738 40656
rect 14274 40644 14280 40656
rect 9732 40616 14280 40644
rect 9732 40604 9738 40616
rect 14274 40604 14280 40616
rect 14332 40604 14338 40656
rect 17865 40647 17923 40653
rect 17865 40613 17877 40647
rect 17911 40644 17923 40647
rect 19518 40644 19524 40656
rect 17911 40616 19524 40644
rect 17911 40613 17923 40616
rect 17865 40607 17923 40613
rect 19518 40604 19524 40616
rect 19576 40604 19582 40656
rect 19978 40644 19984 40656
rect 19628 40616 19984 40644
rect 12986 40536 12992 40588
rect 13044 40576 13050 40588
rect 13173 40579 13231 40585
rect 13173 40576 13185 40579
rect 13044 40548 13185 40576
rect 13044 40536 13050 40548
rect 13173 40545 13185 40548
rect 13219 40545 13231 40579
rect 13173 40539 13231 40545
rect 4045 40511 4103 40517
rect 4045 40505 4057 40511
rect 3988 40477 4057 40505
rect 4091 40477 4103 40511
rect 4045 40471 4103 40477
rect 4154 40505 4212 40511
rect 4154 40471 4166 40505
rect 4200 40471 4212 40505
rect 4154 40465 4212 40471
rect 4246 40468 4252 40520
rect 4304 40517 4310 40520
rect 4304 40508 4312 40517
rect 4433 40511 4491 40517
rect 4304 40480 4349 40508
rect 4304 40471 4312 40480
rect 4433 40477 4445 40511
rect 4479 40508 4491 40511
rect 4798 40508 4804 40520
rect 4479 40480 4804 40508
rect 4479 40477 4491 40480
rect 4433 40471 4491 40477
rect 4304 40468 4310 40471
rect 4798 40468 4804 40480
rect 4856 40468 4862 40520
rect 6086 40508 6092 40520
rect 6047 40480 6092 40508
rect 6086 40468 6092 40480
rect 6144 40468 6150 40520
rect 9950 40508 9956 40520
rect 9911 40480 9956 40508
rect 9950 40468 9956 40480
rect 10008 40468 10014 40520
rect 10045 40511 10103 40517
rect 10045 40477 10057 40511
rect 10091 40477 10103 40511
rect 10045 40471 10103 40477
rect 3786 40372 3792 40384
rect 3747 40344 3792 40372
rect 3786 40332 3792 40344
rect 3844 40332 3850 40384
rect 4172 40372 4200 40465
rect 4890 40440 4896 40452
rect 4851 40412 4896 40440
rect 4890 40400 4896 40412
rect 4948 40400 4954 40452
rect 5810 40400 5816 40452
rect 5868 40440 5874 40452
rect 6334 40443 6392 40449
rect 6334 40440 6346 40443
rect 5868 40412 6346 40440
rect 5868 40400 5874 40412
rect 6334 40409 6346 40412
rect 6380 40409 6392 40443
rect 7190 40440 7196 40452
rect 6334 40403 6392 40409
rect 6472 40412 7196 40440
rect 5442 40372 5448 40384
rect 4172 40344 5448 40372
rect 5442 40332 5448 40344
rect 5500 40332 5506 40384
rect 5629 40375 5687 40381
rect 5629 40341 5641 40375
rect 5675 40372 5687 40375
rect 5718 40372 5724 40384
rect 5675 40344 5724 40372
rect 5675 40341 5687 40344
rect 5629 40335 5687 40341
rect 5718 40332 5724 40344
rect 5776 40372 5782 40384
rect 6472 40372 6500 40412
rect 7190 40400 7196 40412
rect 7248 40400 7254 40452
rect 9858 40400 9864 40452
rect 9916 40440 9922 40452
rect 10060 40440 10088 40471
rect 10134 40468 10140 40520
rect 10192 40508 10198 40520
rect 10321 40511 10379 40517
rect 10192 40480 10237 40508
rect 10192 40468 10198 40480
rect 10321 40477 10333 40511
rect 10367 40508 10379 40511
rect 10410 40508 10416 40520
rect 10367 40480 10416 40508
rect 10367 40477 10379 40480
rect 10321 40471 10379 40477
rect 10410 40468 10416 40480
rect 10468 40468 10474 40520
rect 10870 40468 10876 40520
rect 10928 40508 10934 40520
rect 11149 40511 11207 40517
rect 11149 40508 11161 40511
rect 10928 40480 11161 40508
rect 10928 40468 10934 40480
rect 11149 40477 11161 40480
rect 11195 40477 11207 40511
rect 13449 40511 13507 40517
rect 13449 40508 13461 40511
rect 11149 40471 11207 40477
rect 13188 40480 13461 40508
rect 13188 40452 13216 40480
rect 13449 40477 13461 40480
rect 13495 40477 13507 40511
rect 13449 40471 13507 40477
rect 14458 40468 14464 40520
rect 14516 40508 14522 40520
rect 14553 40511 14611 40517
rect 14553 40508 14565 40511
rect 14516 40480 14565 40508
rect 14516 40468 14522 40480
rect 14553 40477 14565 40480
rect 14599 40477 14611 40511
rect 14553 40471 14611 40477
rect 15381 40511 15439 40517
rect 15381 40477 15393 40511
rect 15427 40508 15439 40511
rect 16114 40508 16120 40520
rect 15427 40480 16120 40508
rect 15427 40477 15439 40480
rect 15381 40471 15439 40477
rect 16114 40468 16120 40480
rect 16172 40468 16178 40520
rect 17954 40468 17960 40520
rect 18012 40508 18018 40520
rect 18509 40511 18567 40517
rect 18509 40508 18521 40511
rect 18012 40480 18521 40508
rect 18012 40468 18018 40480
rect 18509 40477 18521 40480
rect 18555 40477 18567 40511
rect 18509 40471 18567 40477
rect 19426 40468 19432 40520
rect 19484 40508 19490 40520
rect 19628 40517 19656 40616
rect 19978 40604 19984 40616
rect 20036 40644 20042 40656
rect 20346 40644 20352 40656
rect 20036 40616 20352 40644
rect 20036 40604 20042 40616
rect 20346 40604 20352 40616
rect 20404 40604 20410 40656
rect 20622 40536 20628 40588
rect 20680 40576 20686 40588
rect 20717 40579 20775 40585
rect 20717 40576 20729 40579
rect 20680 40548 20729 40576
rect 20680 40536 20686 40548
rect 20717 40545 20729 40548
rect 20763 40545 20775 40579
rect 20717 40539 20775 40545
rect 19521 40511 19579 40517
rect 19521 40508 19533 40511
rect 19484 40480 19533 40508
rect 19484 40468 19490 40480
rect 19521 40477 19533 40480
rect 19567 40477 19579 40511
rect 19521 40471 19579 40477
rect 19613 40511 19671 40517
rect 19613 40477 19625 40511
rect 19659 40477 19671 40511
rect 19613 40471 19671 40477
rect 19705 40511 19763 40517
rect 19705 40477 19717 40511
rect 19751 40508 19763 40511
rect 19794 40508 19800 40520
rect 19751 40480 19800 40508
rect 19751 40477 19763 40480
rect 19705 40471 19763 40477
rect 9916 40412 10088 40440
rect 9916 40400 9922 40412
rect 10502 40400 10508 40452
rect 10560 40440 10566 40452
rect 10965 40443 11023 40449
rect 10965 40440 10977 40443
rect 10560 40412 10977 40440
rect 10560 40400 10566 40412
rect 10965 40409 10977 40412
rect 11011 40409 11023 40443
rect 13170 40440 13176 40452
rect 10965 40403 11023 40409
rect 12406 40412 13176 40440
rect 5776 40344 6500 40372
rect 5776 40332 5782 40344
rect 6914 40332 6920 40384
rect 6972 40372 6978 40384
rect 7469 40375 7527 40381
rect 7469 40372 7481 40375
rect 6972 40344 7481 40372
rect 6972 40332 6978 40344
rect 7469 40341 7481 40344
rect 7515 40372 7527 40375
rect 8110 40372 8116 40384
rect 7515 40344 8116 40372
rect 7515 40341 7527 40344
rect 7469 40335 7527 40341
rect 8110 40332 8116 40344
rect 8168 40332 8174 40384
rect 9674 40372 9680 40384
rect 9635 40344 9680 40372
rect 9674 40332 9680 40344
rect 9732 40332 9738 40384
rect 10778 40372 10784 40384
rect 10739 40344 10784 40372
rect 10778 40332 10784 40344
rect 10836 40332 10842 40384
rect 11054 40332 11060 40384
rect 11112 40372 11118 40384
rect 12069 40375 12127 40381
rect 12069 40372 12081 40375
rect 11112 40344 12081 40372
rect 11112 40332 11118 40344
rect 12069 40341 12081 40344
rect 12115 40372 12127 40375
rect 12406 40372 12434 40412
rect 13170 40400 13176 40412
rect 13228 40400 13234 40452
rect 14734 40440 14740 40452
rect 14695 40412 14740 40440
rect 14734 40400 14740 40412
rect 14792 40400 14798 40452
rect 15654 40449 15660 40452
rect 15648 40403 15660 40449
rect 15712 40440 15718 40452
rect 18325 40443 18383 40449
rect 15712 40412 15748 40440
rect 15654 40400 15660 40403
rect 15712 40400 15718 40412
rect 18325 40409 18337 40443
rect 18371 40440 18383 40443
rect 19536 40440 19564 40471
rect 19794 40468 19800 40480
rect 19852 40468 19858 40520
rect 19886 40468 19892 40520
rect 19944 40508 19950 40520
rect 20438 40508 20444 40520
rect 19944 40480 20444 40508
rect 19944 40468 19950 40480
rect 20438 40468 20444 40480
rect 20496 40468 20502 40520
rect 22278 40468 22284 40520
rect 22336 40508 22342 40520
rect 22557 40511 22615 40517
rect 22557 40508 22569 40511
rect 22336 40480 22569 40508
rect 22336 40468 22342 40480
rect 22557 40477 22569 40480
rect 22603 40477 22615 40511
rect 22738 40508 22744 40520
rect 22699 40480 22744 40508
rect 22557 40471 22615 40477
rect 22738 40468 22744 40480
rect 22796 40468 22802 40520
rect 22833 40511 22891 40517
rect 22833 40477 22845 40511
rect 22879 40477 22891 40511
rect 22833 40471 22891 40477
rect 22925 40511 22983 40517
rect 22925 40477 22937 40511
rect 22971 40508 22983 40511
rect 23014 40508 23020 40520
rect 22971 40480 23020 40508
rect 22971 40477 22983 40480
rect 22925 40471 22983 40477
rect 20346 40440 20352 40452
rect 18371 40412 19472 40440
rect 19536 40412 20352 40440
rect 18371 40409 18383 40412
rect 18325 40403 18383 40409
rect 16758 40372 16764 40384
rect 12115 40344 12434 40372
rect 16719 40344 16764 40372
rect 12115 40341 12127 40344
rect 12069 40335 12127 40341
rect 16758 40332 16764 40344
rect 16816 40332 16822 40384
rect 19242 40372 19248 40384
rect 19203 40344 19248 40372
rect 19242 40332 19248 40344
rect 19300 40332 19306 40384
rect 19444 40372 19472 40412
rect 20346 40400 20352 40412
rect 20404 40400 20410 40452
rect 20984 40443 21042 40449
rect 20984 40409 20996 40443
rect 21030 40440 21042 40443
rect 21358 40440 21364 40452
rect 21030 40412 21364 40440
rect 21030 40409 21042 40412
rect 20984 40403 21042 40409
rect 21358 40400 21364 40412
rect 21416 40400 21422 40452
rect 21910 40400 21916 40452
rect 21968 40440 21974 40452
rect 22848 40440 22876 40471
rect 23014 40468 23020 40480
rect 23072 40468 23078 40520
rect 27246 40508 27252 40520
rect 27207 40480 27252 40508
rect 27246 40468 27252 40480
rect 27304 40468 27310 40520
rect 58158 40508 58164 40520
rect 58119 40480 58164 40508
rect 58158 40468 58164 40480
rect 58216 40468 58222 40520
rect 21968 40412 22876 40440
rect 21968 40400 21974 40412
rect 27154 40400 27160 40452
rect 27212 40440 27218 40452
rect 27494 40443 27552 40449
rect 27494 40440 27506 40443
rect 27212 40412 27506 40440
rect 27212 40400 27218 40412
rect 27494 40409 27506 40412
rect 27540 40409 27552 40443
rect 27494 40403 27552 40409
rect 20714 40372 20720 40384
rect 19444 40344 20720 40372
rect 20714 40332 20720 40344
rect 20772 40332 20778 40384
rect 22097 40375 22155 40381
rect 22097 40341 22109 40375
rect 22143 40372 22155 40375
rect 22554 40372 22560 40384
rect 22143 40344 22560 40372
rect 22143 40341 22155 40344
rect 22097 40335 22155 40341
rect 22554 40332 22560 40344
rect 22612 40332 22618 40384
rect 23201 40375 23259 40381
rect 23201 40341 23213 40375
rect 23247 40372 23259 40375
rect 23474 40372 23480 40384
rect 23247 40344 23480 40372
rect 23247 40341 23259 40344
rect 23201 40335 23259 40341
rect 23474 40332 23480 40344
rect 23532 40332 23538 40384
rect 23658 40372 23664 40384
rect 23619 40344 23664 40372
rect 23658 40332 23664 40344
rect 23716 40332 23722 40384
rect 28166 40332 28172 40384
rect 28224 40372 28230 40384
rect 28629 40375 28687 40381
rect 28629 40372 28641 40375
rect 28224 40344 28641 40372
rect 28224 40332 28230 40344
rect 28629 40341 28641 40344
rect 28675 40341 28687 40375
rect 28629 40335 28687 40341
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 3881 40171 3939 40177
rect 3881 40137 3893 40171
rect 3927 40137 3939 40171
rect 3881 40131 3939 40137
rect 2768 40103 2826 40109
rect 2768 40069 2780 40103
rect 2814 40100 2826 40103
rect 3786 40100 3792 40112
rect 2814 40072 3792 40100
rect 2814 40069 2826 40072
rect 2768 40063 2826 40069
rect 3786 40060 3792 40072
rect 3844 40060 3850 40112
rect 3896 40100 3924 40131
rect 4246 40128 4252 40180
rect 4304 40168 4310 40180
rect 4341 40171 4399 40177
rect 4341 40168 4353 40171
rect 4304 40140 4353 40168
rect 4304 40128 4310 40140
rect 4341 40137 4353 40140
rect 4387 40137 4399 40171
rect 5810 40168 5816 40180
rect 4341 40131 4399 40137
rect 5368 40140 5580 40168
rect 5771 40140 5816 40168
rect 4525 40103 4583 40109
rect 4525 40100 4537 40103
rect 3896 40072 4537 40100
rect 4525 40069 4537 40072
rect 4571 40100 4583 40103
rect 4982 40100 4988 40112
rect 4571 40072 4988 40100
rect 4571 40069 4583 40072
rect 4525 40063 4583 40069
rect 4982 40060 4988 40072
rect 5040 40060 5046 40112
rect 5368 40047 5396 40140
rect 5552 40100 5580 40140
rect 5810 40128 5816 40140
rect 5868 40128 5874 40180
rect 12526 40128 12532 40180
rect 12584 40168 12590 40180
rect 12894 40168 12900 40180
rect 12584 40140 12900 40168
rect 12584 40128 12590 40140
rect 12894 40128 12900 40140
rect 12952 40128 12958 40180
rect 13538 40128 13544 40180
rect 13596 40168 13602 40180
rect 14734 40168 14740 40180
rect 13596 40140 14740 40168
rect 13596 40128 13602 40140
rect 14734 40128 14740 40140
rect 14792 40128 14798 40180
rect 19242 40128 19248 40180
rect 19300 40168 19306 40180
rect 19518 40168 19524 40180
rect 19300 40140 19524 40168
rect 19300 40128 19306 40140
rect 19518 40128 19524 40140
rect 19576 40128 19582 40180
rect 22094 40168 22100 40180
rect 20916 40140 22100 40168
rect 6365 40103 6423 40109
rect 6365 40100 6377 40103
rect 5552 40072 6377 40100
rect 6365 40069 6377 40072
rect 6411 40069 6423 40103
rect 6365 40063 6423 40069
rect 6549 40103 6607 40109
rect 6549 40069 6561 40103
rect 6595 40100 6607 40103
rect 6914 40100 6920 40112
rect 6595 40072 6920 40100
rect 6595 40069 6607 40072
rect 6549 40063 6607 40069
rect 6914 40060 6920 40072
rect 6972 40060 6978 40112
rect 9858 40060 9864 40112
rect 9916 40100 9922 40112
rect 10778 40100 10784 40112
rect 9916 40072 10180 40100
rect 9916 40060 9922 40072
rect 4706 40032 4712 40044
rect 4667 40004 4712 40032
rect 4706 39992 4712 40004
rect 4764 39992 4770 40044
rect 4798 39992 4804 40044
rect 4856 40032 4862 40044
rect 5332 40041 5396 40047
rect 5193 40038 5251 40041
rect 5092 40035 5251 40038
rect 5092 40032 5205 40035
rect 4856 40010 5205 40032
rect 4856 40004 5120 40010
rect 5184 40004 5205 40010
rect 4856 39992 4862 40004
rect 5193 40001 5205 40004
rect 5239 40001 5251 40035
rect 5332 40007 5344 40041
rect 5378 40010 5396 40041
rect 5378 40007 5390 40010
rect 5332 40001 5390 40007
rect 5193 39995 5251 40001
rect 5442 39992 5448 40044
rect 5500 40032 5506 40044
rect 5583 40035 5641 40041
rect 5500 40004 5545 40032
rect 5500 39992 5506 40004
rect 5583 40001 5595 40035
rect 5629 40032 5641 40035
rect 5718 40032 5724 40044
rect 5629 40004 5724 40032
rect 5629 40001 5641 40004
rect 5583 39995 5641 40001
rect 5718 39992 5724 40004
rect 5776 39992 5782 40044
rect 6730 40032 6736 40044
rect 6691 40004 6736 40032
rect 6730 39992 6736 40004
rect 6788 39992 6794 40044
rect 7460 40035 7518 40041
rect 7460 40001 7472 40035
rect 7506 40032 7518 40035
rect 8938 40032 8944 40044
rect 7506 40004 8944 40032
rect 7506 40001 7518 40004
rect 7460 39995 7518 40001
rect 8938 39992 8944 40004
rect 8996 39992 9002 40044
rect 10152 40041 10180 40072
rect 10244 40072 10784 40100
rect 10244 40041 10272 40072
rect 10778 40060 10784 40072
rect 10836 40060 10842 40112
rect 11790 40109 11796 40112
rect 11784 40100 11796 40109
rect 11751 40072 11796 40100
rect 11784 40063 11796 40072
rect 11790 40060 11796 40063
rect 11848 40060 11854 40112
rect 15378 40060 15384 40112
rect 15436 40100 15442 40112
rect 15850 40103 15908 40109
rect 15850 40100 15862 40103
rect 15436 40072 15862 40100
rect 15436 40060 15442 40072
rect 15850 40069 15862 40072
rect 15896 40069 15908 40103
rect 15850 40063 15908 40069
rect 17402 40060 17408 40112
rect 17460 40100 17466 40112
rect 20916 40109 20944 40140
rect 22094 40128 22100 40140
rect 22152 40128 22158 40180
rect 22186 40128 22192 40180
rect 22244 40168 22250 40180
rect 23658 40168 23664 40180
rect 22244 40140 23664 40168
rect 22244 40128 22250 40140
rect 17957 40103 18015 40109
rect 17957 40100 17969 40103
rect 17460 40072 17969 40100
rect 17460 40060 17466 40072
rect 17957 40069 17969 40072
rect 18003 40069 18015 40103
rect 17957 40063 18015 40069
rect 20901 40103 20959 40109
rect 20901 40069 20913 40103
rect 20947 40069 20959 40103
rect 20901 40063 20959 40069
rect 21085 40103 21143 40109
rect 21085 40069 21097 40103
rect 21131 40100 21143 40103
rect 22554 40100 22560 40112
rect 21131 40072 22094 40100
rect 21131 40069 21143 40072
rect 21085 40063 21143 40069
rect 10045 40035 10103 40041
rect 10045 40001 10057 40035
rect 10091 40001 10103 40035
rect 10045 39995 10103 40001
rect 10137 40035 10195 40041
rect 10137 40001 10149 40035
rect 10183 40001 10195 40035
rect 10137 39995 10195 40001
rect 10229 40035 10287 40041
rect 10229 40001 10241 40035
rect 10275 40001 10287 40035
rect 10410 40032 10416 40044
rect 10371 40004 10416 40032
rect 10229 39995 10287 40001
rect 1854 39924 1860 39976
rect 1912 39964 1918 39976
rect 2501 39967 2559 39973
rect 2501 39964 2513 39967
rect 1912 39936 2513 39964
rect 1912 39924 1918 39936
rect 2501 39933 2513 39936
rect 2547 39933 2559 39967
rect 2501 39927 2559 39933
rect 6086 39924 6092 39976
rect 6144 39964 6150 39976
rect 7193 39967 7251 39973
rect 7193 39964 7205 39967
rect 6144 39936 7205 39964
rect 6144 39924 6150 39936
rect 7193 39933 7205 39936
rect 7239 39933 7251 39967
rect 10060 39964 10088 39995
rect 10410 39992 10416 40004
rect 10468 39992 10474 40044
rect 16114 40032 16120 40044
rect 16075 40004 16120 40032
rect 16114 39992 16120 40004
rect 16172 39992 16178 40044
rect 22066 40032 22094 40072
rect 22204 40072 22560 40100
rect 22204 40032 22232 40072
rect 22554 40060 22560 40072
rect 22612 40060 22618 40112
rect 22066 40004 22232 40032
rect 22278 39992 22284 40044
rect 22336 40032 22342 40044
rect 22465 40035 22523 40041
rect 22465 40032 22477 40035
rect 22336 40004 22477 40032
rect 22336 39992 22342 40004
rect 22465 40001 22477 40004
rect 22511 40001 22523 40035
rect 22646 40032 22652 40044
rect 22607 40004 22652 40032
rect 22465 39995 22523 40001
rect 22646 39992 22652 40004
rect 22704 39992 22710 40044
rect 22848 40041 22876 40140
rect 23658 40128 23664 40140
rect 23716 40128 23722 40180
rect 30834 40128 30840 40180
rect 30892 40168 30898 40180
rect 30892 40140 30972 40168
rect 30892 40128 30898 40140
rect 28166 40100 28172 40112
rect 28127 40072 28172 40100
rect 28166 40060 28172 40072
rect 28224 40060 28230 40112
rect 28353 40103 28411 40109
rect 28353 40069 28365 40103
rect 28399 40100 28411 40103
rect 29178 40100 29184 40112
rect 28399 40072 29184 40100
rect 28399 40069 28411 40072
rect 28353 40063 28411 40069
rect 29178 40060 29184 40072
rect 29236 40060 29242 40112
rect 30944 40100 30972 40140
rect 30852 40072 30972 40100
rect 22741 40035 22799 40041
rect 22741 40001 22753 40035
rect 22787 40001 22799 40035
rect 22741 39995 22799 40001
rect 22833 40035 22891 40041
rect 22833 40001 22845 40035
rect 22879 40001 22891 40035
rect 24682 40035 24740 40041
rect 24682 40032 24694 40035
rect 22833 39995 22891 40001
rect 23124 40004 24694 40032
rect 11517 39967 11575 39973
rect 10060 39936 11008 39964
rect 7193 39927 7251 39933
rect 10980 39840 11008 39936
rect 11517 39933 11529 39967
rect 11563 39933 11575 39967
rect 11517 39927 11575 39933
rect 8570 39828 8576 39840
rect 8531 39800 8576 39828
rect 8570 39788 8576 39800
rect 8628 39788 8634 39840
rect 9766 39828 9772 39840
rect 9727 39800 9772 39828
rect 9766 39788 9772 39800
rect 9824 39788 9830 39840
rect 10962 39828 10968 39840
rect 10923 39800 10968 39828
rect 10962 39788 10968 39800
rect 11020 39788 11026 39840
rect 11532 39828 11560 39927
rect 21910 39924 21916 39976
rect 21968 39964 21974 39976
rect 22756 39964 22784 39995
rect 23124 39973 23152 40004
rect 24682 40001 24694 40004
rect 24728 40001 24740 40035
rect 30558 40032 30564 40044
rect 30519 40004 30564 40032
rect 24682 39995 24740 40001
rect 30558 39992 30564 40004
rect 30616 39992 30622 40044
rect 30724 40041 30782 40047
rect 30852 40041 30880 40072
rect 31018 40041 31024 40044
rect 30724 40038 30736 40041
rect 30714 40007 30736 40038
rect 30770 40007 30782 40041
rect 30714 40001 30782 40007
rect 30837 40035 30895 40041
rect 30837 40001 30849 40035
rect 30883 40001 30895 40035
rect 21968 39936 22784 39964
rect 23109 39967 23167 39973
rect 21968 39924 21974 39936
rect 23109 39933 23121 39967
rect 23155 39933 23167 39967
rect 23109 39927 23167 39933
rect 24949 39967 25007 39973
rect 24949 39933 24961 39967
rect 24995 39964 25007 39967
rect 25038 39964 25044 39976
rect 24995 39936 25044 39964
rect 24995 39933 25007 39936
rect 24949 39927 25007 39933
rect 25038 39924 25044 39936
rect 25096 39924 25102 39976
rect 30714 39896 30742 40001
rect 30837 39995 30895 40001
rect 30975 40035 31024 40041
rect 30975 40001 30987 40035
rect 31021 40001 31024 40035
rect 30975 39995 31024 40001
rect 31018 39992 31024 39995
rect 31076 39992 31082 40044
rect 31110 39896 31116 39908
rect 30714 39868 31116 39896
rect 31110 39856 31116 39868
rect 31168 39856 31174 39908
rect 12618 39828 12624 39840
rect 11532 39800 12624 39828
rect 12618 39788 12624 39800
rect 12676 39788 12682 39840
rect 17402 39828 17408 39840
rect 17363 39800 17408 39828
rect 17402 39788 17408 39800
rect 17460 39788 17466 39840
rect 19242 39828 19248 39840
rect 19203 39800 19248 39828
rect 19242 39788 19248 39800
rect 19300 39788 19306 39840
rect 20257 39831 20315 39837
rect 20257 39797 20269 39831
rect 20303 39828 20315 39831
rect 20346 39828 20352 39840
rect 20303 39800 20352 39828
rect 20303 39797 20315 39800
rect 20257 39791 20315 39797
rect 20346 39788 20352 39800
rect 20404 39788 20410 39840
rect 21269 39831 21327 39837
rect 21269 39797 21281 39831
rect 21315 39828 21327 39831
rect 21818 39828 21824 39840
rect 21315 39800 21824 39828
rect 21315 39797 21327 39800
rect 21269 39791 21327 39797
rect 21818 39788 21824 39800
rect 21876 39788 21882 39840
rect 23382 39788 23388 39840
rect 23440 39828 23446 39840
rect 23569 39831 23627 39837
rect 23569 39828 23581 39831
rect 23440 39800 23581 39828
rect 23440 39788 23446 39800
rect 23569 39797 23581 39800
rect 23615 39797 23627 39831
rect 23569 39791 23627 39797
rect 27614 39788 27620 39840
rect 27672 39828 27678 39840
rect 27985 39831 28043 39837
rect 27985 39828 27997 39831
rect 27672 39800 27997 39828
rect 27672 39788 27678 39800
rect 27985 39797 27997 39800
rect 28031 39797 28043 39831
rect 30006 39828 30012 39840
rect 29967 39800 30012 39828
rect 27985 39791 28043 39797
rect 30006 39788 30012 39800
rect 30064 39828 30070 39840
rect 31018 39828 31024 39840
rect 30064 39800 31024 39828
rect 30064 39788 30070 39800
rect 31018 39788 31024 39800
rect 31076 39788 31082 39840
rect 31205 39831 31263 39837
rect 31205 39797 31217 39831
rect 31251 39828 31263 39831
rect 31294 39828 31300 39840
rect 31251 39800 31300 39828
rect 31251 39797 31263 39800
rect 31205 39791 31263 39797
rect 31294 39788 31300 39800
rect 31352 39788 31358 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 11054 39624 11060 39636
rect 7576 39596 11060 39624
rect 5810 39448 5816 39500
rect 5868 39488 5874 39500
rect 7576 39497 7604 39596
rect 11054 39584 11060 39596
rect 11112 39584 11118 39636
rect 11241 39627 11299 39633
rect 11241 39593 11253 39627
rect 11287 39624 11299 39627
rect 11698 39624 11704 39636
rect 11287 39596 11704 39624
rect 11287 39593 11299 39596
rect 11241 39587 11299 39593
rect 11698 39584 11704 39596
rect 11756 39584 11762 39636
rect 15470 39624 15476 39636
rect 15431 39596 15476 39624
rect 15470 39584 15476 39596
rect 15528 39584 15534 39636
rect 21358 39624 21364 39636
rect 21319 39596 21364 39624
rect 21358 39584 21364 39596
rect 21416 39584 21422 39636
rect 32674 39624 32680 39636
rect 31036 39596 32680 39624
rect 31036 39497 31064 39596
rect 32674 39584 32680 39596
rect 32732 39584 32738 39636
rect 6273 39491 6331 39497
rect 5868 39460 6224 39488
rect 5868 39448 5874 39460
rect 1854 39380 1860 39432
rect 1912 39420 1918 39432
rect 4433 39423 4491 39429
rect 4433 39420 4445 39423
rect 1912 39392 4445 39420
rect 1912 39380 1918 39392
rect 4433 39389 4445 39392
rect 4479 39420 4491 39423
rect 6086 39420 6092 39432
rect 4479 39392 6092 39420
rect 4479 39389 4491 39392
rect 4433 39383 4491 39389
rect 6086 39380 6092 39392
rect 6144 39380 6150 39432
rect 6196 39420 6224 39460
rect 6273 39457 6285 39491
rect 6319 39488 6331 39491
rect 7561 39491 7619 39497
rect 7561 39488 7573 39491
rect 6319 39460 7573 39488
rect 6319 39457 6331 39460
rect 6273 39451 6331 39457
rect 7561 39457 7573 39460
rect 7607 39457 7619 39491
rect 7561 39451 7619 39457
rect 31021 39491 31079 39497
rect 31021 39457 31033 39491
rect 31067 39457 31079 39491
rect 31021 39451 31079 39457
rect 6549 39423 6607 39429
rect 6549 39420 6561 39423
rect 6196 39392 6561 39420
rect 6549 39389 6561 39392
rect 6595 39389 6607 39423
rect 6549 39383 6607 39389
rect 9030 39380 9036 39432
rect 9088 39420 9094 39432
rect 9125 39423 9183 39429
rect 9125 39420 9137 39423
rect 9088 39392 9137 39420
rect 9088 39380 9094 39392
rect 9125 39389 9137 39392
rect 9171 39389 9183 39423
rect 9125 39383 9183 39389
rect 9392 39423 9450 39429
rect 9392 39389 9404 39423
rect 9438 39420 9450 39423
rect 9766 39420 9772 39432
rect 9438 39392 9772 39420
rect 9438 39389 9450 39392
rect 9392 39383 9450 39389
rect 9766 39380 9772 39392
rect 9824 39380 9830 39432
rect 12342 39420 12348 39432
rect 12400 39429 12406 39432
rect 12312 39392 12348 39420
rect 12342 39380 12348 39392
rect 12400 39383 12412 39429
rect 12618 39420 12624 39432
rect 12531 39392 12624 39420
rect 12400 39380 12406 39383
rect 12618 39380 12624 39392
rect 12676 39420 12682 39432
rect 13262 39420 13268 39432
rect 12676 39392 13268 39420
rect 12676 39380 12682 39392
rect 13262 39380 13268 39392
rect 13320 39380 13326 39432
rect 16114 39380 16120 39432
rect 16172 39420 16178 39432
rect 16853 39423 16911 39429
rect 16853 39420 16865 39423
rect 16172 39392 16865 39420
rect 16172 39380 16178 39392
rect 16853 39389 16865 39392
rect 16899 39420 16911 39423
rect 18138 39420 18144 39432
rect 16899 39392 18144 39420
rect 16899 39389 16911 39392
rect 16853 39383 16911 39389
rect 18138 39380 18144 39392
rect 18196 39420 18202 39432
rect 19242 39420 19248 39432
rect 18196 39392 19248 39420
rect 18196 39380 18202 39392
rect 19242 39380 19248 39392
rect 19300 39380 19306 39432
rect 19518 39429 19524 39432
rect 19512 39420 19524 39429
rect 19479 39392 19524 39420
rect 19512 39383 19524 39392
rect 19518 39380 19524 39383
rect 19576 39380 19582 39432
rect 21634 39420 21640 39432
rect 21595 39392 21640 39420
rect 21634 39380 21640 39392
rect 21692 39380 21698 39432
rect 21729 39423 21787 39429
rect 21729 39389 21741 39423
rect 21775 39389 21787 39423
rect 21729 39383 21787 39389
rect 4700 39355 4758 39361
rect 4700 39321 4712 39355
rect 4746 39352 4758 39355
rect 5166 39352 5172 39364
rect 4746 39324 5172 39352
rect 4746 39321 4758 39324
rect 4700 39315 4758 39321
rect 5166 39312 5172 39324
rect 5224 39312 5230 39364
rect 16574 39352 16580 39364
rect 16632 39361 16638 39364
rect 16544 39324 16580 39352
rect 16574 39312 16580 39324
rect 16632 39315 16644 39361
rect 21744 39352 21772 39383
rect 21818 39380 21824 39432
rect 21876 39420 21882 39432
rect 22005 39423 22063 39429
rect 21876 39392 21921 39420
rect 21876 39380 21882 39392
rect 22005 39389 22017 39423
rect 22051 39420 22063 39423
rect 22278 39420 22284 39432
rect 22051 39392 22284 39420
rect 22051 39389 22063 39392
rect 22005 39383 22063 39389
rect 22278 39380 22284 39392
rect 22336 39380 22342 39432
rect 23845 39423 23903 39429
rect 23845 39389 23857 39423
rect 23891 39420 23903 39423
rect 25038 39420 25044 39432
rect 23891 39392 25044 39420
rect 23891 39389 23903 39392
rect 23845 39383 23903 39389
rect 25038 39380 25044 39392
rect 25096 39380 25102 39432
rect 27157 39423 27215 39429
rect 27157 39389 27169 39423
rect 27203 39420 27215 39423
rect 27246 39420 27252 39432
rect 27203 39392 27252 39420
rect 27203 39389 27215 39392
rect 27157 39383 27215 39389
rect 27246 39380 27252 39392
rect 27304 39380 27310 39432
rect 31294 39429 31300 39432
rect 31288 39420 31300 39429
rect 31255 39392 31300 39420
rect 31288 39383 31300 39392
rect 31294 39380 31300 39383
rect 31352 39380 31358 39432
rect 21910 39352 21916 39364
rect 21744 39324 21916 39352
rect 16632 39312 16638 39315
rect 21910 39312 21916 39324
rect 21968 39312 21974 39364
rect 23474 39312 23480 39364
rect 23532 39352 23538 39364
rect 23578 39355 23636 39361
rect 23578 39352 23590 39355
rect 23532 39324 23590 39352
rect 23532 39312 23538 39324
rect 23578 39321 23590 39324
rect 23624 39321 23636 39355
rect 23578 39315 23636 39321
rect 27424 39355 27482 39361
rect 27424 39321 27436 39355
rect 27470 39352 27482 39355
rect 27522 39352 27528 39364
rect 27470 39324 27528 39352
rect 27470 39321 27482 39324
rect 27424 39315 27482 39321
rect 27522 39312 27528 39324
rect 27580 39312 27586 39364
rect 30558 39312 30564 39364
rect 30616 39352 30622 39364
rect 31018 39352 31024 39364
rect 30616 39324 31024 39352
rect 30616 39312 30622 39324
rect 31018 39312 31024 39324
rect 31076 39312 31082 39364
rect 5813 39287 5871 39293
rect 5813 39253 5825 39287
rect 5859 39284 5871 39287
rect 6638 39284 6644 39296
rect 5859 39256 6644 39284
rect 5859 39253 5871 39256
rect 5813 39247 5871 39253
rect 6638 39244 6644 39256
rect 6696 39244 6702 39296
rect 10502 39284 10508 39296
rect 10463 39256 10508 39284
rect 10502 39244 10508 39256
rect 10560 39244 10566 39296
rect 20070 39244 20076 39296
rect 20128 39284 20134 39296
rect 20625 39287 20683 39293
rect 20625 39284 20637 39287
rect 20128 39256 20637 39284
rect 20128 39244 20134 39256
rect 20625 39253 20637 39256
rect 20671 39253 20683 39287
rect 20625 39247 20683 39253
rect 22465 39287 22523 39293
rect 22465 39253 22477 39287
rect 22511 39284 22523 39287
rect 22646 39284 22652 39296
rect 22511 39256 22652 39284
rect 22511 39253 22523 39256
rect 22465 39247 22523 39253
rect 22646 39244 22652 39256
rect 22704 39244 22710 39296
rect 28537 39287 28595 39293
rect 28537 39253 28549 39287
rect 28583 39284 28595 39287
rect 28810 39284 28816 39296
rect 28583 39256 28816 39284
rect 28583 39253 28595 39256
rect 28537 39247 28595 39253
rect 28810 39244 28816 39256
rect 28868 39244 28874 39296
rect 28994 39244 29000 39296
rect 29052 39284 29058 39296
rect 29733 39287 29791 39293
rect 29733 39284 29745 39287
rect 29052 39256 29745 39284
rect 29052 39244 29058 39256
rect 29733 39253 29745 39256
rect 29779 39253 29791 39287
rect 30374 39284 30380 39296
rect 30335 39256 30380 39284
rect 29733 39247 29791 39253
rect 30374 39244 30380 39256
rect 30432 39244 30438 39296
rect 31294 39244 31300 39296
rect 31352 39284 31358 39296
rect 32401 39287 32459 39293
rect 32401 39284 32413 39287
rect 31352 39256 32413 39284
rect 31352 39244 31358 39256
rect 32401 39253 32413 39256
rect 32447 39253 32459 39287
rect 32401 39247 32459 39253
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 5166 39080 5172 39092
rect 5127 39052 5172 39080
rect 5166 39040 5172 39052
rect 5224 39040 5230 39092
rect 5258 39040 5264 39092
rect 5316 39080 5322 39092
rect 5316 39052 9812 39080
rect 5316 39040 5322 39052
rect 4709 39015 4767 39021
rect 4709 38981 4721 39015
rect 4755 39012 4767 39015
rect 5994 39012 6000 39024
rect 4755 38984 6000 39012
rect 4755 38981 4767 38984
rect 4709 38975 4767 38981
rect 3047 38953 3053 38956
rect 2941 38947 2999 38953
rect 2941 38944 2953 38947
rect 2884 38916 2953 38944
rect 2884 38820 2912 38916
rect 2941 38913 2953 38916
rect 2987 38913 2999 38947
rect 2941 38907 2999 38913
rect 3034 38947 3053 38953
rect 3034 38913 3046 38947
rect 3034 38907 3053 38913
rect 3047 38904 3053 38907
rect 3105 38904 3111 38956
rect 3142 38904 3148 38956
rect 3200 38953 3206 38956
rect 3200 38944 3208 38953
rect 3326 38944 3332 38956
rect 3200 38916 3245 38944
rect 3287 38916 3332 38944
rect 3200 38907 3208 38916
rect 3200 38904 3206 38907
rect 3326 38904 3332 38916
rect 3384 38904 3390 38956
rect 5276 38950 5304 38984
rect 5994 38972 6000 38984
rect 6052 38972 6058 39024
rect 6086 38972 6092 39024
rect 6144 39012 6150 39024
rect 9030 39012 9036 39024
rect 6144 38984 9036 39012
rect 6144 38972 6150 38984
rect 5445 38950 5503 38953
rect 5276 38947 5503 38950
rect 5276 38922 5457 38947
rect 5445 38913 5457 38922
rect 5491 38913 5503 38947
rect 5445 38907 5503 38913
rect 5534 38947 5592 38953
rect 5534 38913 5546 38947
rect 5580 38913 5592 38947
rect 5534 38907 5592 38913
rect 5629 38947 5687 38953
rect 5629 38913 5641 38947
rect 5675 38913 5687 38947
rect 5629 38907 5687 38913
rect 3068 38876 3096 38904
rect 5549 38876 5577 38907
rect 3068 38848 5577 38876
rect 5644 38876 5672 38907
rect 5810 38904 5816 38956
rect 5868 38944 5874 38956
rect 6549 38947 6607 38953
rect 5868 38916 5913 38944
rect 5868 38904 5874 38916
rect 6549 38913 6561 38947
rect 6595 38944 6607 38947
rect 6638 38944 6644 38956
rect 6595 38916 6644 38944
rect 6595 38913 6607 38916
rect 6549 38907 6607 38913
rect 6638 38904 6644 38916
rect 6696 38904 6702 38956
rect 6730 38904 6736 38956
rect 6788 38944 6794 38956
rect 8956 38953 8984 38984
rect 9030 38972 9036 38984
rect 9088 38972 9094 39024
rect 9208 39015 9266 39021
rect 9208 38981 9220 39015
rect 9254 39012 9266 39015
rect 9674 39012 9680 39024
rect 9254 38984 9680 39012
rect 9254 38981 9266 38984
rect 9208 38975 9266 38981
rect 9674 38972 9680 38984
rect 9732 38972 9738 39024
rect 9784 39012 9812 39052
rect 12434 39040 12440 39092
rect 12492 39080 12498 39092
rect 12621 39083 12679 39089
rect 12621 39080 12633 39083
rect 12492 39052 12633 39080
rect 12492 39040 12498 39052
rect 12621 39049 12633 39052
rect 12667 39049 12679 39083
rect 12621 39043 12679 39049
rect 22094 39040 22100 39092
rect 22152 39080 22158 39092
rect 22152 39052 22508 39080
rect 22152 39040 22158 39052
rect 22480 39021 22508 39052
rect 22738 39040 22744 39092
rect 22796 39080 22802 39092
rect 22833 39083 22891 39089
rect 22833 39080 22845 39083
rect 22796 39052 22845 39080
rect 22796 39040 22802 39052
rect 22833 39049 22845 39052
rect 22879 39049 22891 39083
rect 27154 39080 27160 39092
rect 27115 39052 27160 39080
rect 22833 39043 22891 39049
rect 27154 39040 27160 39052
rect 27212 39040 27218 39092
rect 27890 39080 27896 39092
rect 27586 39052 27896 39080
rect 22465 39015 22523 39021
rect 9784 38984 22094 39012
rect 8941 38947 8999 38953
rect 6788 38916 6833 38944
rect 7668 38916 8892 38944
rect 6788 38904 6794 38916
rect 7668 38888 7696 38916
rect 6365 38879 6423 38885
rect 6365 38876 6377 38879
rect 5644 38848 6377 38876
rect 2866 38768 2872 38820
rect 2924 38808 2930 38820
rect 3881 38811 3939 38817
rect 3881 38808 3893 38811
rect 2924 38780 3893 38808
rect 2924 38768 2930 38780
rect 3881 38777 3893 38780
rect 3927 38808 3939 38811
rect 5258 38808 5264 38820
rect 3927 38780 5264 38808
rect 3927 38777 3939 38780
rect 3881 38771 3939 38777
rect 5258 38768 5264 38780
rect 5316 38768 5322 38820
rect 5442 38768 5448 38820
rect 5500 38808 5506 38820
rect 5549 38808 5577 38848
rect 6365 38845 6377 38848
rect 6411 38845 6423 38879
rect 6365 38839 6423 38845
rect 7469 38879 7527 38885
rect 7469 38845 7481 38879
rect 7515 38876 7527 38879
rect 7650 38876 7656 38888
rect 7515 38848 7656 38876
rect 7515 38845 7527 38848
rect 7469 38839 7527 38845
rect 7650 38836 7656 38848
rect 7708 38836 7714 38888
rect 7745 38879 7803 38885
rect 7745 38845 7757 38879
rect 7791 38845 7803 38879
rect 8864 38876 8892 38916
rect 8941 38913 8953 38947
rect 8987 38913 8999 38947
rect 12437 38947 12495 38953
rect 8941 38907 8999 38913
rect 9048 38916 9996 38944
rect 9048 38876 9076 38916
rect 8864 38848 9076 38876
rect 9968 38876 9996 38916
rect 12437 38913 12449 38947
rect 12483 38944 12495 38947
rect 12526 38944 12532 38956
rect 12483 38916 12532 38944
rect 12483 38913 12495 38916
rect 12437 38907 12495 38913
rect 12526 38904 12532 38916
rect 12584 38904 12590 38956
rect 13449 38947 13507 38953
rect 13449 38913 13461 38947
rect 13495 38944 13507 38947
rect 15562 38944 15568 38956
rect 13495 38916 15568 38944
rect 13495 38913 13507 38916
rect 13449 38907 13507 38913
rect 15562 38904 15568 38916
rect 15620 38904 15626 38956
rect 13173 38879 13231 38885
rect 13173 38876 13185 38879
rect 9968 38848 13185 38876
rect 7745 38839 7803 38845
rect 13173 38845 13185 38848
rect 13219 38845 13231 38879
rect 22066 38876 22094 38984
rect 22465 38981 22477 39015
rect 22511 39012 22523 39015
rect 23014 39012 23020 39024
rect 22511 38984 23020 39012
rect 22511 38981 22523 38984
rect 22465 38975 22523 38981
rect 23014 38972 23020 38984
rect 23072 38972 23078 39024
rect 24946 38972 24952 39024
rect 25004 39012 25010 39024
rect 27586 39012 27614 39052
rect 27890 39040 27896 39052
rect 27948 39080 27954 39092
rect 30834 39080 30840 39092
rect 27948 39052 30840 39080
rect 27948 39040 27954 39052
rect 30834 39040 30840 39052
rect 30892 39040 30898 39092
rect 32125 39015 32183 39021
rect 32125 39012 32137 39015
rect 25004 38984 25544 39012
rect 25004 38972 25010 38984
rect 22646 38904 22652 38956
rect 22704 38944 22710 38956
rect 23290 38944 23296 38956
rect 22704 38916 23296 38944
rect 22704 38904 22710 38916
rect 23290 38904 23296 38916
rect 23348 38904 23354 38956
rect 24578 38904 24584 38956
rect 24636 38944 24642 38956
rect 25225 38947 25283 38953
rect 25225 38944 25237 38947
rect 24636 38916 25237 38944
rect 24636 38904 24642 38916
rect 25225 38913 25237 38916
rect 25271 38913 25283 38947
rect 25406 38944 25412 38956
rect 25367 38916 25412 38944
rect 25225 38907 25283 38913
rect 25406 38904 25412 38916
rect 25464 38904 25470 38956
rect 25516 38953 25544 38984
rect 27540 38984 27614 39012
rect 30944 38984 32137 39012
rect 25501 38947 25559 38953
rect 25501 38913 25513 38947
rect 25547 38913 25559 38947
rect 25501 38907 25559 38913
rect 25590 38904 25596 38956
rect 25648 38944 25654 38956
rect 27540 38953 27568 38984
rect 30944 38956 30972 38984
rect 32125 38981 32137 38984
rect 32171 38981 32183 39015
rect 32125 38975 32183 38981
rect 27433 38947 27491 38953
rect 27433 38944 27445 38947
rect 25648 38916 25693 38944
rect 26344 38916 27445 38944
rect 25648 38904 25654 38916
rect 26344 38885 26372 38916
rect 27433 38913 27445 38916
rect 27479 38913 27491 38947
rect 27433 38907 27491 38913
rect 27525 38947 27583 38953
rect 27525 38913 27537 38947
rect 27571 38913 27583 38947
rect 27525 38907 27583 38913
rect 26329 38879 26387 38885
rect 26329 38876 26341 38879
rect 22066 38848 26341 38876
rect 13173 38839 13231 38845
rect 26329 38845 26341 38848
rect 26375 38845 26387 38879
rect 27448 38876 27476 38907
rect 27614 38904 27620 38956
rect 27672 38944 27678 38956
rect 27801 38947 27859 38953
rect 27672 38916 27717 38944
rect 27672 38904 27678 38916
rect 27801 38913 27813 38947
rect 27847 38944 27859 38947
rect 28074 38944 28080 38956
rect 27847 38916 28080 38944
rect 27847 38913 27859 38916
rect 27801 38907 27859 38913
rect 28074 38904 28080 38916
rect 28132 38904 28138 38956
rect 28261 38947 28319 38953
rect 28261 38913 28273 38947
rect 28307 38944 28319 38947
rect 28994 38944 29000 38956
rect 28307 38916 29000 38944
rect 28307 38913 28319 38916
rect 28261 38907 28319 38913
rect 28994 38904 29000 38916
rect 29052 38904 29058 38956
rect 30374 38904 30380 38956
rect 30432 38944 30438 38956
rect 30725 38947 30783 38953
rect 30725 38944 30737 38947
rect 30432 38916 30737 38944
rect 30432 38904 30438 38916
rect 30725 38913 30737 38916
rect 30771 38913 30783 38947
rect 30725 38907 30783 38913
rect 30834 38947 30892 38953
rect 30834 38913 30846 38947
rect 30880 38913 30892 38947
rect 30834 38907 30892 38913
rect 30929 38950 30987 38956
rect 30929 38916 30941 38950
rect 30975 38916 30987 38950
rect 30929 38910 30987 38916
rect 27706 38876 27712 38888
rect 27448 38848 27712 38876
rect 26329 38839 26387 38845
rect 7760 38808 7788 38839
rect 27706 38836 27712 38848
rect 27764 38836 27770 38888
rect 30852 38820 30880 38907
rect 31018 38904 31024 38956
rect 31076 38944 31082 38956
rect 31113 38947 31171 38953
rect 31113 38944 31125 38947
rect 31076 38916 31125 38944
rect 31076 38904 31082 38916
rect 31113 38913 31125 38916
rect 31159 38944 31171 38947
rect 31570 38944 31576 38956
rect 31159 38916 31576 38944
rect 31159 38913 31171 38916
rect 31113 38907 31171 38913
rect 31570 38904 31576 38916
rect 31628 38904 31634 38956
rect 31754 38904 31760 38956
rect 31812 38944 31818 38956
rect 32309 38947 32367 38953
rect 32309 38944 32321 38947
rect 31812 38916 32321 38944
rect 31812 38904 31818 38916
rect 32309 38913 32321 38916
rect 32355 38913 32367 38947
rect 32309 38907 32367 38913
rect 32493 38947 32551 38953
rect 32493 38913 32505 38947
rect 32539 38944 32551 38947
rect 32766 38944 32772 38956
rect 32539 38916 32772 38944
rect 32539 38913 32551 38916
rect 32493 38907 32551 38913
rect 32766 38904 32772 38916
rect 32824 38904 32830 38956
rect 16298 38808 16304 38820
rect 5500 38780 7788 38808
rect 13740 38780 16304 38808
rect 5500 38768 5506 38780
rect 2682 38740 2688 38752
rect 2643 38712 2688 38740
rect 2682 38700 2688 38712
rect 2740 38700 2746 38752
rect 3326 38700 3332 38752
rect 3384 38740 3390 38752
rect 4798 38740 4804 38752
rect 3384 38712 4804 38740
rect 3384 38700 3390 38712
rect 4798 38700 4804 38712
rect 4856 38740 4862 38752
rect 5810 38740 5816 38752
rect 4856 38712 5816 38740
rect 4856 38700 4862 38712
rect 5810 38700 5816 38712
rect 5868 38700 5874 38752
rect 10318 38740 10324 38752
rect 10279 38712 10324 38740
rect 10318 38700 10324 38712
rect 10376 38700 10382 38752
rect 10962 38700 10968 38752
rect 11020 38740 11026 38752
rect 13740 38740 13768 38780
rect 16298 38768 16304 38780
rect 16356 38808 16362 38820
rect 20622 38808 20628 38820
rect 16356 38780 20628 38808
rect 16356 38768 16362 38780
rect 20622 38768 20628 38780
rect 20680 38768 20686 38820
rect 30834 38768 30840 38820
rect 30892 38768 30898 38820
rect 58158 38808 58164 38820
rect 58119 38780 58164 38808
rect 58158 38768 58164 38780
rect 58216 38768 58222 38820
rect 11020 38712 13768 38740
rect 11020 38700 11026 38712
rect 13814 38700 13820 38752
rect 13872 38740 13878 38752
rect 19426 38740 19432 38752
rect 13872 38712 19432 38740
rect 13872 38700 13878 38712
rect 19426 38700 19432 38712
rect 19484 38700 19490 38752
rect 21634 38700 21640 38752
rect 21692 38740 21698 38752
rect 21913 38743 21971 38749
rect 21913 38740 21925 38743
rect 21692 38712 21925 38740
rect 21692 38700 21698 38712
rect 21913 38709 21925 38712
rect 21959 38709 21971 38743
rect 24762 38740 24768 38752
rect 24675 38712 24768 38740
rect 21913 38703 21971 38709
rect 24762 38700 24768 38712
rect 24820 38740 24826 38752
rect 25222 38740 25228 38752
rect 24820 38712 25228 38740
rect 24820 38700 24826 38712
rect 25222 38700 25228 38712
rect 25280 38740 25286 38752
rect 25590 38740 25596 38752
rect 25280 38712 25596 38740
rect 25280 38700 25286 38712
rect 25590 38700 25596 38712
rect 25648 38700 25654 38752
rect 25869 38743 25927 38749
rect 25869 38709 25881 38743
rect 25915 38740 25927 38743
rect 25958 38740 25964 38752
rect 25915 38712 25964 38740
rect 25915 38709 25927 38712
rect 25869 38703 25927 38709
rect 25958 38700 25964 38712
rect 26016 38700 26022 38752
rect 29086 38700 29092 38752
rect 29144 38740 29150 38752
rect 29549 38743 29607 38749
rect 29549 38740 29561 38743
rect 29144 38712 29561 38740
rect 29144 38700 29150 38712
rect 29549 38709 29561 38712
rect 29595 38709 29607 38743
rect 30466 38740 30472 38752
rect 30427 38712 30472 38740
rect 29549 38703 29607 38709
rect 30466 38700 30472 38712
rect 30524 38700 30530 38752
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 6086 38496 6092 38548
rect 6144 38536 6150 38548
rect 6549 38539 6607 38545
rect 6549 38536 6561 38539
rect 6144 38508 6561 38536
rect 6144 38496 6150 38508
rect 6549 38505 6561 38508
rect 6595 38505 6607 38539
rect 6549 38499 6607 38505
rect 6730 38496 6736 38548
rect 6788 38536 6794 38548
rect 7929 38539 7987 38545
rect 7929 38536 7941 38539
rect 6788 38508 7941 38536
rect 6788 38496 6794 38508
rect 7929 38505 7941 38508
rect 7975 38505 7987 38539
rect 7929 38499 7987 38505
rect 9125 38539 9183 38545
rect 9125 38505 9137 38539
rect 9171 38536 9183 38539
rect 9398 38536 9404 38548
rect 9171 38508 9404 38536
rect 9171 38505 9183 38508
rect 9125 38499 9183 38505
rect 9398 38496 9404 38508
rect 9456 38496 9462 38548
rect 27522 38536 27528 38548
rect 27483 38508 27528 38536
rect 27522 38496 27528 38508
rect 27580 38496 27586 38548
rect 14645 38471 14703 38477
rect 14645 38437 14657 38471
rect 14691 38468 14703 38471
rect 19242 38468 19248 38480
rect 14691 38440 19248 38468
rect 14691 38437 14703 38440
rect 14645 38431 14703 38437
rect 19242 38428 19248 38440
rect 19300 38428 19306 38480
rect 19889 38471 19947 38477
rect 19889 38437 19901 38471
rect 19935 38468 19947 38471
rect 21082 38468 21088 38480
rect 19935 38440 21088 38468
rect 19935 38437 19947 38440
rect 19889 38431 19947 38437
rect 21082 38428 21088 38440
rect 21140 38428 21146 38480
rect 24946 38468 24952 38480
rect 24872 38440 24952 38468
rect 12526 38400 12532 38412
rect 8128 38372 12532 38400
rect 1854 38332 1860 38344
rect 1815 38304 1860 38332
rect 1854 38292 1860 38304
rect 1912 38292 1918 38344
rect 2124 38335 2182 38341
rect 2124 38301 2136 38335
rect 2170 38332 2182 38335
rect 2682 38332 2688 38344
rect 2170 38304 2688 38332
rect 2170 38301 2182 38304
rect 2124 38295 2182 38301
rect 2682 38292 2688 38304
rect 2740 38292 2746 38344
rect 8128 38341 8156 38372
rect 12526 38360 12532 38372
rect 12584 38360 12590 38412
rect 19150 38400 19156 38412
rect 18893 38372 19156 38400
rect 8113 38335 8171 38341
rect 8113 38301 8125 38335
rect 8159 38301 8171 38335
rect 8113 38295 8171 38301
rect 8570 38292 8576 38344
rect 8628 38332 8634 38344
rect 9306 38332 9312 38344
rect 8628 38304 9312 38332
rect 8628 38292 8634 38304
rect 9306 38292 9312 38304
rect 9364 38292 9370 38344
rect 10318 38292 10324 38344
rect 10376 38332 10382 38344
rect 14093 38335 14151 38341
rect 14093 38332 14105 38335
rect 10376 38304 14105 38332
rect 10376 38292 10382 38304
rect 14093 38301 14105 38304
rect 14139 38301 14151 38335
rect 14461 38335 14519 38341
rect 14461 38332 14473 38335
rect 14093 38295 14151 38301
rect 14200 38304 14473 38332
rect 5261 38267 5319 38273
rect 5261 38233 5273 38267
rect 5307 38264 5319 38267
rect 6730 38264 6736 38276
rect 5307 38236 6736 38264
rect 5307 38233 5319 38236
rect 5261 38227 5319 38233
rect 6730 38224 6736 38236
rect 6788 38224 6794 38276
rect 9493 38267 9551 38273
rect 9493 38233 9505 38267
rect 9539 38264 9551 38267
rect 9674 38264 9680 38276
rect 9539 38236 9680 38264
rect 9539 38233 9551 38236
rect 9493 38227 9551 38233
rect 9674 38224 9680 38236
rect 9732 38264 9738 38276
rect 10870 38264 10876 38276
rect 9732 38236 10876 38264
rect 9732 38224 9738 38236
rect 10870 38224 10876 38236
rect 10928 38224 10934 38276
rect 13630 38224 13636 38276
rect 13688 38264 13694 38276
rect 14200 38264 14228 38304
rect 14461 38301 14473 38304
rect 14507 38301 14519 38335
rect 17586 38332 17592 38344
rect 17547 38304 17592 38332
rect 14461 38295 14519 38301
rect 17586 38292 17592 38304
rect 17644 38292 17650 38344
rect 17678 38292 17684 38344
rect 17736 38332 17742 38344
rect 17954 38332 17960 38344
rect 17736 38304 17781 38332
rect 17915 38304 17960 38332
rect 17736 38292 17742 38304
rect 17954 38292 17960 38304
rect 18012 38292 18018 38344
rect 18095 38335 18153 38341
rect 18095 38301 18107 38335
rect 18141 38332 18153 38335
rect 18893 38332 18921 38372
rect 19150 38360 19156 38372
rect 19208 38400 19214 38412
rect 19208 38372 19564 38400
rect 19208 38360 19214 38372
rect 19242 38332 19248 38344
rect 18141 38304 18921 38332
rect 19203 38304 19248 38332
rect 18141 38301 18153 38304
rect 18095 38295 18153 38301
rect 19242 38292 19248 38304
rect 19300 38292 19306 38344
rect 19334 38292 19340 38344
rect 19392 38332 19398 38344
rect 19536 38332 19564 38372
rect 19710 38335 19768 38341
rect 19710 38332 19722 38335
rect 19392 38304 19437 38332
rect 19536 38304 19722 38332
rect 19392 38292 19398 38304
rect 19710 38301 19722 38304
rect 19756 38301 19768 38335
rect 19710 38295 19768 38301
rect 20346 38292 20352 38344
rect 20404 38332 20410 38344
rect 24578 38332 24584 38344
rect 20404 38304 22094 38332
rect 24539 38304 24584 38332
rect 20404 38292 20410 38304
rect 13688 38236 14228 38264
rect 14277 38267 14335 38273
rect 13688 38224 13694 38236
rect 14277 38233 14289 38267
rect 14323 38233 14335 38267
rect 14277 38227 14335 38233
rect 14369 38267 14427 38273
rect 14369 38233 14381 38267
rect 14415 38264 14427 38267
rect 15470 38264 15476 38276
rect 14415 38236 15476 38264
rect 14415 38233 14427 38236
rect 14369 38227 14427 38233
rect 3237 38199 3295 38205
rect 3237 38165 3249 38199
rect 3283 38196 3295 38199
rect 5074 38196 5080 38208
rect 3283 38168 5080 38196
rect 3283 38165 3295 38168
rect 3237 38159 3295 38165
rect 5074 38156 5080 38168
rect 5132 38156 5138 38208
rect 13722 38156 13728 38208
rect 13780 38196 13786 38208
rect 14292 38196 14320 38227
rect 15470 38224 15476 38236
rect 15528 38224 15534 38276
rect 17865 38267 17923 38273
rect 17865 38233 17877 38267
rect 17911 38264 17923 38267
rect 19521 38267 19579 38273
rect 19521 38264 19533 38267
rect 17911 38236 19533 38264
rect 17911 38233 17923 38236
rect 17865 38227 17923 38233
rect 19260 38208 19288 38236
rect 19521 38233 19533 38236
rect 19567 38233 19579 38267
rect 19521 38227 19579 38233
rect 19613 38267 19671 38273
rect 19613 38233 19625 38267
rect 19659 38264 19671 38267
rect 20070 38264 20076 38276
rect 19659 38236 20076 38264
rect 19659 38233 19671 38236
rect 19613 38227 19671 38233
rect 20070 38224 20076 38236
rect 20128 38224 20134 38276
rect 20530 38264 20536 38276
rect 20491 38236 20536 38264
rect 20530 38224 20536 38236
rect 20588 38224 20594 38276
rect 20714 38264 20720 38276
rect 20675 38236 20720 38264
rect 20714 38224 20720 38236
rect 20772 38224 20778 38276
rect 13780 38168 14320 38196
rect 18233 38199 18291 38205
rect 13780 38156 13786 38168
rect 18233 38165 18245 38199
rect 18279 38196 18291 38199
rect 18598 38196 18604 38208
rect 18279 38168 18604 38196
rect 18279 38165 18291 38168
rect 18233 38159 18291 38165
rect 18598 38156 18604 38168
rect 18656 38156 18662 38208
rect 19242 38156 19248 38208
rect 19300 38156 19306 38208
rect 20162 38156 20168 38208
rect 20220 38196 20226 38208
rect 20349 38199 20407 38205
rect 20349 38196 20361 38199
rect 20220 38168 20361 38196
rect 20220 38156 20226 38168
rect 20349 38165 20361 38168
rect 20395 38165 20407 38199
rect 22066 38196 22094 38304
rect 24578 38292 24584 38304
rect 24636 38292 24642 38344
rect 24762 38332 24768 38344
rect 24723 38304 24768 38332
rect 24762 38292 24768 38304
rect 24820 38292 24826 38344
rect 24872 38341 24900 38440
rect 24946 38428 24952 38440
rect 25004 38428 25010 38480
rect 27890 38428 27896 38480
rect 27948 38428 27954 38480
rect 24857 38335 24915 38341
rect 24857 38301 24869 38335
rect 24903 38301 24915 38335
rect 24857 38295 24915 38301
rect 24949 38335 25007 38341
rect 24949 38301 24961 38335
rect 24995 38301 25007 38335
rect 25682 38332 25688 38344
rect 25643 38304 25688 38332
rect 24949 38295 25007 38301
rect 24964 38264 24992 38295
rect 25682 38292 25688 38304
rect 25740 38292 25746 38344
rect 25958 38341 25964 38344
rect 25952 38332 25964 38341
rect 25919 38304 25964 38332
rect 25952 38295 25964 38304
rect 25958 38292 25964 38295
rect 26016 38292 26022 38344
rect 27338 38292 27344 38344
rect 27396 38332 27402 38344
rect 27905 38341 27933 38428
rect 29086 38360 29092 38412
rect 29144 38400 29150 38412
rect 30193 38403 30251 38409
rect 30193 38400 30205 38403
rect 29144 38372 30205 38400
rect 29144 38360 29150 38372
rect 30193 38369 30205 38372
rect 30239 38369 30251 38403
rect 30193 38363 30251 38369
rect 27801 38335 27859 38341
rect 27801 38332 27813 38335
rect 27396 38304 27813 38332
rect 27396 38292 27402 38304
rect 27801 38301 27813 38304
rect 27847 38301 27859 38335
rect 27801 38295 27859 38301
rect 27890 38335 27948 38341
rect 27890 38301 27902 38335
rect 27936 38301 27948 38335
rect 27890 38295 27948 38301
rect 27985 38335 28043 38341
rect 27985 38301 27997 38335
rect 28031 38301 28043 38335
rect 27985 38295 28043 38301
rect 24688 38236 24992 38264
rect 28000 38264 28028 38295
rect 28074 38292 28080 38344
rect 28132 38332 28138 38344
rect 28169 38335 28227 38341
rect 28169 38332 28181 38335
rect 28132 38304 28181 38332
rect 28132 38292 28138 38304
rect 28169 38301 28181 38304
rect 28215 38332 28227 38335
rect 28997 38335 29055 38341
rect 28215 38304 28948 38332
rect 28215 38301 28227 38304
rect 28169 38295 28227 38301
rect 28629 38267 28687 38273
rect 28629 38264 28641 38267
rect 28000 38236 28641 38264
rect 24688 38208 24716 38236
rect 28629 38233 28641 38236
rect 28675 38233 28687 38267
rect 28810 38264 28816 38276
rect 28771 38236 28816 38264
rect 28629 38227 28687 38233
rect 28810 38224 28816 38236
rect 28868 38224 28874 38276
rect 28920 38264 28948 38304
rect 28997 38301 29009 38335
rect 29043 38332 29055 38335
rect 29178 38332 29184 38344
rect 29043 38304 29184 38332
rect 29043 38301 29055 38304
rect 28997 38295 29055 38301
rect 29178 38292 29184 38304
rect 29236 38292 29242 38344
rect 30466 38341 30472 38344
rect 30460 38332 30472 38341
rect 30427 38304 30472 38332
rect 30460 38295 30472 38304
rect 30466 38292 30472 38295
rect 30524 38292 30530 38344
rect 32674 38332 32680 38344
rect 32587 38304 32680 38332
rect 32674 38292 32680 38304
rect 32732 38332 32738 38344
rect 32732 38304 33180 38332
rect 32732 38292 32738 38304
rect 33152 38276 33180 38304
rect 30558 38264 30564 38276
rect 28920 38236 30564 38264
rect 30558 38224 30564 38236
rect 30616 38224 30622 38276
rect 32944 38267 33002 38273
rect 32944 38233 32956 38267
rect 32990 38264 33002 38267
rect 33042 38264 33048 38276
rect 32990 38236 33048 38264
rect 32990 38233 33002 38236
rect 32944 38227 33002 38233
rect 33042 38224 33048 38236
rect 33100 38224 33106 38276
rect 33134 38224 33140 38276
rect 33192 38224 33198 38276
rect 23845 38199 23903 38205
rect 23845 38196 23857 38199
rect 22066 38168 23857 38196
rect 20349 38159 20407 38165
rect 23845 38165 23857 38168
rect 23891 38196 23903 38199
rect 24670 38196 24676 38208
rect 23891 38168 24676 38196
rect 23891 38165 23903 38168
rect 23845 38159 23903 38165
rect 24670 38156 24676 38168
rect 24728 38156 24734 38208
rect 25225 38199 25283 38205
rect 25225 38165 25237 38199
rect 25271 38196 25283 38199
rect 25314 38196 25320 38208
rect 25271 38168 25320 38196
rect 25271 38165 25283 38168
rect 25225 38159 25283 38165
rect 25314 38156 25320 38168
rect 25372 38156 25378 38208
rect 26326 38156 26332 38208
rect 26384 38196 26390 38208
rect 27065 38199 27123 38205
rect 27065 38196 27077 38199
rect 26384 38168 27077 38196
rect 26384 38156 26390 38168
rect 27065 38165 27077 38168
rect 27111 38165 27123 38199
rect 27065 38159 27123 38165
rect 31573 38199 31631 38205
rect 31573 38165 31585 38199
rect 31619 38196 31631 38199
rect 31754 38196 31760 38208
rect 31619 38168 31760 38196
rect 31619 38165 31631 38168
rect 31573 38159 31631 38165
rect 31754 38156 31760 38168
rect 31812 38156 31818 38208
rect 33502 38156 33508 38208
rect 33560 38196 33566 38208
rect 34057 38199 34115 38205
rect 34057 38196 34069 38199
rect 33560 38168 34069 38196
rect 33560 38156 33566 38168
rect 34057 38165 34069 38168
rect 34103 38165 34115 38199
rect 34057 38159 34115 38165
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 3050 37992 3056 38004
rect 3049 37952 3056 37992
rect 3108 37952 3114 38004
rect 3142 37952 3148 38004
rect 3200 37992 3206 38004
rect 4617 37995 4675 38001
rect 4617 37992 4629 37995
rect 3200 37964 4629 37992
rect 3200 37952 3206 37964
rect 4617 37961 4629 37964
rect 4663 37961 4675 37995
rect 4617 37955 4675 37961
rect 11698 37952 11704 38004
rect 11756 37992 11762 38004
rect 14369 37995 14427 38001
rect 11756 37964 11836 37992
rect 11756 37952 11762 37964
rect 3049 37871 3077 37952
rect 4157 37927 4215 37933
rect 4157 37893 4169 37927
rect 4203 37924 4215 37927
rect 4706 37924 4712 37936
rect 4203 37896 4712 37924
rect 4203 37893 4215 37896
rect 4157 37887 4215 37893
rect 4706 37884 4712 37896
rect 4764 37924 4770 37936
rect 11808 37933 11836 37964
rect 14369 37961 14381 37995
rect 14415 37992 14427 37995
rect 17586 37992 17592 38004
rect 14415 37964 17592 37992
rect 14415 37961 14427 37964
rect 14369 37955 14427 37961
rect 17586 37952 17592 37964
rect 17644 37952 17650 38004
rect 17770 37952 17776 38004
rect 17828 37992 17834 38004
rect 20346 37992 20352 38004
rect 17828 37964 20352 37992
rect 17828 37952 17834 37964
rect 20346 37952 20352 37964
rect 20404 37952 20410 38004
rect 25406 37952 25412 38004
rect 25464 37992 25470 38004
rect 26053 37995 26111 38001
rect 26053 37992 26065 37995
rect 25464 37964 26065 37992
rect 25464 37952 25470 37964
rect 26053 37961 26065 37964
rect 26099 37961 26111 37995
rect 26053 37955 26111 37961
rect 29178 37952 29184 38004
rect 29236 37952 29242 38004
rect 31110 37992 31116 38004
rect 31071 37964 31116 37992
rect 31110 37952 31116 37964
rect 31168 37952 31174 38004
rect 32766 37992 32772 38004
rect 31726 37964 32772 37992
rect 4985 37927 5043 37933
rect 4985 37924 4997 37927
rect 4764 37896 4997 37924
rect 4764 37884 4770 37896
rect 4985 37893 4997 37896
rect 5031 37893 5043 37927
rect 4985 37887 5043 37893
rect 11793 37927 11851 37933
rect 11793 37893 11805 37927
rect 11839 37893 11851 37927
rect 11793 37887 11851 37893
rect 13354 37884 13360 37936
rect 13412 37924 13418 37936
rect 13722 37924 13728 37936
rect 13412 37896 13728 37924
rect 13412 37884 13418 37896
rect 13722 37884 13728 37896
rect 13780 37924 13786 37936
rect 14001 37927 14059 37933
rect 14001 37924 14013 37927
rect 13780 37896 14013 37924
rect 13780 37884 13786 37896
rect 14001 37893 14013 37896
rect 14047 37893 14059 37927
rect 14001 37887 14059 37893
rect 14093 37927 14151 37933
rect 14093 37893 14105 37927
rect 14139 37924 14151 37927
rect 16758 37924 16764 37936
rect 14139 37896 16764 37924
rect 14139 37893 14151 37896
rect 14093 37887 14151 37893
rect 16758 37884 16764 37896
rect 16816 37884 16822 37936
rect 19426 37884 19432 37936
rect 19484 37924 19490 37936
rect 21085 37927 21143 37933
rect 21085 37924 21097 37927
rect 19484 37896 21097 37924
rect 19484 37884 19490 37896
rect 2774 37816 2780 37868
rect 2832 37856 2838 37868
rect 3034 37865 3092 37871
rect 2915 37859 2973 37865
rect 2915 37856 2927 37859
rect 2832 37828 2927 37856
rect 2832 37816 2838 37828
rect 2915 37825 2927 37828
rect 2961 37825 2973 37859
rect 3034 37831 3046 37865
rect 3080 37831 3092 37865
rect 3034 37825 3092 37831
rect 3150 37859 3208 37865
rect 3150 37825 3162 37859
rect 3196 37825 3208 37859
rect 3326 37856 3332 37868
rect 3287 37828 3332 37856
rect 2915 37819 2973 37825
rect 3150 37819 3208 37825
rect 3160 37788 3188 37819
rect 3326 37816 3332 37828
rect 3384 37816 3390 37868
rect 3418 37816 3424 37868
rect 3476 37856 3482 37868
rect 3973 37859 4031 37865
rect 3973 37856 3985 37859
rect 3476 37828 3985 37856
rect 3476 37816 3482 37828
rect 3973 37825 3985 37828
rect 4019 37825 4031 37859
rect 3973 37819 4031 37825
rect 4801 37859 4859 37865
rect 4801 37825 4813 37859
rect 4847 37856 4859 37859
rect 5074 37856 5080 37868
rect 4847 37828 5080 37856
rect 4847 37825 4859 37828
rect 4801 37819 4859 37825
rect 5074 37816 5080 37828
rect 5132 37816 5138 37868
rect 9306 37816 9312 37868
rect 9364 37856 9370 37868
rect 11517 37859 11575 37865
rect 11517 37856 11529 37859
rect 9364 37828 11529 37856
rect 9364 37816 9370 37828
rect 11517 37825 11529 37828
rect 11563 37825 11575 37859
rect 11698 37856 11704 37868
rect 11659 37828 11704 37856
rect 11517 37819 11575 37825
rect 11698 37816 11704 37828
rect 11756 37816 11762 37868
rect 11885 37859 11943 37865
rect 11885 37825 11897 37859
rect 11931 37856 11943 37859
rect 12250 37856 12256 37868
rect 11931 37828 12256 37856
rect 11931 37825 11943 37828
rect 11885 37819 11943 37825
rect 12250 37816 12256 37828
rect 12308 37816 12314 37868
rect 13817 37859 13875 37865
rect 13817 37856 13829 37859
rect 12406 37828 13829 37856
rect 3789 37791 3847 37797
rect 3789 37788 3801 37791
rect 3160 37760 3801 37788
rect 3789 37757 3801 37760
rect 3835 37757 3847 37791
rect 3789 37751 3847 37757
rect 10502 37748 10508 37800
rect 10560 37788 10566 37800
rect 12406 37788 12434 37828
rect 13817 37825 13829 37828
rect 13863 37825 13875 37859
rect 13817 37819 13875 37825
rect 14185 37859 14243 37865
rect 14185 37825 14197 37859
rect 14231 37825 14243 37859
rect 18138 37856 18144 37868
rect 18099 37828 18144 37856
rect 14185 37819 14243 37825
rect 10560 37760 12434 37788
rect 10560 37748 10566 37760
rect 12250 37680 12256 37732
rect 12308 37720 12314 37732
rect 13630 37720 13636 37732
rect 12308 37692 13636 37720
rect 12308 37680 12314 37692
rect 13630 37680 13636 37692
rect 13688 37720 13694 37732
rect 14200 37720 14228 37819
rect 18138 37816 18144 37828
rect 18196 37816 18202 37868
rect 18230 37816 18236 37868
rect 18288 37856 18294 37868
rect 18397 37859 18455 37865
rect 18397 37856 18409 37859
rect 18288 37828 18409 37856
rect 18288 37816 18294 37828
rect 18397 37825 18409 37828
rect 18443 37825 18455 37859
rect 18397 37819 18455 37825
rect 19150 37816 19156 37868
rect 19208 37856 19214 37868
rect 19702 37856 19708 37868
rect 19208 37828 19708 37856
rect 19208 37816 19214 37828
rect 19702 37816 19708 37828
rect 19760 37816 19766 37868
rect 19981 37859 20039 37865
rect 19981 37825 19993 37859
rect 20027 37825 20039 37859
rect 20162 37856 20168 37868
rect 20123 37828 20168 37856
rect 19981 37819 20039 37825
rect 19996 37788 20024 37819
rect 20162 37816 20168 37828
rect 20220 37816 20226 37868
rect 20364 37865 20392 37896
rect 21085 37893 21097 37896
rect 21131 37924 21143 37927
rect 23658 37924 23664 37936
rect 21131 37896 23664 37924
rect 21131 37893 21143 37896
rect 21085 37887 21143 37893
rect 23658 37884 23664 37896
rect 23716 37884 23722 37936
rect 25038 37884 25044 37936
rect 25096 37924 25102 37936
rect 25682 37924 25688 37936
rect 25096 37896 25688 37924
rect 25096 37884 25102 37896
rect 20257 37859 20315 37865
rect 20257 37825 20269 37859
rect 20303 37825 20315 37859
rect 20257 37819 20315 37825
rect 20349 37859 20407 37865
rect 20349 37825 20361 37859
rect 20395 37825 20407 37859
rect 20349 37819 20407 37825
rect 20272 37788 20300 37819
rect 25314 37816 25320 37868
rect 25372 37865 25378 37868
rect 25608 37865 25636 37896
rect 25682 37884 25688 37896
rect 25740 37884 25746 37936
rect 26142 37884 26148 37936
rect 26200 37924 26206 37936
rect 26421 37927 26479 37933
rect 26421 37924 26433 37927
rect 26200 37896 26433 37924
rect 26200 37884 26206 37896
rect 26421 37893 26433 37896
rect 26467 37893 26479 37927
rect 29196 37924 29224 37952
rect 31481 37927 31539 37933
rect 31481 37924 31493 37927
rect 29196 37896 31493 37924
rect 26421 37887 26479 37893
rect 31481 37893 31493 37896
rect 31527 37924 31539 37927
rect 31726 37924 31754 37964
rect 32766 37952 32772 37964
rect 32824 37952 32830 38004
rect 33042 37992 33048 38004
rect 33003 37964 33048 37992
rect 33042 37952 33048 37964
rect 33100 37952 33106 38004
rect 31527 37896 31754 37924
rect 31527 37893 31539 37896
rect 31481 37887 31539 37893
rect 25372 37856 25384 37865
rect 25593 37859 25651 37865
rect 25372 37828 25417 37856
rect 25372 37819 25384 37828
rect 25593 37825 25605 37859
rect 25639 37825 25651 37859
rect 25593 37819 25651 37825
rect 26237 37859 26295 37865
rect 26237 37825 26249 37859
rect 26283 37856 26295 37859
rect 26326 37856 26332 37868
rect 26283 37828 26332 37856
rect 26283 37825 26295 37828
rect 26237 37819 26295 37825
rect 25372 37816 25378 37819
rect 26326 37816 26332 37828
rect 26384 37816 26390 37868
rect 29178 37816 29184 37868
rect 29236 37856 29242 37868
rect 29345 37859 29403 37865
rect 29345 37856 29357 37859
rect 29236 37828 29357 37856
rect 29236 37816 29242 37828
rect 29345 37825 29357 37828
rect 29391 37825 29403 37859
rect 31294 37856 31300 37868
rect 31255 37828 31300 37856
rect 29345 37819 29403 37825
rect 31294 37816 31300 37828
rect 31352 37816 31358 37868
rect 31570 37816 31576 37868
rect 31628 37856 31634 37868
rect 32401 37859 32459 37865
rect 32401 37856 32413 37859
rect 31628 37828 32413 37856
rect 31628 37816 31634 37828
rect 32401 37825 32413 37828
rect 32447 37825 32459 37859
rect 32582 37856 32588 37868
rect 32543 37828 32588 37856
rect 32401 37819 32459 37825
rect 32582 37816 32588 37828
rect 32640 37816 32646 37868
rect 32677 37859 32735 37865
rect 32677 37825 32689 37859
rect 32723 37825 32735 37859
rect 32677 37819 32735 37825
rect 32769 37859 32827 37865
rect 32769 37825 32781 37859
rect 32815 37856 32827 37859
rect 33042 37856 33048 37868
rect 32815 37828 33048 37856
rect 32815 37825 32827 37828
rect 32769 37819 32827 37825
rect 19996 37760 20116 37788
rect 13688 37692 14228 37720
rect 13688 37680 13694 37692
rect 20088 37664 20116 37760
rect 20180 37760 20300 37788
rect 20180 37732 20208 37760
rect 20622 37748 20628 37800
rect 20680 37788 20686 37800
rect 22186 37788 22192 37800
rect 20680 37760 22192 37788
rect 20680 37748 20686 37760
rect 22186 37748 22192 37760
rect 22244 37748 22250 37800
rect 27430 37748 27436 37800
rect 27488 37788 27494 37800
rect 29086 37788 29092 37800
rect 27488 37760 29092 37788
rect 27488 37748 27494 37760
rect 29086 37748 29092 37760
rect 29144 37748 29150 37800
rect 32692 37788 32720 37819
rect 33042 37816 33048 37828
rect 33100 37816 33106 37868
rect 33778 37788 33784 37800
rect 32692 37760 33784 37788
rect 33778 37748 33784 37760
rect 33836 37748 33842 37800
rect 20162 37680 20168 37732
rect 20220 37680 20226 37732
rect 2682 37652 2688 37664
rect 2643 37624 2688 37652
rect 2682 37612 2688 37624
rect 2740 37612 2746 37664
rect 6730 37612 6736 37664
rect 6788 37652 6794 37664
rect 7193 37655 7251 37661
rect 7193 37652 7205 37655
rect 6788 37624 7205 37652
rect 6788 37612 6794 37624
rect 7193 37621 7205 37624
rect 7239 37652 7251 37655
rect 11330 37652 11336 37664
rect 7239 37624 11336 37652
rect 7239 37621 7251 37624
rect 7193 37615 7251 37621
rect 11330 37612 11336 37624
rect 11388 37612 11394 37664
rect 12069 37655 12127 37661
rect 12069 37621 12081 37655
rect 12115 37652 12127 37655
rect 13722 37652 13728 37664
rect 12115 37624 13728 37652
rect 12115 37621 12127 37624
rect 12069 37615 12127 37621
rect 13722 37612 13728 37624
rect 13780 37612 13786 37664
rect 17770 37612 17776 37664
rect 17828 37652 17834 37664
rect 19334 37652 19340 37664
rect 17828 37624 19340 37652
rect 17828 37612 17834 37624
rect 19334 37612 19340 37624
rect 19392 37652 19398 37664
rect 19521 37655 19579 37661
rect 19521 37652 19533 37655
rect 19392 37624 19533 37652
rect 19392 37612 19398 37624
rect 19521 37621 19533 37624
rect 19567 37621 19579 37655
rect 19521 37615 19579 37621
rect 20070 37612 20076 37664
rect 20128 37652 20134 37664
rect 20438 37652 20444 37664
rect 20128 37624 20444 37652
rect 20128 37612 20134 37624
rect 20438 37612 20444 37624
rect 20496 37612 20502 37664
rect 20625 37655 20683 37661
rect 20625 37621 20637 37655
rect 20671 37652 20683 37655
rect 20990 37652 20996 37664
rect 20671 37624 20996 37652
rect 20671 37621 20683 37624
rect 20625 37615 20683 37621
rect 20990 37612 20996 37624
rect 21048 37612 21054 37664
rect 24210 37652 24216 37664
rect 24171 37624 24216 37652
rect 24210 37612 24216 37624
rect 24268 37612 24274 37664
rect 27338 37652 27344 37664
rect 27299 37624 27344 37652
rect 27338 37612 27344 37624
rect 27396 37612 27402 37664
rect 30374 37612 30380 37664
rect 30432 37652 30438 37664
rect 30469 37655 30527 37661
rect 30469 37652 30481 37655
rect 30432 37624 30481 37652
rect 30432 37612 30438 37624
rect 30469 37621 30481 37624
rect 30515 37621 30527 37655
rect 30469 37615 30527 37621
rect 33042 37612 33048 37664
rect 33100 37652 33106 37664
rect 33505 37655 33563 37661
rect 33505 37652 33517 37655
rect 33100 37624 33517 37652
rect 33100 37612 33106 37624
rect 33505 37621 33517 37624
rect 33551 37621 33563 37655
rect 33505 37615 33563 37621
rect 34149 37655 34207 37661
rect 34149 37621 34161 37655
rect 34195 37652 34207 37655
rect 34330 37652 34336 37664
rect 34195 37624 34336 37652
rect 34195 37621 34207 37624
rect 34149 37615 34207 37621
rect 34330 37612 34336 37624
rect 34388 37612 34394 37664
rect 58158 37652 58164 37664
rect 58119 37624 58164 37652
rect 58158 37612 58164 37624
rect 58216 37612 58222 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 2774 37408 2780 37460
rect 2832 37448 2838 37460
rect 3789 37451 3847 37457
rect 3789 37448 3801 37451
rect 2832 37420 3801 37448
rect 2832 37408 2838 37420
rect 3789 37417 3801 37420
rect 3835 37448 3847 37451
rect 4062 37448 4068 37460
rect 3835 37420 4068 37448
rect 3835 37417 3847 37420
rect 3789 37411 3847 37417
rect 4062 37408 4068 37420
rect 4120 37408 4126 37460
rect 12342 37408 12348 37460
rect 12400 37448 12406 37460
rect 17402 37448 17408 37460
rect 12400 37420 17408 37448
rect 12400 37408 12406 37420
rect 17402 37408 17408 37420
rect 17460 37408 17466 37460
rect 18049 37451 18107 37457
rect 18049 37417 18061 37451
rect 18095 37448 18107 37451
rect 18230 37448 18236 37460
rect 18095 37420 18236 37448
rect 18095 37417 18107 37420
rect 18049 37411 18107 37417
rect 18230 37408 18236 37420
rect 18288 37408 18294 37460
rect 18506 37448 18512 37460
rect 18467 37420 18512 37448
rect 18506 37408 18512 37420
rect 18564 37408 18570 37460
rect 20441 37451 20499 37457
rect 20441 37417 20453 37451
rect 20487 37448 20499 37451
rect 20530 37448 20536 37460
rect 20487 37420 20536 37448
rect 20487 37417 20499 37420
rect 20441 37411 20499 37417
rect 16669 37383 16727 37389
rect 16669 37349 16681 37383
rect 16715 37380 16727 37383
rect 16850 37380 16856 37392
rect 16715 37352 16856 37380
rect 16715 37349 16727 37352
rect 16669 37343 16727 37349
rect 16850 37340 16856 37352
rect 16908 37380 16914 37392
rect 17678 37380 17684 37392
rect 16908 37352 17684 37380
rect 16908 37340 16914 37352
rect 17678 37340 17684 37352
rect 17736 37340 17742 37392
rect 1854 37312 1860 37324
rect 1815 37284 1860 37312
rect 1854 37272 1860 37284
rect 1912 37272 1918 37324
rect 14642 37272 14648 37324
rect 14700 37312 14706 37324
rect 14737 37315 14795 37321
rect 14737 37312 14749 37315
rect 14700 37284 14749 37312
rect 14700 37272 14706 37284
rect 14737 37281 14749 37284
rect 14783 37281 14795 37315
rect 20456 37312 20484 37411
rect 20530 37408 20536 37420
rect 20588 37408 20594 37460
rect 24673 37451 24731 37457
rect 24673 37417 24685 37451
rect 24719 37448 24731 37451
rect 24762 37448 24768 37460
rect 24719 37420 24768 37448
rect 24719 37417 24731 37420
rect 24673 37411 24731 37417
rect 24762 37408 24768 37420
rect 24820 37408 24826 37460
rect 30469 37451 30527 37457
rect 30469 37417 30481 37451
rect 30515 37448 30527 37451
rect 31478 37448 31484 37460
rect 30515 37420 31484 37448
rect 30515 37417 30527 37420
rect 30469 37411 30527 37417
rect 31478 37408 31484 37420
rect 31536 37408 31542 37460
rect 32582 37408 32588 37460
rect 32640 37448 32646 37460
rect 33045 37451 33103 37457
rect 33045 37448 33057 37451
rect 32640 37420 33057 37448
rect 32640 37408 32646 37420
rect 33045 37417 33057 37420
rect 33091 37417 33103 37451
rect 33045 37411 33103 37417
rect 31496 37380 31524 37408
rect 31496 37352 31754 37380
rect 14737 37275 14795 37281
rect 17328 37284 17724 37312
rect 2124 37247 2182 37253
rect 2124 37213 2136 37247
rect 2170 37244 2182 37247
rect 2682 37244 2688 37256
rect 2170 37216 2688 37244
rect 2170 37213 2182 37216
rect 2124 37207 2182 37213
rect 2682 37204 2688 37216
rect 2740 37204 2746 37256
rect 5997 37247 6055 37253
rect 5997 37213 6009 37247
rect 6043 37244 6055 37247
rect 6086 37244 6092 37256
rect 6043 37216 6092 37244
rect 6043 37213 6055 37216
rect 5997 37207 6055 37213
rect 6086 37204 6092 37216
rect 6144 37204 6150 37256
rect 7837 37247 7895 37253
rect 7837 37244 7849 37247
rect 7392 37216 7849 37244
rect 6264 37179 6322 37185
rect 6264 37145 6276 37179
rect 6310 37176 6322 37179
rect 7098 37176 7104 37188
rect 6310 37148 7104 37176
rect 6310 37145 6322 37148
rect 6264 37139 6322 37145
rect 7098 37136 7104 37148
rect 7156 37136 7162 37188
rect 3237 37111 3295 37117
rect 3237 37077 3249 37111
rect 3283 37108 3295 37111
rect 3326 37108 3332 37120
rect 3283 37080 3332 37108
rect 3283 37077 3295 37080
rect 3237 37071 3295 37077
rect 3326 37068 3332 37080
rect 3384 37068 3390 37120
rect 7392 37117 7420 37216
rect 7837 37213 7849 37216
rect 7883 37213 7895 37247
rect 8110 37244 8116 37256
rect 8071 37216 8116 37244
rect 7837 37207 7895 37213
rect 8110 37204 8116 37216
rect 8168 37204 8174 37256
rect 8202 37204 8208 37256
rect 8260 37244 8266 37256
rect 11698 37244 11704 37256
rect 8260 37216 8305 37244
rect 11164 37216 11704 37244
rect 8260 37204 8266 37216
rect 8018 37176 8024 37188
rect 7979 37148 8024 37176
rect 8018 37136 8024 37148
rect 8076 37176 8082 37188
rect 11164 37176 11192 37216
rect 11698 37204 11704 37216
rect 11756 37204 11762 37256
rect 15289 37247 15347 37253
rect 15289 37244 15301 37247
rect 13280 37216 15301 37244
rect 8076 37148 11192 37176
rect 8076 37136 8082 37148
rect 11330 37136 11336 37188
rect 11388 37176 11394 37188
rect 11793 37179 11851 37185
rect 11793 37176 11805 37179
rect 11388 37148 11805 37176
rect 11388 37136 11394 37148
rect 11793 37145 11805 37148
rect 11839 37176 11851 37179
rect 12342 37176 12348 37188
rect 11839 37148 12348 37176
rect 11839 37145 11851 37148
rect 11793 37139 11851 37145
rect 12342 37136 12348 37148
rect 12400 37136 12406 37188
rect 13280 37120 13308 37216
rect 15289 37213 15301 37216
rect 15335 37213 15347 37247
rect 17328 37244 17356 37284
rect 15289 37207 15347 37213
rect 15488 37216 17356 37244
rect 14366 37176 14372 37188
rect 14327 37148 14372 37176
rect 14366 37136 14372 37148
rect 14424 37136 14430 37188
rect 14550 37176 14556 37188
rect 14511 37148 14556 37176
rect 14550 37136 14556 37148
rect 14608 37136 14614 37188
rect 14660 37148 14872 37176
rect 7377 37111 7435 37117
rect 7377 37077 7389 37111
rect 7423 37108 7435 37111
rect 7558 37108 7564 37120
rect 7423 37080 7564 37108
rect 7423 37077 7435 37080
rect 7377 37071 7435 37077
rect 7558 37068 7564 37080
rect 7616 37068 7622 37120
rect 8389 37111 8447 37117
rect 8389 37077 8401 37111
rect 8435 37108 8447 37111
rect 8938 37108 8944 37120
rect 8435 37080 8944 37108
rect 8435 37077 8447 37080
rect 8389 37071 8447 37077
rect 8938 37068 8944 37080
rect 8996 37068 9002 37120
rect 13262 37108 13268 37120
rect 13223 37080 13268 37108
rect 13262 37068 13268 37080
rect 13320 37068 13326 37120
rect 13722 37068 13728 37120
rect 13780 37108 13786 37120
rect 14660 37108 14688 37148
rect 13780 37080 14688 37108
rect 14844 37108 14872 37148
rect 15194 37136 15200 37188
rect 15252 37176 15258 37188
rect 15488 37176 15516 37216
rect 17402 37204 17408 37256
rect 17460 37244 17466 37256
rect 17586 37244 17592 37256
rect 17460 37216 17505 37244
rect 17547 37216 17592 37244
rect 17460 37204 17466 37216
rect 17586 37204 17592 37216
rect 17644 37204 17650 37256
rect 17696 37253 17724 37284
rect 19628 37284 20484 37312
rect 31481 37315 31539 37321
rect 17681 37247 17739 37253
rect 17681 37213 17693 37247
rect 17727 37213 17739 37247
rect 17681 37207 17739 37213
rect 17773 37247 17831 37253
rect 17773 37213 17785 37247
rect 17819 37244 17831 37247
rect 18506 37244 18512 37256
rect 17819 37216 18512 37244
rect 17819 37213 17831 37216
rect 17773 37207 17831 37213
rect 18506 37204 18512 37216
rect 18564 37204 18570 37256
rect 19245 37247 19303 37253
rect 19245 37213 19257 37247
rect 19291 37213 19303 37247
rect 19245 37207 19303 37213
rect 15562 37185 15568 37188
rect 15252 37148 15516 37176
rect 15252 37136 15258 37148
rect 15556 37139 15568 37185
rect 15620 37176 15626 37188
rect 19260 37176 19288 37207
rect 19334 37204 19340 37256
rect 19392 37244 19398 37256
rect 19628 37253 19656 37284
rect 31481 37281 31493 37315
rect 31527 37312 31539 37315
rect 31570 37312 31576 37324
rect 31527 37284 31576 37312
rect 31527 37281 31539 37284
rect 31481 37275 31539 37281
rect 31570 37272 31576 37284
rect 31628 37272 31634 37324
rect 31726 37321 31754 37352
rect 31711 37315 31769 37321
rect 31711 37281 31723 37315
rect 31757 37281 31769 37315
rect 31711 37275 31769 37281
rect 33318 37272 33324 37324
rect 33376 37312 33382 37324
rect 34238 37312 34244 37324
rect 33376 37284 33548 37312
rect 33376 37272 33382 37284
rect 19613 37247 19671 37253
rect 19392 37216 19437 37244
rect 19392 37204 19398 37216
rect 19613 37213 19625 37247
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 19702 37204 19708 37256
rect 19760 37253 19766 37256
rect 19760 37244 19768 37253
rect 19760 37216 19805 37244
rect 19760 37207 19768 37216
rect 19760 37204 19766 37207
rect 20990 37204 20996 37256
rect 21048 37244 21054 37256
rect 21554 37247 21612 37253
rect 21554 37244 21566 37247
rect 21048 37216 21566 37244
rect 21048 37204 21054 37216
rect 21554 37213 21566 37216
rect 21600 37213 21612 37247
rect 21818 37244 21824 37256
rect 21779 37216 21824 37244
rect 21554 37207 21612 37213
rect 21818 37204 21824 37216
rect 21876 37204 21882 37256
rect 32677 37247 32735 37253
rect 32677 37213 32689 37247
rect 32723 37244 32735 37247
rect 33410 37244 33416 37256
rect 32723 37216 33416 37244
rect 32723 37213 32735 37216
rect 32677 37207 32735 37213
rect 33410 37204 33416 37216
rect 33468 37204 33474 37256
rect 33520 37253 33548 37284
rect 33796 37284 34244 37312
rect 33796 37256 33824 37284
rect 34238 37272 34244 37284
rect 34296 37272 34302 37324
rect 33505 37247 33563 37253
rect 33505 37213 33517 37247
rect 33551 37213 33563 37247
rect 33686 37244 33692 37256
rect 33647 37216 33692 37244
rect 33505 37207 33563 37213
rect 33686 37204 33692 37216
rect 33744 37204 33750 37256
rect 33778 37204 33784 37256
rect 33836 37244 33842 37256
rect 33919 37247 33977 37253
rect 33836 37216 33881 37244
rect 33836 37204 33842 37216
rect 33919 37213 33931 37247
rect 33965 37244 33977 37247
rect 34330 37244 34336 37256
rect 33965 37216 34336 37244
rect 33965 37213 33977 37216
rect 33919 37207 33977 37213
rect 34330 37204 34336 37216
rect 34388 37204 34394 37256
rect 36081 37247 36139 37253
rect 36081 37213 36093 37247
rect 36127 37244 36139 37247
rect 36722 37244 36728 37256
rect 36127 37216 36728 37244
rect 36127 37213 36139 37216
rect 36081 37207 36139 37213
rect 36722 37204 36728 37216
rect 36780 37204 36786 37256
rect 15620 37148 15656 37176
rect 15764 37148 19288 37176
rect 15562 37136 15568 37139
rect 15620 37136 15626 37148
rect 15764 37108 15792 37148
rect 19426 37136 19432 37188
rect 19484 37176 19490 37188
rect 19521 37179 19579 37185
rect 19521 37176 19533 37179
rect 19484 37148 19533 37176
rect 19484 37136 19490 37148
rect 19521 37145 19533 37148
rect 19567 37145 19579 37179
rect 19521 37139 19579 37145
rect 24210 37136 24216 37188
rect 24268 37176 24274 37188
rect 24857 37179 24915 37185
rect 24857 37176 24869 37179
rect 24268 37148 24869 37176
rect 24268 37136 24274 37148
rect 24857 37145 24869 37148
rect 24903 37145 24915 37179
rect 24857 37139 24915 37145
rect 24946 37136 24952 37188
rect 25004 37176 25010 37188
rect 25041 37179 25099 37185
rect 25041 37176 25053 37179
rect 25004 37148 25053 37176
rect 25004 37136 25010 37148
rect 25041 37145 25053 37148
rect 25087 37176 25099 37179
rect 26142 37176 26148 37188
rect 25087 37148 26148 37176
rect 25087 37145 25099 37148
rect 25041 37139 25099 37145
rect 26142 37136 26148 37148
rect 26200 37136 26206 37188
rect 32861 37179 32919 37185
rect 32861 37145 32873 37179
rect 32907 37176 32919 37179
rect 34149 37179 34207 37185
rect 32907 37148 33548 37176
rect 32907 37145 32919 37148
rect 32861 37139 32919 37145
rect 33520 37120 33548 37148
rect 34149 37145 34161 37179
rect 34195 37176 34207 37179
rect 35814 37179 35872 37185
rect 35814 37176 35826 37179
rect 34195 37148 35826 37176
rect 34195 37145 34207 37148
rect 34149 37139 34207 37145
rect 35814 37145 35826 37148
rect 35860 37145 35872 37179
rect 35814 37139 35872 37145
rect 14844 37080 15792 37108
rect 13780 37068 13786 37080
rect 16114 37068 16120 37120
rect 16172 37108 16178 37120
rect 17402 37108 17408 37120
rect 16172 37080 17408 37108
rect 16172 37068 16178 37080
rect 17402 37068 17408 37080
rect 17460 37068 17466 37120
rect 19150 37068 19156 37120
rect 19208 37108 19214 37120
rect 19702 37108 19708 37120
rect 19208 37080 19708 37108
rect 19208 37068 19214 37080
rect 19702 37068 19708 37080
rect 19760 37068 19766 37120
rect 19889 37111 19947 37117
rect 19889 37077 19901 37111
rect 19935 37108 19947 37111
rect 20898 37108 20904 37120
rect 19935 37080 20904 37108
rect 19935 37077 19947 37080
rect 19889 37071 19947 37077
rect 20898 37068 20904 37080
rect 20956 37068 20962 37120
rect 22830 37068 22836 37120
rect 22888 37108 22894 37120
rect 23385 37111 23443 37117
rect 23385 37108 23397 37111
rect 22888 37080 23397 37108
rect 22888 37068 22894 37080
rect 23385 37077 23397 37080
rect 23431 37077 23443 37111
rect 23385 37071 23443 37077
rect 33502 37068 33508 37120
rect 33560 37068 33566 37120
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 34701 37111 34759 37117
rect 34701 37108 34713 37111
rect 34572 37080 34713 37108
rect 34572 37068 34578 37080
rect 34701 37077 34713 37080
rect 34747 37077 34759 37111
rect 34701 37071 34759 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 8202 36904 8208 36916
rect 6748 36876 8208 36904
rect 6638 36836 6644 36848
rect 6599 36808 6644 36836
rect 6638 36796 6644 36808
rect 6696 36796 6702 36848
rect 5166 36728 5172 36780
rect 5224 36768 5230 36780
rect 6748 36777 6776 36876
rect 8202 36864 8208 36876
rect 8260 36904 8266 36916
rect 12250 36904 12256 36916
rect 8260 36876 12256 36904
rect 8260 36864 8266 36876
rect 12250 36864 12256 36876
rect 12308 36904 12314 36916
rect 12897 36907 12955 36913
rect 12897 36904 12909 36907
rect 12308 36876 12909 36904
rect 12308 36864 12314 36876
rect 12897 36873 12909 36876
rect 12943 36873 12955 36907
rect 12897 36867 12955 36873
rect 14366 36864 14372 36916
rect 14424 36904 14430 36916
rect 15473 36907 15531 36913
rect 14424 36876 15056 36904
rect 14424 36864 14430 36876
rect 7558 36836 7564 36848
rect 7519 36808 7564 36836
rect 7558 36796 7564 36808
rect 7616 36796 7622 36848
rect 11698 36796 11704 36848
rect 11756 36836 11762 36848
rect 12710 36836 12716 36848
rect 11756 36808 12716 36836
rect 11756 36796 11762 36808
rect 12710 36796 12716 36808
rect 12768 36836 12774 36848
rect 13354 36836 13360 36848
rect 12768 36808 13360 36836
rect 12768 36796 12774 36808
rect 13354 36796 13360 36808
rect 13412 36796 13418 36848
rect 15028 36836 15056 36876
rect 15473 36873 15485 36907
rect 15519 36904 15531 36907
rect 15562 36904 15568 36916
rect 15519 36876 15568 36904
rect 15519 36873 15531 36876
rect 15473 36867 15531 36873
rect 15562 36864 15568 36876
rect 15620 36864 15626 36916
rect 17586 36864 17592 36916
rect 17644 36904 17650 36916
rect 18049 36907 18107 36913
rect 18049 36904 18061 36907
rect 17644 36876 18061 36904
rect 17644 36864 17650 36876
rect 18049 36873 18061 36876
rect 18095 36873 18107 36907
rect 18049 36867 18107 36873
rect 19242 36864 19248 36916
rect 19300 36904 19306 36916
rect 19889 36907 19947 36913
rect 19889 36904 19901 36907
rect 19300 36876 19901 36904
rect 19300 36864 19306 36876
rect 19889 36873 19901 36876
rect 19935 36904 19947 36907
rect 20070 36904 20076 36916
rect 19935 36876 20076 36904
rect 19935 36873 19947 36876
rect 19889 36867 19947 36873
rect 20070 36864 20076 36876
rect 20128 36864 20134 36916
rect 16850 36836 16856 36848
rect 15028 36808 16252 36836
rect 16811 36808 16856 36836
rect 6365 36771 6423 36777
rect 6365 36768 6377 36771
rect 5224 36740 6377 36768
rect 5224 36728 5230 36740
rect 6365 36737 6377 36740
rect 6411 36737 6423 36771
rect 6365 36731 6423 36737
rect 6549 36771 6607 36777
rect 6549 36737 6561 36771
rect 6595 36737 6607 36771
rect 6549 36731 6607 36737
rect 6733 36771 6791 36777
rect 6733 36737 6745 36771
rect 6779 36737 6791 36771
rect 6733 36731 6791 36737
rect 6564 36700 6592 36731
rect 7282 36728 7288 36780
rect 7340 36768 7346 36780
rect 7377 36771 7435 36777
rect 7377 36768 7389 36771
rect 7340 36740 7389 36768
rect 7340 36728 7346 36740
rect 7377 36737 7389 36740
rect 7423 36737 7435 36771
rect 7377 36731 7435 36737
rect 10226 36728 10232 36780
rect 10284 36768 10290 36780
rect 10781 36771 10839 36777
rect 10781 36768 10793 36771
rect 10284 36740 10793 36768
rect 10284 36728 10290 36740
rect 10781 36737 10793 36740
rect 10827 36768 10839 36771
rect 12161 36771 12219 36777
rect 12161 36768 12173 36771
rect 10827 36740 12173 36768
rect 10827 36737 10839 36740
rect 10781 36731 10839 36737
rect 12161 36737 12173 36740
rect 12207 36737 12219 36771
rect 12161 36731 12219 36737
rect 12802 36728 12808 36780
rect 12860 36768 12866 36780
rect 12989 36771 13047 36777
rect 12989 36768 13001 36771
rect 12860 36740 13001 36768
rect 12860 36728 12866 36740
rect 12989 36737 13001 36740
rect 13035 36737 13047 36771
rect 12989 36731 13047 36737
rect 13808 36771 13866 36777
rect 13808 36737 13820 36771
rect 13854 36768 13866 36771
rect 14090 36768 14096 36780
rect 13854 36740 14096 36768
rect 13854 36737 13866 36740
rect 13808 36731 13866 36737
rect 14090 36728 14096 36740
rect 14148 36728 14154 36780
rect 15746 36768 15752 36780
rect 15707 36740 15752 36768
rect 15746 36728 15752 36740
rect 15804 36728 15810 36780
rect 15841 36771 15899 36777
rect 15841 36737 15853 36771
rect 15887 36737 15899 36771
rect 15841 36731 15899 36737
rect 15933 36771 15991 36777
rect 15933 36737 15945 36771
rect 15979 36737 15991 36771
rect 16114 36768 16120 36780
rect 16075 36740 16120 36768
rect 15933 36731 15991 36737
rect 8018 36700 8024 36712
rect 6564 36672 8024 36700
rect 8018 36660 8024 36672
rect 8076 36660 8082 36712
rect 9766 36660 9772 36712
rect 9824 36700 9830 36712
rect 10410 36700 10416 36712
rect 9824 36672 10416 36700
rect 9824 36660 9830 36672
rect 10410 36660 10416 36672
rect 10468 36700 10474 36712
rect 10505 36703 10563 36709
rect 10505 36700 10517 36703
rect 10468 36672 10517 36700
rect 10468 36660 10474 36672
rect 10505 36669 10517 36672
rect 10551 36669 10563 36703
rect 10505 36663 10563 36669
rect 13262 36660 13268 36712
rect 13320 36700 13326 36712
rect 13541 36703 13599 36709
rect 13541 36700 13553 36703
rect 13320 36672 13553 36700
rect 13320 36660 13326 36672
rect 13541 36669 13553 36672
rect 13587 36669 13599 36703
rect 13541 36663 13599 36669
rect 15194 36660 15200 36712
rect 15252 36700 15258 36712
rect 15856 36700 15884 36731
rect 15252 36672 15884 36700
rect 15948 36700 15976 36731
rect 16114 36728 16120 36740
rect 16172 36728 16178 36780
rect 16224 36768 16252 36808
rect 16850 36796 16856 36808
rect 16908 36796 16914 36848
rect 17770 36796 17776 36848
rect 17828 36836 17834 36848
rect 17865 36839 17923 36845
rect 17865 36836 17877 36839
rect 17828 36808 17877 36836
rect 17828 36796 17834 36808
rect 17865 36805 17877 36808
rect 17911 36805 17923 36839
rect 17865 36799 17923 36805
rect 23017 36839 23075 36845
rect 23017 36805 23029 36839
rect 23063 36836 23075 36839
rect 24210 36836 24216 36848
rect 23063 36808 24216 36836
rect 23063 36805 23075 36808
rect 23017 36799 23075 36805
rect 24210 36796 24216 36808
rect 24268 36796 24274 36848
rect 17037 36771 17095 36777
rect 17037 36768 17049 36771
rect 16224 36740 17049 36768
rect 17037 36737 17049 36740
rect 17083 36768 17095 36771
rect 17678 36768 17684 36780
rect 17083 36740 17684 36768
rect 17083 36737 17095 36740
rect 17037 36731 17095 36737
rect 17678 36728 17684 36740
rect 17736 36728 17742 36780
rect 22830 36728 22836 36780
rect 22888 36768 22894 36780
rect 22925 36771 22983 36777
rect 22925 36768 22937 36771
rect 22888 36740 22937 36768
rect 22888 36728 22894 36740
rect 22925 36737 22937 36740
rect 22971 36737 22983 36771
rect 22925 36731 22983 36737
rect 23109 36771 23167 36777
rect 23109 36737 23121 36771
rect 23155 36737 23167 36771
rect 23290 36768 23296 36780
rect 23251 36740 23296 36768
rect 23109 36731 23167 36737
rect 16669 36703 16727 36709
rect 16669 36700 16681 36703
rect 15948 36672 16681 36700
rect 15252 36660 15258 36672
rect 16669 36669 16681 36672
rect 16715 36669 16727 36703
rect 23124 36700 23152 36731
rect 23290 36728 23296 36740
rect 23348 36728 23354 36780
rect 23753 36771 23811 36777
rect 23753 36737 23765 36771
rect 23799 36768 23811 36771
rect 25961 36771 26019 36777
rect 25961 36768 25973 36771
rect 23799 36740 25973 36768
rect 23799 36737 23811 36740
rect 23753 36731 23811 36737
rect 25961 36737 25973 36740
rect 26007 36768 26019 36771
rect 28994 36768 29000 36780
rect 26007 36740 29000 36768
rect 26007 36737 26019 36740
rect 25961 36731 26019 36737
rect 28994 36728 29000 36740
rect 29052 36728 29058 36780
rect 34241 36771 34299 36777
rect 34241 36737 34253 36771
rect 34287 36768 34299 36771
rect 34422 36768 34428 36780
rect 34287 36740 34428 36768
rect 34287 36737 34299 36740
rect 34241 36731 34299 36737
rect 34422 36728 34428 36740
rect 34480 36728 34486 36780
rect 35342 36728 35348 36780
rect 35400 36768 35406 36780
rect 36458 36771 36516 36777
rect 36458 36768 36470 36771
rect 35400 36740 36470 36768
rect 35400 36728 35406 36740
rect 36458 36737 36470 36740
rect 36504 36737 36516 36771
rect 36458 36731 36516 36737
rect 36722 36700 36728 36712
rect 16669 36663 16727 36669
rect 22388 36672 23152 36700
rect 36683 36672 36728 36700
rect 14550 36592 14556 36644
rect 14608 36632 14614 36644
rect 14921 36635 14979 36641
rect 14921 36632 14933 36635
rect 14608 36604 14933 36632
rect 14608 36592 14614 36604
rect 14921 36601 14933 36604
rect 14967 36632 14979 36635
rect 19334 36632 19340 36644
rect 14967 36604 19340 36632
rect 14967 36601 14979 36604
rect 14921 36595 14979 36601
rect 19334 36592 19340 36604
rect 19392 36592 19398 36644
rect 22388 36576 22416 36672
rect 36722 36660 36728 36672
rect 36780 36660 36786 36712
rect 6914 36564 6920 36576
rect 6875 36536 6920 36564
rect 6914 36524 6920 36536
rect 6972 36524 6978 36576
rect 7650 36524 7656 36576
rect 7708 36564 7714 36576
rect 7745 36567 7803 36573
rect 7745 36564 7757 36567
rect 7708 36536 7757 36564
rect 7708 36524 7714 36536
rect 7745 36533 7757 36536
rect 7791 36533 7803 36567
rect 7745 36527 7803 36533
rect 12253 36567 12311 36573
rect 12253 36533 12265 36567
rect 12299 36564 12311 36567
rect 12618 36564 12624 36576
rect 12299 36536 12624 36564
rect 12299 36533 12311 36536
rect 12253 36527 12311 36533
rect 12618 36524 12624 36536
rect 12676 36524 12682 36576
rect 22281 36567 22339 36573
rect 22281 36533 22293 36567
rect 22327 36564 22339 36567
rect 22370 36564 22376 36576
rect 22327 36536 22376 36564
rect 22327 36533 22339 36536
rect 22281 36527 22339 36533
rect 22370 36524 22376 36536
rect 22428 36524 22434 36576
rect 22741 36567 22799 36573
rect 22741 36533 22753 36567
rect 22787 36564 22799 36567
rect 22922 36564 22928 36576
rect 22787 36536 22928 36564
rect 22787 36533 22799 36536
rect 22741 36527 22799 36533
rect 22922 36524 22928 36536
rect 22980 36524 22986 36576
rect 25038 36564 25044 36576
rect 24999 36536 25044 36564
rect 25038 36524 25044 36536
rect 25096 36524 25102 36576
rect 27522 36524 27528 36576
rect 27580 36564 27586 36576
rect 27985 36567 28043 36573
rect 27985 36564 27997 36567
rect 27580 36536 27997 36564
rect 27580 36524 27586 36536
rect 27985 36533 27997 36536
rect 28031 36533 28043 36567
rect 27985 36527 28043 36533
rect 32953 36567 33011 36573
rect 32953 36533 32965 36567
rect 32999 36564 33011 36567
rect 33134 36564 33140 36576
rect 32999 36536 33140 36564
rect 32999 36533 33011 36536
rect 32953 36527 33011 36533
rect 33134 36524 33140 36536
rect 33192 36524 33198 36576
rect 34790 36564 34796 36576
rect 34751 36536 34796 36564
rect 34790 36524 34796 36536
rect 34848 36524 34854 36576
rect 35345 36567 35403 36573
rect 35345 36533 35357 36567
rect 35391 36564 35403 36567
rect 35434 36564 35440 36576
rect 35391 36536 35440 36564
rect 35391 36533 35403 36536
rect 35345 36527 35403 36533
rect 35434 36524 35440 36536
rect 35492 36524 35498 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 5166 36360 5172 36372
rect 5127 36332 5172 36360
rect 5166 36320 5172 36332
rect 5224 36320 5230 36372
rect 7098 36360 7104 36372
rect 7059 36332 7104 36360
rect 7098 36320 7104 36332
rect 7156 36320 7162 36372
rect 14090 36360 14096 36372
rect 14051 36332 14096 36360
rect 14090 36320 14096 36332
rect 14148 36320 14154 36372
rect 15746 36320 15752 36372
rect 15804 36360 15810 36372
rect 16298 36360 16304 36372
rect 15804 36332 16304 36360
rect 15804 36320 15810 36332
rect 16298 36320 16304 36332
rect 16356 36320 16362 36372
rect 28994 36320 29000 36372
rect 29052 36360 29058 36372
rect 29730 36360 29736 36372
rect 29052 36332 29736 36360
rect 29052 36320 29058 36332
rect 29730 36320 29736 36332
rect 29788 36360 29794 36372
rect 29788 36332 32444 36360
rect 29788 36320 29794 36332
rect 8110 36292 8116 36304
rect 7481 36264 8116 36292
rect 1854 36184 1860 36236
rect 1912 36224 1918 36236
rect 3789 36227 3847 36233
rect 3789 36224 3801 36227
rect 1912 36196 3801 36224
rect 1912 36184 1918 36196
rect 3789 36193 3801 36196
rect 3835 36193 3847 36227
rect 3789 36187 3847 36193
rect 7374 36156 7380 36168
rect 7335 36128 7380 36156
rect 7374 36116 7380 36128
rect 7432 36116 7438 36168
rect 7481 36165 7509 36264
rect 8110 36252 8116 36264
rect 8168 36252 8174 36304
rect 27890 36292 27896 36304
rect 27803 36264 27896 36292
rect 27890 36252 27896 36264
rect 27948 36292 27954 36304
rect 28718 36292 28724 36304
rect 27948 36264 28724 36292
rect 27948 36252 27954 36264
rect 28718 36252 28724 36264
rect 28776 36252 28782 36304
rect 9766 36224 9772 36236
rect 7760 36196 9772 36224
rect 7466 36159 7524 36165
rect 7466 36125 7478 36159
rect 7512 36125 7524 36159
rect 7466 36119 7524 36125
rect 7561 36156 7619 36162
rect 7650 36156 7656 36168
rect 7561 36122 7573 36156
rect 7607 36128 7656 36156
rect 7607 36122 7619 36128
rect 7561 36116 7619 36122
rect 7650 36116 7656 36128
rect 7708 36116 7714 36168
rect 7760 36165 7788 36196
rect 9766 36184 9772 36196
rect 9824 36184 9830 36236
rect 12710 36224 12716 36236
rect 12671 36196 12716 36224
rect 12710 36184 12716 36196
rect 12768 36184 12774 36236
rect 15197 36227 15255 36233
rect 15197 36224 15209 36227
rect 14384 36196 15209 36224
rect 7745 36159 7803 36165
rect 7745 36125 7757 36159
rect 7791 36125 7803 36159
rect 7745 36119 7803 36125
rect 8202 36116 8208 36168
rect 8260 36156 8266 36168
rect 9401 36159 9459 36165
rect 9401 36156 9413 36159
rect 8260 36128 9413 36156
rect 8260 36116 8266 36128
rect 9401 36125 9413 36128
rect 9447 36125 9459 36159
rect 9401 36119 9459 36125
rect 10045 36159 10103 36165
rect 10045 36125 10057 36159
rect 10091 36156 10103 36159
rect 10091 36128 11008 36156
rect 10091 36125 10103 36128
rect 10045 36119 10103 36125
rect 4056 36091 4114 36097
rect 4056 36057 4068 36091
rect 4102 36088 4114 36091
rect 4706 36088 4712 36100
rect 4102 36060 4712 36088
rect 4102 36057 4114 36060
rect 4056 36051 4114 36057
rect 4706 36048 4712 36060
rect 4764 36048 4770 36100
rect 7392 36088 7420 36116
rect 10428 36100 10456 36128
rect 10318 36097 10324 36100
rect 8297 36091 8355 36097
rect 8297 36088 8309 36091
rect 7392 36060 8309 36088
rect 8297 36057 8309 36060
rect 8343 36057 8355 36091
rect 10312 36088 10324 36097
rect 10279 36060 10324 36088
rect 8297 36051 8355 36057
rect 10312 36051 10324 36060
rect 10318 36048 10324 36051
rect 10376 36048 10382 36100
rect 10410 36048 10416 36100
rect 10468 36048 10474 36100
rect 10980 36088 11008 36128
rect 12434 36116 12440 36168
rect 12492 36156 12498 36168
rect 12492 36128 12537 36156
rect 12492 36116 12498 36128
rect 14274 36116 14280 36168
rect 14332 36156 14338 36168
rect 14384 36165 14412 36196
rect 15197 36193 15209 36196
rect 15243 36224 15255 36227
rect 21634 36224 21640 36236
rect 15243 36196 21640 36224
rect 15243 36193 15255 36196
rect 15197 36187 15255 36193
rect 21634 36184 21640 36196
rect 21692 36224 21698 36236
rect 22094 36224 22100 36236
rect 21692 36196 22100 36224
rect 21692 36184 21698 36196
rect 22094 36184 22100 36196
rect 22152 36184 22158 36236
rect 24762 36224 24768 36236
rect 22296 36196 24768 36224
rect 14369 36159 14427 36165
rect 14369 36156 14381 36159
rect 14332 36128 14381 36156
rect 14332 36116 14338 36128
rect 14369 36125 14381 36128
rect 14415 36125 14427 36159
rect 14369 36119 14427 36125
rect 14461 36159 14519 36165
rect 14461 36125 14473 36159
rect 14507 36125 14519 36159
rect 14461 36119 14519 36125
rect 14553 36159 14611 36165
rect 14553 36125 14565 36159
rect 14599 36156 14611 36159
rect 14642 36156 14648 36168
rect 14599 36128 14648 36156
rect 14599 36125 14611 36128
rect 14553 36119 14611 36125
rect 13262 36088 13268 36100
rect 10980 36060 13268 36088
rect 13262 36048 13268 36060
rect 13320 36048 13326 36100
rect 14476 36088 14504 36119
rect 14642 36116 14648 36128
rect 14700 36116 14706 36168
rect 14734 36116 14740 36168
rect 14792 36156 14798 36168
rect 22186 36156 22192 36168
rect 14792 36128 14837 36156
rect 22147 36128 22192 36156
rect 14792 36116 14798 36128
rect 22186 36116 22192 36128
rect 22244 36116 22250 36168
rect 22296 36165 22324 36196
rect 24762 36184 24768 36196
rect 24820 36184 24826 36236
rect 28442 36184 28448 36236
rect 28500 36224 28506 36236
rect 28997 36227 29055 36233
rect 28500 36196 28672 36224
rect 28500 36184 28506 36196
rect 22281 36159 22339 36165
rect 22281 36125 22293 36159
rect 22327 36125 22339 36159
rect 22554 36156 22560 36168
rect 22515 36128 22560 36156
rect 22281 36119 22339 36125
rect 22554 36116 22560 36128
rect 22612 36116 22618 36168
rect 22830 36116 22836 36168
rect 22888 36156 22894 36168
rect 24397 36159 24455 36165
rect 24397 36156 24409 36159
rect 22888 36128 24409 36156
rect 22888 36116 22894 36128
rect 24397 36125 24409 36128
rect 24443 36125 24455 36159
rect 27522 36156 27528 36168
rect 24397 36119 24455 36125
rect 27080 36128 27528 36156
rect 15194 36088 15200 36100
rect 14476 36060 15200 36088
rect 15194 36048 15200 36060
rect 15252 36048 15258 36100
rect 22370 36088 22376 36100
rect 22283 36060 22376 36088
rect 22370 36048 22376 36060
rect 22428 36088 22434 36100
rect 22428 36060 23336 36088
rect 22428 36048 22434 36060
rect 23308 36032 23336 36060
rect 27080 36032 27108 36128
rect 27522 36116 27528 36128
rect 27580 36156 27586 36168
rect 28644 36165 28672 36196
rect 28997 36193 29009 36227
rect 29043 36224 29055 36227
rect 29178 36224 29184 36236
rect 29043 36196 29184 36224
rect 29043 36193 29055 36196
rect 28997 36187 29055 36193
rect 29178 36184 29184 36196
rect 29236 36184 29242 36236
rect 28353 36159 28411 36165
rect 28353 36156 28365 36159
rect 27580 36128 28365 36156
rect 27580 36116 27586 36128
rect 28353 36125 28365 36128
rect 28399 36125 28411 36159
rect 28537 36159 28595 36165
rect 28537 36156 28549 36159
rect 28353 36119 28411 36125
rect 28460 36128 28549 36156
rect 28460 36088 28488 36128
rect 28537 36125 28549 36128
rect 28583 36125 28595 36159
rect 28537 36119 28595 36125
rect 28629 36159 28687 36165
rect 28629 36125 28641 36159
rect 28675 36125 28687 36159
rect 28629 36119 28687 36125
rect 28718 36116 28724 36168
rect 28776 36156 28782 36168
rect 29733 36159 29791 36165
rect 28776 36128 28821 36156
rect 28776 36116 28782 36128
rect 29733 36125 29745 36159
rect 29779 36156 29791 36159
rect 30374 36156 30380 36168
rect 29779 36128 30380 36156
rect 29779 36125 29791 36128
rect 29733 36119 29791 36125
rect 30374 36116 30380 36128
rect 30432 36116 30438 36168
rect 32416 36165 32444 36332
rect 33686 36320 33692 36372
rect 33744 36360 33750 36372
rect 33781 36363 33839 36369
rect 33781 36360 33793 36363
rect 33744 36332 33793 36360
rect 33744 36320 33750 36332
rect 33781 36329 33793 36332
rect 33827 36329 33839 36363
rect 35342 36360 35348 36372
rect 35303 36332 35348 36360
rect 33781 36323 33839 36329
rect 35342 36320 35348 36332
rect 35400 36320 35406 36372
rect 33318 36184 33324 36236
rect 33376 36224 33382 36236
rect 33376 36196 34744 36224
rect 33376 36184 33382 36196
rect 32401 36159 32459 36165
rect 32401 36125 32413 36159
rect 32447 36156 32459 36159
rect 34422 36156 34428 36168
rect 32447 36128 34428 36156
rect 32447 36125 32459 36128
rect 32401 36119 32459 36125
rect 34422 36116 34428 36128
rect 34480 36116 34486 36168
rect 34716 36165 34744 36196
rect 34790 36184 34796 36236
rect 34848 36224 34854 36236
rect 34848 36196 35112 36224
rect 34848 36184 34854 36196
rect 34701 36159 34759 36165
rect 34701 36125 34713 36159
rect 34747 36125 34759 36159
rect 34882 36156 34888 36168
rect 34843 36128 34888 36156
rect 34701 36119 34759 36125
rect 34882 36116 34888 36128
rect 34940 36116 34946 36168
rect 35084 36165 35112 36196
rect 34977 36159 35035 36165
rect 34977 36125 34989 36159
rect 35023 36125 35035 36159
rect 34977 36119 35035 36125
rect 35069 36159 35127 36165
rect 35069 36125 35081 36159
rect 35115 36156 35127 36159
rect 36630 36156 36636 36168
rect 35115 36128 36636 36156
rect 35115 36125 35127 36128
rect 35069 36119 35127 36125
rect 29549 36091 29607 36097
rect 29549 36088 29561 36091
rect 28460 36060 29561 36088
rect 29549 36057 29561 36060
rect 29595 36057 29607 36091
rect 29917 36091 29975 36097
rect 29917 36088 29929 36091
rect 29549 36051 29607 36057
rect 29656 36060 29929 36088
rect 29656 36032 29684 36060
rect 29917 36057 29929 36060
rect 29963 36057 29975 36091
rect 33410 36088 33416 36100
rect 33371 36060 33416 36088
rect 29917 36051 29975 36057
rect 33410 36048 33416 36060
rect 33468 36048 33474 36100
rect 33597 36091 33655 36097
rect 33597 36057 33609 36091
rect 33643 36088 33655 36091
rect 34514 36088 34520 36100
rect 33643 36060 34520 36088
rect 33643 36057 33655 36060
rect 33597 36051 33655 36057
rect 34514 36048 34520 36060
rect 34572 36048 34578 36100
rect 9585 36023 9643 36029
rect 9585 35989 9597 36023
rect 9631 36020 9643 36023
rect 9674 36020 9680 36032
rect 9631 35992 9680 36020
rect 9631 35989 9643 35992
rect 9585 35983 9643 35989
rect 9674 35980 9680 35992
rect 9732 35980 9738 36032
rect 11422 36020 11428 36032
rect 11383 35992 11428 36020
rect 11422 35980 11428 35992
rect 11480 35980 11486 36032
rect 21726 35980 21732 36032
rect 21784 36020 21790 36032
rect 22005 36023 22063 36029
rect 22005 36020 22017 36023
rect 21784 35992 22017 36020
rect 21784 35980 21790 35992
rect 22005 35989 22017 35992
rect 22051 35989 22063 36023
rect 22005 35983 22063 35989
rect 22186 35980 22192 36032
rect 22244 36020 22250 36032
rect 22830 36020 22836 36032
rect 22244 35992 22836 36020
rect 22244 35980 22250 35992
rect 22830 35980 22836 35992
rect 22888 36020 22894 36032
rect 23109 36023 23167 36029
rect 23109 36020 23121 36023
rect 22888 35992 23121 36020
rect 22888 35980 22894 35992
rect 23109 35989 23121 35992
rect 23155 35989 23167 36023
rect 23109 35983 23167 35989
rect 23290 35980 23296 36032
rect 23348 36020 23354 36032
rect 23661 36023 23719 36029
rect 23661 36020 23673 36023
rect 23348 35992 23673 36020
rect 23348 35980 23354 35992
rect 23661 35989 23673 35992
rect 23707 35989 23719 36023
rect 27062 36020 27068 36032
rect 27023 35992 27068 36020
rect 23661 35983 23719 35989
rect 27062 35980 27068 35992
rect 27120 35980 27126 36032
rect 29638 35980 29644 36032
rect 29696 35980 29702 36032
rect 34238 35980 34244 36032
rect 34296 36020 34302 36032
rect 34992 36020 35020 36119
rect 36630 36116 36636 36128
rect 36688 36116 36694 36168
rect 58158 36156 58164 36168
rect 58119 36128 58164 36156
rect 58158 36116 58164 36128
rect 58216 36116 58222 36168
rect 34296 35992 35020 36020
rect 34296 35980 34302 35992
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 11422 35776 11428 35828
rect 11480 35816 11486 35828
rect 12250 35816 12256 35828
rect 11480 35788 12256 35816
rect 11480 35776 11486 35788
rect 12250 35776 12256 35788
rect 12308 35816 12314 35828
rect 13357 35819 13415 35825
rect 12308 35788 12572 35816
rect 12308 35776 12314 35788
rect 4985 35751 5043 35757
rect 4985 35717 4997 35751
rect 5031 35748 5043 35751
rect 5166 35748 5172 35760
rect 5031 35720 5172 35748
rect 5031 35717 5043 35720
rect 4985 35711 5043 35717
rect 5166 35708 5172 35720
rect 5224 35708 5230 35760
rect 9674 35708 9680 35760
rect 9732 35748 9738 35760
rect 12544 35757 12572 35788
rect 13357 35785 13369 35819
rect 13403 35816 13415 35819
rect 13722 35816 13728 35828
rect 13403 35788 13728 35816
rect 13403 35785 13415 35788
rect 13357 35779 13415 35785
rect 13722 35776 13728 35788
rect 13780 35816 13786 35828
rect 27062 35816 27068 35828
rect 13780 35788 27068 35816
rect 13780 35776 13786 35788
rect 27062 35776 27068 35788
rect 27120 35776 27126 35828
rect 34882 35776 34888 35828
rect 34940 35816 34946 35828
rect 35069 35819 35127 35825
rect 35069 35816 35081 35819
rect 34940 35788 35081 35816
rect 34940 35776 34946 35788
rect 35069 35785 35081 35788
rect 35115 35785 35127 35819
rect 35069 35779 35127 35785
rect 11885 35751 11943 35757
rect 11885 35748 11897 35751
rect 9732 35720 11897 35748
rect 9732 35708 9738 35720
rect 11885 35717 11897 35720
rect 11931 35748 11943 35751
rect 12345 35751 12403 35757
rect 12345 35748 12357 35751
rect 11931 35720 12357 35748
rect 11931 35717 11943 35720
rect 11885 35711 11943 35717
rect 12345 35717 12357 35720
rect 12391 35717 12403 35751
rect 12345 35711 12403 35717
rect 12529 35751 12587 35757
rect 12529 35717 12541 35751
rect 12575 35717 12587 35751
rect 12529 35711 12587 35717
rect 16114 35708 16120 35760
rect 16172 35748 16178 35760
rect 16172 35720 17632 35748
rect 16172 35708 16178 35720
rect 3602 35640 3608 35692
rect 3660 35680 3666 35692
rect 4801 35683 4859 35689
rect 4801 35680 4813 35683
rect 3660 35652 4813 35680
rect 3660 35640 3666 35652
rect 4801 35649 4813 35652
rect 4847 35680 4859 35683
rect 7282 35680 7288 35692
rect 4847 35652 7288 35680
rect 4847 35649 4859 35652
rect 4801 35643 4859 35649
rect 7282 35640 7288 35652
rect 7340 35680 7346 35692
rect 8297 35683 8355 35689
rect 8297 35680 8309 35683
rect 7340 35652 8309 35680
rect 7340 35640 7346 35652
rect 8297 35649 8309 35652
rect 8343 35649 8355 35683
rect 9858 35680 9864 35692
rect 9819 35652 9864 35680
rect 8297 35643 8355 35649
rect 9858 35640 9864 35652
rect 9916 35640 9922 35692
rect 11701 35683 11759 35689
rect 11701 35649 11713 35683
rect 11747 35680 11759 35683
rect 11790 35680 11796 35692
rect 11747 35652 11796 35680
rect 11747 35649 11759 35652
rect 11701 35643 11759 35649
rect 11790 35640 11796 35652
rect 11848 35640 11854 35692
rect 13170 35640 13176 35692
rect 13228 35680 13234 35692
rect 13265 35683 13323 35689
rect 13265 35680 13277 35683
rect 13228 35652 13277 35680
rect 13228 35640 13234 35652
rect 13265 35649 13277 35652
rect 13311 35680 13323 35683
rect 14461 35683 14519 35689
rect 14461 35680 14473 35683
rect 13311 35652 14473 35680
rect 13311 35649 13323 35652
rect 13265 35643 13323 35649
rect 14461 35649 14473 35652
rect 14507 35649 14519 35683
rect 17126 35680 17132 35692
rect 14461 35643 14519 35649
rect 15212 35652 17132 35680
rect 8021 35615 8079 35621
rect 8021 35581 8033 35615
rect 8067 35612 8079 35615
rect 8202 35612 8208 35624
rect 8067 35584 8208 35612
rect 8067 35581 8079 35584
rect 8021 35575 8079 35581
rect 8202 35572 8208 35584
rect 8260 35572 8266 35624
rect 9214 35572 9220 35624
rect 9272 35612 9278 35624
rect 9585 35615 9643 35621
rect 9585 35612 9597 35615
rect 9272 35584 9597 35612
rect 9272 35572 9278 35584
rect 9585 35581 9597 35584
rect 9631 35581 9643 35615
rect 10962 35612 10968 35624
rect 10875 35584 10968 35612
rect 9585 35575 9643 35581
rect 10962 35572 10968 35584
rect 11020 35612 11026 35624
rect 15212 35612 15240 35652
rect 17126 35640 17132 35652
rect 17184 35680 17190 35692
rect 17221 35683 17279 35689
rect 17221 35680 17233 35683
rect 17184 35652 17233 35680
rect 17184 35640 17190 35652
rect 17221 35649 17233 35652
rect 17267 35649 17279 35683
rect 17221 35643 17279 35649
rect 17313 35683 17371 35689
rect 17313 35649 17325 35683
rect 17359 35649 17371 35683
rect 17313 35643 17371 35649
rect 17328 35612 17356 35643
rect 17402 35640 17408 35692
rect 17460 35680 17466 35692
rect 17604 35689 17632 35720
rect 21818 35708 21824 35760
rect 21876 35748 21882 35760
rect 25038 35748 25044 35760
rect 21876 35720 25044 35748
rect 21876 35708 21882 35720
rect 24228 35692 24256 35720
rect 25038 35708 25044 35720
rect 25096 35708 25102 35760
rect 27798 35708 27804 35760
rect 27856 35748 27862 35760
rect 28442 35748 28448 35760
rect 27856 35720 28448 35748
rect 27856 35708 27862 35720
rect 28442 35708 28448 35720
rect 28500 35748 28506 35760
rect 30650 35748 30656 35760
rect 28500 35720 30656 35748
rect 28500 35708 28506 35720
rect 17589 35683 17647 35689
rect 17460 35652 17505 35680
rect 17460 35640 17466 35652
rect 17589 35649 17601 35683
rect 17635 35649 17647 35683
rect 17589 35643 17647 35649
rect 22186 35640 22192 35692
rect 22244 35680 22250 35692
rect 22649 35683 22707 35689
rect 22649 35680 22661 35683
rect 22244 35652 22661 35680
rect 22244 35640 22250 35652
rect 22649 35649 22661 35652
rect 22695 35649 22707 35683
rect 22649 35643 22707 35649
rect 22741 35683 22799 35689
rect 22741 35649 22753 35683
rect 22787 35649 22799 35683
rect 22741 35643 22799 35649
rect 11020 35584 15240 35612
rect 17052 35584 17356 35612
rect 11020 35572 11026 35584
rect 9490 35504 9496 35556
rect 9548 35544 9554 35556
rect 11517 35547 11575 35553
rect 11517 35544 11529 35547
rect 9548 35516 11529 35544
rect 9548 35504 9554 35516
rect 11517 35513 11529 35516
rect 11563 35513 11575 35547
rect 11517 35507 11575 35513
rect 12618 35504 12624 35556
rect 12676 35544 12682 35556
rect 13909 35547 13967 35553
rect 13909 35544 13921 35547
rect 12676 35516 13921 35544
rect 12676 35504 12682 35516
rect 13909 35513 13921 35516
rect 13955 35544 13967 35547
rect 14734 35544 14740 35556
rect 13955 35516 14740 35544
rect 13955 35513 13967 35516
rect 13909 35507 13967 35513
rect 14734 35504 14740 35516
rect 14792 35504 14798 35556
rect 15194 35504 15200 35556
rect 15252 35544 15258 35556
rect 17052 35544 17080 35584
rect 15252 35516 17080 35544
rect 15252 35504 15258 35516
rect 17126 35504 17132 35556
rect 17184 35544 17190 35556
rect 18049 35547 18107 35553
rect 18049 35544 18061 35547
rect 17184 35516 18061 35544
rect 17184 35504 17190 35516
rect 18049 35513 18061 35516
rect 18095 35544 18107 35547
rect 21174 35544 21180 35556
rect 18095 35516 21180 35544
rect 18095 35513 18107 35516
rect 18049 35507 18107 35513
rect 21174 35504 21180 35516
rect 21232 35504 21238 35556
rect 22756 35544 22784 35643
rect 22830 35640 22836 35692
rect 22888 35680 22894 35692
rect 23017 35683 23075 35689
rect 22888 35652 22933 35680
rect 22888 35640 22894 35652
rect 23017 35649 23029 35683
rect 23063 35680 23075 35683
rect 23382 35680 23388 35692
rect 23063 35652 23388 35680
rect 23063 35649 23075 35652
rect 23017 35643 23075 35649
rect 23382 35640 23388 35652
rect 23440 35640 23446 35692
rect 24210 35680 24216 35692
rect 24123 35652 24216 35680
rect 24210 35640 24216 35652
rect 24268 35640 24274 35692
rect 24302 35640 24308 35692
rect 24360 35680 24366 35692
rect 24469 35683 24527 35689
rect 24469 35680 24481 35683
rect 24360 35652 24481 35680
rect 24360 35640 24366 35652
rect 24469 35649 24481 35652
rect 24515 35649 24527 35683
rect 24469 35643 24527 35649
rect 27341 35683 27399 35689
rect 27341 35649 27353 35683
rect 27387 35680 27399 35683
rect 27430 35680 27436 35692
rect 27387 35652 27436 35680
rect 27387 35649 27399 35652
rect 27341 35643 27399 35649
rect 27430 35640 27436 35652
rect 27488 35640 27494 35692
rect 27614 35689 27620 35692
rect 27608 35643 27620 35689
rect 27672 35680 27678 35692
rect 30101 35683 30159 35689
rect 27672 35652 27708 35680
rect 27614 35640 27620 35643
rect 27672 35640 27678 35652
rect 30101 35649 30113 35683
rect 30147 35649 30159 35683
rect 30282 35680 30288 35692
rect 30243 35652 30288 35680
rect 30101 35643 30159 35649
rect 22848 35612 22876 35640
rect 23290 35612 23296 35624
rect 22848 35584 23296 35612
rect 23290 35572 23296 35584
rect 23348 35612 23354 35624
rect 23477 35615 23535 35621
rect 23477 35612 23489 35615
rect 23348 35584 23489 35612
rect 23348 35572 23354 35584
rect 23477 35581 23489 35584
rect 23523 35581 23535 35615
rect 30116 35612 30144 35643
rect 30282 35640 30288 35652
rect 30340 35640 30346 35692
rect 30392 35689 30420 35720
rect 30650 35708 30656 35720
rect 30708 35708 30714 35760
rect 30377 35683 30435 35689
rect 30377 35649 30389 35683
rect 30423 35649 30435 35683
rect 30377 35643 30435 35649
rect 30466 35640 30472 35692
rect 30524 35680 30530 35692
rect 30524 35652 30569 35680
rect 30524 35640 30530 35652
rect 33410 35640 33416 35692
rect 33468 35680 33474 35692
rect 34701 35683 34759 35689
rect 34701 35680 34713 35683
rect 33468 35652 34713 35680
rect 33468 35640 33474 35652
rect 34701 35649 34713 35652
rect 34747 35649 34759 35683
rect 34701 35643 34759 35649
rect 34885 35683 34943 35689
rect 34885 35649 34897 35683
rect 34931 35680 34943 35683
rect 35342 35680 35348 35692
rect 34931 35652 35348 35680
rect 34931 35649 34943 35652
rect 34885 35643 34943 35649
rect 35342 35640 35348 35652
rect 35400 35640 35406 35692
rect 30926 35612 30932 35624
rect 30116 35584 30932 35612
rect 23477 35575 23535 35581
rect 30926 35572 30932 35584
rect 30984 35572 30990 35624
rect 32125 35615 32183 35621
rect 32125 35612 32137 35615
rect 31726 35584 32137 35612
rect 29549 35547 29607 35553
rect 29549 35544 29561 35547
rect 22756 35516 24256 35544
rect 5166 35476 5172 35488
rect 5127 35448 5172 35476
rect 5166 35436 5172 35448
rect 5224 35436 5230 35488
rect 10778 35436 10784 35488
rect 10836 35476 10842 35488
rect 12713 35479 12771 35485
rect 12713 35476 12725 35479
rect 10836 35448 12725 35476
rect 10836 35436 10842 35448
rect 12713 35445 12725 35448
rect 12759 35445 12771 35479
rect 12713 35439 12771 35445
rect 16945 35479 17003 35485
rect 16945 35445 16957 35479
rect 16991 35476 17003 35479
rect 17218 35476 17224 35488
rect 16991 35448 17224 35476
rect 16991 35445 17003 35448
rect 16945 35439 17003 35445
rect 17218 35436 17224 35448
rect 17276 35436 17282 35488
rect 22462 35476 22468 35488
rect 22423 35448 22468 35476
rect 22462 35436 22468 35448
rect 22520 35436 22526 35488
rect 24228 35476 24256 35516
rect 28368 35516 29561 35544
rect 25593 35479 25651 35485
rect 25593 35476 25605 35479
rect 24228 35448 25605 35476
rect 25593 35445 25605 35448
rect 25639 35476 25651 35479
rect 26418 35476 26424 35488
rect 25639 35448 26424 35476
rect 25639 35445 25651 35448
rect 25593 35439 25651 35445
rect 26418 35436 26424 35448
rect 26476 35436 26482 35488
rect 27522 35436 27528 35488
rect 27580 35476 27586 35488
rect 28368 35476 28396 35516
rect 29549 35513 29561 35516
rect 29595 35544 29607 35547
rect 30466 35544 30472 35556
rect 29595 35516 30472 35544
rect 29595 35513 29607 35516
rect 29549 35507 29607 35513
rect 30466 35504 30472 35516
rect 30524 35504 30530 35556
rect 27580 35448 28396 35476
rect 27580 35436 27586 35448
rect 28442 35436 28448 35488
rect 28500 35476 28506 35488
rect 28721 35479 28779 35485
rect 28721 35476 28733 35479
rect 28500 35448 28733 35476
rect 28500 35436 28506 35448
rect 28721 35445 28733 35448
rect 28767 35445 28779 35479
rect 30742 35476 30748 35488
rect 30703 35448 30748 35476
rect 28721 35439 28779 35445
rect 30742 35436 30748 35448
rect 30800 35436 30806 35488
rect 31478 35476 31484 35488
rect 31439 35448 31484 35476
rect 31478 35436 31484 35448
rect 31536 35476 31542 35488
rect 31726 35476 31754 35584
rect 32125 35581 32137 35584
rect 32171 35581 32183 35615
rect 32125 35575 32183 35581
rect 32401 35615 32459 35621
rect 32401 35581 32413 35615
rect 32447 35612 32459 35615
rect 33318 35612 33324 35624
rect 32447 35584 33324 35612
rect 32447 35581 32459 35584
rect 32401 35575 32459 35581
rect 33318 35572 33324 35584
rect 33376 35572 33382 35624
rect 31536 35448 31754 35476
rect 31536 35436 31542 35448
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 4706 35272 4712 35284
rect 4667 35244 4712 35272
rect 4706 35232 4712 35244
rect 4764 35232 4770 35284
rect 11790 35272 11796 35284
rect 5092 35244 8156 35272
rect 11751 35244 11796 35272
rect 2682 35096 2688 35148
rect 2740 35136 2746 35148
rect 5092 35136 5120 35244
rect 8128 35216 8156 35244
rect 11790 35232 11796 35244
rect 11848 35232 11854 35284
rect 17310 35232 17316 35284
rect 17368 35272 17374 35284
rect 21085 35275 21143 35281
rect 21085 35272 21097 35275
rect 17368 35244 21097 35272
rect 17368 35232 17374 35244
rect 8110 35204 8116 35216
rect 8071 35176 8116 35204
rect 8110 35164 8116 35176
rect 8168 35164 8174 35216
rect 9766 35136 9772 35148
rect 2740 35108 5120 35136
rect 2740 35096 2746 35108
rect 5092 35077 5120 35108
rect 9324 35108 9772 35136
rect 4985 35071 5043 35077
rect 4985 35037 4997 35071
rect 5031 35037 5043 35071
rect 4985 35031 5043 35037
rect 5077 35071 5135 35077
rect 5077 35037 5089 35071
rect 5123 35037 5135 35071
rect 5077 35031 5135 35037
rect 5000 35000 5028 35031
rect 5166 35028 5172 35080
rect 5224 35068 5230 35080
rect 5353 35071 5411 35077
rect 5224 35040 5269 35068
rect 5224 35028 5230 35040
rect 5353 35037 5365 35071
rect 5399 35037 5411 35071
rect 5353 35031 5411 35037
rect 6089 35071 6147 35077
rect 6089 35037 6101 35071
rect 6135 35068 6147 35071
rect 6822 35068 6828 35080
rect 6135 35040 6828 35068
rect 6135 35037 6147 35040
rect 6089 35031 6147 35037
rect 5258 35000 5264 35012
rect 5000 34972 5264 35000
rect 5258 34960 5264 34972
rect 5316 34960 5322 35012
rect 2958 34892 2964 34944
rect 3016 34932 3022 34944
rect 5368 34932 5396 35031
rect 6822 35028 6828 35040
rect 6880 35028 6886 35080
rect 8297 35071 8355 35077
rect 8297 35037 8309 35071
rect 8343 35068 8355 35071
rect 9214 35068 9220 35080
rect 8343 35040 9220 35068
rect 8343 35037 8355 35040
rect 8297 35031 8355 35037
rect 9214 35028 9220 35040
rect 9272 35028 9278 35080
rect 9324 35077 9352 35108
rect 9766 35096 9772 35108
rect 9824 35096 9830 35148
rect 10410 35136 10416 35148
rect 10371 35108 10416 35136
rect 10410 35096 10416 35108
rect 10468 35096 10474 35148
rect 9309 35071 9367 35077
rect 9309 35037 9321 35071
rect 9355 35037 9367 35071
rect 9490 35068 9496 35080
rect 9451 35040 9496 35068
rect 9309 35031 9367 35037
rect 9490 35028 9496 35040
rect 9548 35028 9554 35080
rect 9585 35071 9643 35077
rect 9585 35037 9597 35071
rect 9631 35037 9643 35071
rect 9585 35031 9643 35037
rect 9677 35071 9735 35077
rect 9677 35037 9689 35071
rect 9723 35068 9735 35071
rect 10962 35068 10968 35080
rect 9723 35040 10968 35068
rect 9723 35037 9735 35040
rect 9677 35031 9735 35037
rect 6356 35003 6414 35009
rect 6356 34969 6368 35003
rect 6402 35000 6414 35003
rect 7006 35000 7012 35012
rect 6402 34972 7012 35000
rect 6402 34969 6414 34972
rect 6356 34963 6414 34969
rect 7006 34960 7012 34972
rect 7064 34960 7070 35012
rect 9600 35000 9628 35031
rect 10962 35028 10968 35040
rect 11020 35028 11026 35080
rect 11808 35068 11836 35232
rect 13538 35136 13544 35148
rect 13280 35108 13544 35136
rect 13280 35077 13308 35108
rect 13538 35096 13544 35108
rect 13596 35096 13602 35148
rect 12989 35071 13047 35077
rect 12989 35068 13001 35071
rect 11808 35040 13001 35068
rect 12989 35037 13001 35040
rect 13035 35037 13047 35071
rect 12989 35031 13047 35037
rect 13265 35071 13323 35077
rect 13265 35037 13277 35071
rect 13311 35037 13323 35071
rect 13265 35031 13323 35037
rect 13357 35071 13415 35077
rect 13357 35037 13369 35071
rect 13403 35037 13415 35071
rect 17126 35068 17132 35080
rect 17087 35040 17132 35068
rect 13357 35031 13415 35037
rect 9858 35000 9864 35012
rect 9600 34972 9864 35000
rect 9858 34960 9864 34972
rect 9916 34960 9922 35012
rect 9953 35003 10011 35009
rect 9953 34969 9965 35003
rect 9999 35000 10011 35003
rect 10658 35003 10716 35009
rect 10658 35000 10670 35003
rect 9999 34972 10670 35000
rect 9999 34969 10011 34972
rect 9953 34963 10011 34969
rect 10658 34969 10670 34972
rect 10704 34969 10716 35003
rect 10658 34963 10716 34969
rect 12434 34960 12440 35012
rect 12492 35000 12498 35012
rect 13173 35003 13231 35009
rect 13173 35000 13185 35003
rect 12492 34972 13185 35000
rect 12492 34960 12498 34972
rect 13173 34969 13185 34972
rect 13219 34969 13231 35003
rect 13173 34963 13231 34969
rect 3016 34904 5396 34932
rect 7469 34935 7527 34941
rect 3016 34892 3022 34904
rect 7469 34901 7481 34935
rect 7515 34932 7527 34935
rect 7558 34932 7564 34944
rect 7515 34904 7564 34932
rect 7515 34901 7527 34904
rect 7469 34895 7527 34901
rect 7558 34892 7564 34904
rect 7616 34892 7622 34944
rect 12802 34892 12808 34944
rect 12860 34932 12866 34944
rect 13372 34932 13400 35031
rect 17126 35028 17132 35040
rect 17184 35028 17190 35080
rect 17218 35028 17224 35080
rect 17276 35068 17282 35080
rect 17385 35071 17443 35077
rect 17385 35068 17397 35071
rect 17276 35040 17397 35068
rect 17276 35028 17282 35040
rect 17385 35037 17397 35040
rect 17431 35037 17443 35071
rect 17385 35031 17443 35037
rect 19889 35071 19947 35077
rect 19889 35037 19901 35071
rect 19935 35068 19947 35071
rect 20070 35068 20076 35080
rect 19935 35040 20076 35068
rect 19935 35037 19947 35040
rect 19889 35031 19947 35037
rect 20070 35028 20076 35040
rect 20128 35028 20134 35080
rect 20732 35068 20760 35244
rect 21085 35241 21097 35244
rect 21131 35241 21143 35275
rect 21085 35235 21143 35241
rect 24762 35232 24768 35284
rect 24820 35272 24826 35284
rect 25774 35272 25780 35284
rect 24820 35244 25780 35272
rect 24820 35232 24826 35244
rect 25774 35232 25780 35244
rect 25832 35232 25838 35284
rect 27433 35275 27491 35281
rect 27433 35241 27445 35275
rect 27479 35272 27491 35275
rect 27614 35272 27620 35284
rect 27479 35244 27620 35272
rect 27479 35241 27491 35244
rect 27433 35235 27491 35241
rect 27614 35232 27620 35244
rect 27672 35232 27678 35284
rect 20806 35164 20812 35216
rect 20864 35204 20870 35216
rect 20864 35176 24164 35204
rect 20864 35164 20870 35176
rect 22741 35139 22799 35145
rect 22741 35136 22753 35139
rect 22112 35108 22753 35136
rect 22112 35077 22140 35108
rect 22741 35105 22753 35108
rect 22787 35105 22799 35139
rect 22741 35099 22799 35105
rect 21913 35071 21971 35077
rect 21913 35068 21925 35071
rect 20732 35040 21925 35068
rect 21913 35037 21925 35040
rect 21959 35037 21971 35071
rect 21913 35031 21971 35037
rect 22005 35071 22063 35077
rect 22005 35037 22017 35071
rect 22051 35037 22063 35071
rect 22005 35031 22063 35037
rect 22097 35071 22155 35077
rect 22097 35037 22109 35071
rect 22143 35037 22155 35071
rect 22097 35031 22155 35037
rect 18690 34960 18696 35012
rect 18748 35000 18754 35012
rect 19705 35003 19763 35009
rect 19705 35000 19717 35003
rect 18748 34972 19717 35000
rect 18748 34960 18754 34972
rect 19705 34969 19717 34972
rect 19751 35000 19763 35003
rect 20714 35000 20720 35012
rect 19751 34972 20720 35000
rect 19751 34969 19763 34972
rect 19705 34963 19763 34969
rect 20714 34960 20720 34972
rect 20772 34960 20778 35012
rect 22020 35000 22048 35031
rect 22278 35028 22284 35080
rect 22336 35068 22342 35080
rect 22554 35068 22560 35080
rect 22336 35040 22560 35068
rect 22336 35028 22342 35040
rect 22554 35028 22560 35040
rect 22612 35028 22618 35080
rect 24136 35068 24164 35176
rect 27062 35164 27068 35216
rect 27120 35204 27126 35216
rect 27120 35176 28028 35204
rect 27120 35164 27126 35176
rect 24210 35096 24216 35148
rect 24268 35136 24274 35148
rect 24397 35139 24455 35145
rect 24397 35136 24409 35139
rect 24268 35108 24409 35136
rect 24268 35096 24274 35108
rect 24397 35105 24409 35108
rect 24443 35105 24455 35139
rect 27522 35136 27528 35148
rect 24397 35099 24455 35105
rect 26252 35108 27528 35136
rect 26252 35068 26280 35108
rect 27522 35096 27528 35108
rect 27580 35096 27586 35148
rect 27614 35096 27620 35148
rect 27672 35136 27678 35148
rect 27672 35108 27841 35136
rect 27672 35096 27678 35108
rect 26418 35068 26424 35080
rect 24136 35040 26280 35068
rect 26379 35040 26424 35068
rect 26418 35028 26424 35040
rect 26476 35028 26482 35080
rect 27706 35068 27712 35080
rect 27667 35040 27712 35068
rect 27706 35028 27712 35040
rect 27764 35028 27770 35080
rect 27813 35074 27841 35108
rect 27798 35068 27856 35074
rect 27798 35034 27810 35068
rect 27844 35034 27856 35068
rect 27798 35028 27856 35034
rect 27893 35071 27951 35077
rect 27893 35037 27905 35071
rect 27939 35037 27951 35071
rect 28000 35068 28028 35176
rect 32033 35139 32091 35145
rect 32033 35105 32045 35139
rect 32079 35136 32091 35139
rect 33134 35136 33140 35148
rect 32079 35108 33140 35136
rect 32079 35105 32091 35108
rect 32033 35099 32091 35105
rect 33134 35096 33140 35108
rect 33192 35096 33198 35148
rect 28077 35071 28135 35077
rect 28077 35068 28089 35071
rect 28000 35040 28089 35068
rect 27893 35031 27951 35037
rect 28077 35037 28089 35040
rect 28123 35037 28135 35071
rect 28077 35031 28135 35037
rect 21928 34972 22048 35000
rect 21928 34944 21956 34972
rect 22738 34960 22744 35012
rect 22796 35000 22802 35012
rect 22925 35003 22983 35009
rect 22925 35000 22937 35003
rect 22796 34972 22937 35000
rect 22796 34960 22802 34972
rect 22925 34969 22937 34972
rect 22971 34969 22983 35003
rect 22925 34963 22983 34969
rect 23014 34960 23020 35012
rect 23072 35000 23078 35012
rect 23109 35003 23167 35009
rect 23109 35000 23121 35003
rect 23072 34972 23121 35000
rect 23072 34960 23078 34972
rect 23109 34969 23121 34972
rect 23155 34969 23167 35003
rect 23109 34963 23167 34969
rect 24486 34960 24492 35012
rect 24544 35000 24550 35012
rect 24642 35003 24700 35009
rect 24642 35000 24654 35003
rect 24544 34972 24654 35000
rect 24544 34960 24550 34972
rect 24642 34969 24654 34972
rect 24688 34969 24700 35003
rect 26605 35003 26663 35009
rect 26605 35000 26617 35003
rect 24642 34963 24700 34969
rect 25976 34972 26617 35000
rect 25976 34944 26004 34972
rect 26605 34969 26617 34972
rect 26651 34969 26663 35003
rect 27908 35000 27936 35031
rect 28442 35028 28448 35080
rect 28500 35068 28506 35080
rect 28721 35071 28779 35077
rect 28721 35068 28733 35071
rect 28500 35040 28733 35068
rect 28500 35028 28506 35040
rect 28721 35037 28733 35040
rect 28767 35037 28779 35071
rect 28721 35031 28779 35037
rect 30742 35028 30748 35080
rect 30800 35068 30806 35080
rect 31766 35071 31824 35077
rect 31766 35068 31778 35071
rect 30800 35040 31778 35068
rect 30800 35028 30806 35040
rect 31766 35037 31778 35040
rect 31812 35037 31824 35071
rect 31766 35031 31824 35037
rect 32122 35028 32128 35080
rect 32180 35068 32186 35080
rect 32493 35071 32551 35077
rect 32493 35068 32505 35071
rect 32180 35040 32505 35068
rect 32180 35028 32186 35040
rect 32493 35037 32505 35040
rect 32539 35037 32551 35071
rect 32766 35068 32772 35080
rect 32727 35040 32772 35068
rect 32493 35031 32551 35037
rect 32766 35028 32772 35040
rect 32824 35028 32830 35080
rect 58158 35068 58164 35080
rect 58119 35040 58164 35068
rect 58158 35028 58164 35040
rect 58216 35028 58222 35080
rect 28537 35003 28595 35009
rect 28537 35000 28549 35003
rect 27908 34972 28549 35000
rect 26605 34963 26663 34969
rect 28537 34969 28549 34972
rect 28583 34969 28595 35003
rect 28537 34963 28595 34969
rect 28905 35003 28963 35009
rect 28905 34969 28917 35003
rect 28951 35000 28963 35003
rect 29546 35000 29552 35012
rect 28951 34972 29552 35000
rect 28951 34969 28963 34972
rect 28905 34963 28963 34969
rect 29546 34960 29552 34972
rect 29604 34960 29610 35012
rect 12860 34904 13400 34932
rect 13541 34935 13599 34941
rect 12860 34892 12866 34904
rect 13541 34901 13553 34935
rect 13587 34932 13599 34935
rect 18322 34932 18328 34944
rect 13587 34904 18328 34932
rect 13587 34901 13599 34904
rect 13541 34895 13599 34901
rect 18322 34892 18328 34904
rect 18380 34892 18386 34944
rect 18506 34932 18512 34944
rect 18467 34904 18512 34932
rect 18506 34892 18512 34904
rect 18564 34892 18570 34944
rect 19978 34892 19984 34944
rect 20036 34932 20042 34944
rect 20073 34935 20131 34941
rect 20073 34932 20085 34935
rect 20036 34904 20085 34932
rect 20036 34892 20042 34904
rect 20073 34901 20085 34904
rect 20119 34901 20131 34935
rect 21634 34932 21640 34944
rect 21595 34904 21640 34932
rect 20073 34895 20131 34901
rect 21634 34892 21640 34904
rect 21692 34892 21698 34944
rect 21910 34892 21916 34944
rect 21968 34892 21974 34944
rect 23842 34932 23848 34944
rect 23803 34904 23848 34932
rect 23842 34892 23848 34904
rect 23900 34892 23906 34944
rect 24210 34892 24216 34944
rect 24268 34932 24274 34944
rect 24946 34932 24952 34944
rect 24268 34904 24952 34932
rect 24268 34892 24274 34904
rect 24946 34892 24952 34904
rect 25004 34932 25010 34944
rect 25958 34932 25964 34944
rect 25004 34904 25964 34932
rect 25004 34892 25010 34904
rect 25958 34892 25964 34904
rect 26016 34892 26022 34944
rect 26234 34932 26240 34944
rect 26195 34904 26240 34932
rect 26234 34892 26240 34904
rect 26292 34892 26298 34944
rect 29638 34892 29644 34944
rect 29696 34932 29702 34944
rect 30101 34935 30159 34941
rect 30101 34932 30113 34935
rect 29696 34904 30113 34932
rect 29696 34892 29702 34904
rect 30101 34901 30113 34904
rect 30147 34901 30159 34935
rect 30101 34895 30159 34901
rect 30190 34892 30196 34944
rect 30248 34932 30254 34944
rect 30653 34935 30711 34941
rect 30653 34932 30665 34935
rect 30248 34904 30665 34932
rect 30248 34892 30254 34904
rect 30653 34901 30665 34904
rect 30699 34932 30711 34935
rect 31110 34932 31116 34944
rect 30699 34904 31116 34932
rect 30699 34901 30711 34904
rect 30653 34895 30711 34901
rect 31110 34892 31116 34904
rect 31168 34892 31174 34944
rect 33873 34935 33931 34941
rect 33873 34901 33885 34935
rect 33919 34932 33931 34935
rect 34054 34932 34060 34944
rect 33919 34904 34060 34932
rect 33919 34901 33931 34904
rect 33873 34895 33931 34901
rect 34054 34892 34060 34904
rect 34112 34892 34118 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 3881 34731 3939 34737
rect 3881 34697 3893 34731
rect 3927 34697 3939 34731
rect 7006 34728 7012 34740
rect 6967 34700 7012 34728
rect 3881 34691 3939 34697
rect 3896 34660 3924 34691
rect 7006 34688 7012 34700
rect 7064 34688 7070 34740
rect 10318 34728 10324 34740
rect 10279 34700 10324 34728
rect 10318 34688 10324 34700
rect 10376 34688 10382 34740
rect 10410 34688 10416 34740
rect 10468 34728 10474 34740
rect 12618 34728 12624 34740
rect 10468 34700 12624 34728
rect 10468 34688 10474 34700
rect 12618 34688 12624 34700
rect 12676 34688 12682 34740
rect 12805 34731 12863 34737
rect 12805 34697 12817 34731
rect 12851 34728 12863 34731
rect 16666 34728 16672 34740
rect 12851 34700 16672 34728
rect 12851 34697 12863 34700
rect 12805 34691 12863 34697
rect 16666 34688 16672 34700
rect 16724 34688 16730 34740
rect 17313 34731 17371 34737
rect 17313 34697 17325 34731
rect 17359 34728 17371 34731
rect 17402 34728 17408 34740
rect 17359 34700 17408 34728
rect 17359 34697 17371 34700
rect 17313 34691 17371 34697
rect 17402 34688 17408 34700
rect 17460 34688 17466 34740
rect 19889 34731 19947 34737
rect 19889 34728 19901 34731
rect 19168 34700 19901 34728
rect 4525 34663 4583 34669
rect 4525 34660 4537 34663
rect 3896 34632 4537 34660
rect 4525 34629 4537 34632
rect 4571 34660 4583 34663
rect 5442 34660 5448 34672
rect 4571 34632 5448 34660
rect 4571 34629 4583 34632
rect 4525 34623 4583 34629
rect 5442 34620 5448 34632
rect 5500 34620 5506 34672
rect 7190 34620 7196 34672
rect 7248 34660 7254 34672
rect 8205 34663 8263 34669
rect 7248 34632 7328 34660
rect 7248 34620 7254 34632
rect 2774 34601 2780 34604
rect 2768 34555 2780 34601
rect 2832 34592 2838 34604
rect 4706 34592 4712 34604
rect 2832 34564 2868 34592
rect 4667 34564 4712 34592
rect 2774 34552 2780 34555
rect 2832 34552 2838 34564
rect 4706 34552 4712 34564
rect 4764 34552 4770 34604
rect 7300 34601 7328 34632
rect 8205 34629 8217 34663
rect 8251 34660 8263 34663
rect 10502 34660 10508 34672
rect 8251 34632 10508 34660
rect 8251 34629 8263 34632
rect 8205 34623 8263 34629
rect 7285 34595 7343 34601
rect 7285 34561 7297 34595
rect 7331 34561 7343 34595
rect 7285 34555 7343 34561
rect 7377 34595 7435 34601
rect 7377 34561 7389 34595
rect 7423 34561 7435 34595
rect 7377 34555 7435 34561
rect 2406 34484 2412 34536
rect 2464 34524 2470 34536
rect 2501 34527 2559 34533
rect 2501 34524 2513 34527
rect 2464 34496 2513 34524
rect 2464 34484 2470 34496
rect 2501 34493 2513 34496
rect 2547 34493 2559 34527
rect 5534 34524 5540 34536
rect 5447 34496 5540 34524
rect 2501 34487 2559 34493
rect 5534 34484 5540 34496
rect 5592 34524 5598 34536
rect 5718 34524 5724 34536
rect 5592 34496 5724 34524
rect 5592 34484 5598 34496
rect 5718 34484 5724 34496
rect 5776 34484 5782 34536
rect 7190 34484 7196 34536
rect 7248 34524 7254 34536
rect 7392 34524 7420 34555
rect 7466 34552 7472 34604
rect 7524 34592 7530 34604
rect 7653 34595 7711 34601
rect 7524 34564 7569 34592
rect 7524 34552 7530 34564
rect 7653 34561 7665 34595
rect 7699 34592 7711 34595
rect 8220 34592 8248 34623
rect 10502 34620 10508 34632
rect 10560 34620 10566 34672
rect 12529 34663 12587 34669
rect 12529 34629 12541 34663
rect 12575 34660 12587 34663
rect 12894 34660 12900 34672
rect 12575 34632 12900 34660
rect 12575 34629 12587 34632
rect 12529 34623 12587 34629
rect 12894 34620 12900 34632
rect 12952 34620 12958 34672
rect 17497 34663 17555 34669
rect 17497 34629 17509 34663
rect 17543 34660 17555 34663
rect 18506 34660 18512 34672
rect 17543 34632 18512 34660
rect 17543 34629 17555 34632
rect 17497 34623 17555 34629
rect 18506 34620 18512 34632
rect 18564 34660 18570 34672
rect 18564 34632 18920 34660
rect 18564 34620 18570 34632
rect 10594 34592 10600 34604
rect 7699 34564 8248 34592
rect 10555 34564 10600 34592
rect 7699 34561 7711 34564
rect 7653 34555 7711 34561
rect 10594 34552 10600 34564
rect 10652 34552 10658 34604
rect 10689 34595 10747 34601
rect 10689 34561 10701 34595
rect 10735 34561 10747 34595
rect 10689 34555 10747 34561
rect 7248 34496 7420 34524
rect 7248 34484 7254 34496
rect 9858 34484 9864 34536
rect 9916 34524 9922 34536
rect 10704 34524 10732 34555
rect 10778 34552 10784 34604
rect 10836 34592 10842 34604
rect 10965 34595 11023 34601
rect 10836 34564 10881 34592
rect 10836 34552 10842 34564
rect 10965 34561 10977 34595
rect 11011 34592 11023 34595
rect 11146 34592 11152 34604
rect 11011 34564 11152 34592
rect 11011 34561 11023 34564
rect 10965 34555 11023 34561
rect 11146 34552 11152 34564
rect 11204 34552 11210 34604
rect 12250 34592 12256 34604
rect 12211 34564 12256 34592
rect 12250 34552 12256 34564
rect 12308 34552 12314 34604
rect 12434 34552 12440 34604
rect 12492 34592 12498 34604
rect 12621 34595 12679 34601
rect 12492 34564 12537 34592
rect 12492 34552 12498 34564
rect 12621 34561 12633 34595
rect 12667 34592 12679 34595
rect 12802 34592 12808 34604
rect 12667 34564 12808 34592
rect 12667 34561 12679 34564
rect 12621 34555 12679 34561
rect 12802 34552 12808 34564
rect 12860 34552 12866 34604
rect 17678 34592 17684 34604
rect 17639 34564 17684 34592
rect 17678 34552 17684 34564
rect 17736 34552 17742 34604
rect 18322 34552 18328 34604
rect 18380 34592 18386 34604
rect 18892 34601 18920 34632
rect 18966 34620 18972 34672
rect 19024 34660 19030 34672
rect 19168 34669 19196 34700
rect 19889 34697 19901 34700
rect 19935 34728 19947 34731
rect 20070 34728 20076 34740
rect 19935 34700 20076 34728
rect 19935 34697 19947 34700
rect 19889 34691 19947 34697
rect 20070 34688 20076 34700
rect 20128 34688 20134 34740
rect 20732 34700 22600 34728
rect 19061 34663 19119 34669
rect 19061 34660 19073 34663
rect 19024 34632 19073 34660
rect 19024 34620 19030 34632
rect 19061 34629 19073 34632
rect 19107 34629 19119 34663
rect 19061 34623 19119 34629
rect 19150 34663 19208 34669
rect 19150 34629 19162 34663
rect 19196 34629 19208 34663
rect 20732 34660 20760 34700
rect 19150 34623 19208 34629
rect 20640 34632 20760 34660
rect 18785 34595 18843 34601
rect 18785 34592 18797 34595
rect 18380 34564 18797 34592
rect 18380 34552 18386 34564
rect 18785 34561 18797 34564
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 18878 34595 18936 34601
rect 18878 34561 18890 34595
rect 18924 34561 18936 34595
rect 19269 34595 19327 34601
rect 19269 34592 19281 34595
rect 18878 34555 18936 34561
rect 19168 34564 19281 34592
rect 19168 34536 19196 34564
rect 19269 34561 19281 34564
rect 19315 34561 19327 34595
rect 20640 34592 20668 34632
rect 21634 34620 21640 34672
rect 21692 34660 21698 34672
rect 22066 34663 22124 34669
rect 22066 34660 22078 34663
rect 21692 34632 22078 34660
rect 21692 34620 21698 34632
rect 22066 34629 22078 34632
rect 22112 34629 22124 34663
rect 22572 34660 22600 34700
rect 22738 34688 22744 34740
rect 22796 34728 22802 34740
rect 23201 34731 23259 34737
rect 23201 34728 23213 34731
rect 22796 34700 23213 34728
rect 22796 34688 22802 34700
rect 23201 34697 23213 34700
rect 23247 34697 23259 34731
rect 24486 34728 24492 34740
rect 24447 34700 24492 34728
rect 23201 34691 23259 34697
rect 24486 34688 24492 34700
rect 24544 34688 24550 34740
rect 27062 34728 27068 34740
rect 24596 34700 26096 34728
rect 27023 34700 27068 34728
rect 23106 34660 23112 34672
rect 22572 34632 23112 34660
rect 22066 34623 22124 34629
rect 23106 34620 23112 34632
rect 23164 34620 23170 34672
rect 23658 34620 23664 34672
rect 23716 34660 23722 34672
rect 24029 34663 24087 34669
rect 24029 34660 24041 34663
rect 23716 34632 24041 34660
rect 23716 34620 23722 34632
rect 24029 34629 24041 34632
rect 24075 34660 24087 34663
rect 24596 34660 24624 34700
rect 25774 34660 25780 34672
rect 24075 34632 24624 34660
rect 25735 34632 25780 34660
rect 24075 34629 24087 34632
rect 24029 34623 24087 34629
rect 19269 34555 19327 34561
rect 19444 34564 20668 34592
rect 9916 34496 10732 34524
rect 9916 34484 9922 34496
rect 19150 34484 19156 34536
rect 19208 34484 19214 34536
rect 19444 34465 19472 34564
rect 20714 34552 20720 34604
rect 20772 34592 20778 34604
rect 21002 34595 21060 34601
rect 21002 34592 21014 34595
rect 20772 34564 21014 34592
rect 20772 34552 20778 34564
rect 21002 34561 21014 34564
rect 21048 34561 21060 34595
rect 21002 34555 21060 34561
rect 21269 34595 21327 34601
rect 21269 34561 21281 34595
rect 21315 34592 21327 34595
rect 21818 34592 21824 34604
rect 21315 34564 21824 34592
rect 21315 34561 21327 34564
rect 21269 34555 21327 34561
rect 21818 34552 21824 34564
rect 21876 34552 21882 34604
rect 24596 34592 24624 34632
rect 25774 34620 25780 34632
rect 25832 34620 25838 34672
rect 25958 34660 25964 34672
rect 25919 34632 25964 34660
rect 25958 34620 25964 34632
rect 26016 34620 26022 34672
rect 26068 34660 26096 34700
rect 27062 34688 27068 34700
rect 27120 34688 27126 34740
rect 27617 34731 27675 34737
rect 27617 34697 27629 34731
rect 27663 34728 27675 34731
rect 27706 34728 27712 34740
rect 27663 34700 27712 34728
rect 27663 34697 27675 34700
rect 27617 34691 27675 34697
rect 27706 34688 27712 34700
rect 27764 34688 27770 34740
rect 29917 34731 29975 34737
rect 29917 34697 29929 34731
rect 29963 34728 29975 34731
rect 30282 34728 30288 34740
rect 29963 34700 30288 34728
rect 29963 34697 29975 34700
rect 29917 34691 29975 34697
rect 30282 34688 30288 34700
rect 30340 34688 30346 34740
rect 32309 34731 32367 34737
rect 32309 34697 32321 34731
rect 32355 34728 32367 34731
rect 34790 34728 34796 34740
rect 32355 34700 33180 34728
rect 32355 34697 32367 34700
rect 32309 34691 32367 34697
rect 29733 34663 29791 34669
rect 26068 34632 29684 34660
rect 24719 34595 24777 34601
rect 24719 34592 24731 34595
rect 24596 34564 24731 34592
rect 24719 34561 24731 34564
rect 24765 34561 24777 34595
rect 24854 34592 24860 34604
rect 24815 34564 24860 34592
rect 24719 34555 24777 34561
rect 24854 34552 24860 34564
rect 24912 34552 24918 34604
rect 24949 34595 25007 34601
rect 24949 34561 24961 34595
rect 24995 34561 25007 34595
rect 25130 34592 25136 34604
rect 25091 34564 25136 34592
rect 24949 34555 25007 34561
rect 24964 34524 24992 34555
rect 25130 34552 25136 34564
rect 25188 34552 25194 34604
rect 29546 34592 29552 34604
rect 29507 34564 29552 34592
rect 29546 34552 29552 34564
rect 29604 34552 29610 34604
rect 29656 34592 29684 34632
rect 29733 34629 29745 34663
rect 29779 34660 29791 34663
rect 30190 34660 30196 34672
rect 29779 34632 30196 34660
rect 29779 34629 29791 34632
rect 29733 34623 29791 34629
rect 30190 34620 30196 34632
rect 30248 34620 30254 34672
rect 33042 34660 33048 34672
rect 30576 34632 33048 34660
rect 30576 34592 30604 34632
rect 33042 34620 33048 34632
rect 33100 34620 33106 34672
rect 30926 34592 30932 34604
rect 29656 34564 30604 34592
rect 30887 34564 30932 34592
rect 30926 34552 30932 34564
rect 30984 34552 30990 34604
rect 32122 34592 32128 34604
rect 32083 34564 32128 34592
rect 32122 34552 32128 34564
rect 32180 34552 32186 34604
rect 33152 34601 33180 34700
rect 33336 34700 34796 34728
rect 33336 34669 33364 34700
rect 34790 34688 34796 34700
rect 34848 34688 34854 34740
rect 33321 34663 33379 34669
rect 33321 34629 33333 34663
rect 33367 34629 33379 34663
rect 33321 34623 33379 34629
rect 33505 34663 33563 34669
rect 33505 34629 33517 34663
rect 33551 34660 33563 34663
rect 33551 34632 34192 34660
rect 33551 34629 33563 34632
rect 33505 34623 33563 34629
rect 33137 34595 33195 34601
rect 33137 34561 33149 34595
rect 33183 34592 33195 34595
rect 33410 34592 33416 34604
rect 33183 34564 33416 34592
rect 33183 34561 33195 34564
rect 33137 34555 33195 34561
rect 33410 34552 33416 34564
rect 33468 34552 33474 34604
rect 34164 34601 34192 34632
rect 33965 34595 34023 34601
rect 33965 34561 33977 34595
rect 34011 34561 34023 34595
rect 33965 34555 34023 34561
rect 34149 34595 34207 34601
rect 34149 34561 34161 34595
rect 34195 34561 34207 34595
rect 34149 34555 34207 34561
rect 34244 34595 34302 34601
rect 34244 34561 34256 34595
rect 34290 34561 34302 34595
rect 34244 34555 34302 34561
rect 34333 34595 34391 34601
rect 34333 34561 34345 34595
rect 34379 34561 34391 34595
rect 34333 34555 34391 34561
rect 25593 34527 25651 34533
rect 25593 34524 25605 34527
rect 24964 34496 25605 34524
rect 25593 34493 25605 34496
rect 25639 34493 25651 34527
rect 25593 34487 25651 34493
rect 29638 34484 29644 34536
rect 29696 34524 29702 34536
rect 31205 34527 31263 34533
rect 31205 34524 31217 34527
rect 29696 34496 31217 34524
rect 29696 34484 29702 34496
rect 31205 34493 31217 34496
rect 31251 34524 31263 34527
rect 31478 34524 31484 34536
rect 31251 34496 31484 34524
rect 31251 34493 31263 34496
rect 31205 34487 31263 34493
rect 31478 34484 31484 34496
rect 31536 34484 31542 34536
rect 33318 34484 33324 34536
rect 33376 34524 33382 34536
rect 33980 34524 34008 34555
rect 33376 34496 34008 34524
rect 33376 34484 33382 34496
rect 34256 34468 34284 34555
rect 19429 34459 19487 34465
rect 19429 34425 19441 34459
rect 19475 34425 19487 34459
rect 19429 34419 19487 34425
rect 34238 34416 34244 34468
rect 34296 34416 34302 34468
rect 3142 34348 3148 34400
rect 3200 34388 3206 34400
rect 4341 34391 4399 34397
rect 4341 34388 4353 34391
rect 3200 34360 4353 34388
rect 3200 34348 3206 34360
rect 4341 34357 4353 34360
rect 4387 34357 4399 34391
rect 4341 34351 4399 34357
rect 10594 34348 10600 34400
rect 10652 34388 10658 34400
rect 11609 34391 11667 34397
rect 11609 34388 11621 34391
rect 10652 34360 11621 34388
rect 10652 34348 10658 34360
rect 11609 34357 11621 34360
rect 11655 34388 11667 34391
rect 15930 34388 15936 34400
rect 11655 34360 15936 34388
rect 11655 34357 11667 34360
rect 11609 34351 11667 34357
rect 15930 34348 15936 34360
rect 15988 34388 15994 34400
rect 16761 34391 16819 34397
rect 16761 34388 16773 34391
rect 15988 34360 16773 34388
rect 15988 34348 15994 34360
rect 16761 34357 16773 34360
rect 16807 34388 16819 34391
rect 17218 34388 17224 34400
rect 16807 34360 17224 34388
rect 16807 34357 16819 34360
rect 16761 34351 16819 34357
rect 17218 34348 17224 34360
rect 17276 34348 17282 34400
rect 34054 34348 34060 34400
rect 34112 34388 34118 34400
rect 34348 34388 34376 34555
rect 34609 34527 34667 34533
rect 34609 34493 34621 34527
rect 34655 34524 34667 34527
rect 35894 34524 35900 34536
rect 34655 34496 35900 34524
rect 34655 34493 34667 34496
rect 34609 34487 34667 34493
rect 35894 34484 35900 34496
rect 35952 34484 35958 34536
rect 34112 34360 34376 34388
rect 34112 34348 34118 34360
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 2593 34187 2651 34193
rect 2593 34153 2605 34187
rect 2639 34184 2651 34187
rect 2774 34184 2780 34196
rect 2639 34156 2780 34184
rect 2639 34153 2651 34156
rect 2593 34147 2651 34153
rect 2774 34144 2780 34156
rect 2832 34144 2838 34196
rect 4062 34144 4068 34196
rect 4120 34184 4126 34196
rect 5534 34184 5540 34196
rect 4120 34156 5540 34184
rect 4120 34144 4126 34156
rect 5534 34144 5540 34156
rect 5592 34144 5598 34196
rect 7377 34187 7435 34193
rect 7377 34153 7389 34187
rect 7423 34184 7435 34187
rect 7466 34184 7472 34196
rect 7423 34156 7472 34184
rect 7423 34153 7435 34156
rect 7377 34147 7435 34153
rect 7466 34144 7472 34156
rect 7524 34144 7530 34196
rect 10502 34144 10508 34196
rect 10560 34184 10566 34196
rect 19242 34184 19248 34196
rect 10560 34156 19248 34184
rect 10560 34144 10566 34156
rect 19242 34144 19248 34156
rect 19300 34144 19306 34196
rect 20349 34187 20407 34193
rect 20349 34153 20361 34187
rect 20395 34184 20407 34187
rect 20714 34184 20720 34196
rect 20395 34156 20720 34184
rect 20395 34153 20407 34156
rect 20349 34147 20407 34153
rect 20714 34144 20720 34156
rect 20772 34144 20778 34196
rect 24302 34144 24308 34196
rect 24360 34184 24366 34196
rect 24397 34187 24455 34193
rect 24397 34184 24409 34187
rect 24360 34156 24409 34184
rect 24360 34144 24366 34156
rect 24397 34153 24409 34156
rect 24443 34153 24455 34187
rect 24397 34147 24455 34153
rect 24486 34144 24492 34196
rect 24544 34184 24550 34196
rect 33045 34187 33103 34193
rect 33045 34184 33057 34187
rect 24544 34156 33057 34184
rect 24544 34144 24550 34156
rect 33045 34153 33057 34156
rect 33091 34184 33103 34187
rect 36262 34184 36268 34196
rect 33091 34156 36268 34184
rect 33091 34153 33103 34156
rect 33045 34147 33103 34153
rect 3252 34088 4752 34116
rect 2866 33980 2872 33992
rect 2746 33952 2872 33980
rect 2133 33915 2191 33921
rect 2133 33881 2145 33915
rect 2179 33912 2191 33915
rect 2746 33912 2774 33952
rect 2866 33940 2872 33952
rect 2924 33940 2930 33992
rect 2961 33983 3019 33989
rect 2961 33949 2973 33983
rect 3007 33949 3019 33983
rect 2961 33943 3019 33949
rect 3053 33983 3111 33989
rect 3053 33949 3065 33983
rect 3099 33980 3111 33983
rect 3142 33980 3148 33992
rect 3099 33952 3148 33980
rect 3099 33949 3111 33952
rect 3053 33943 3111 33949
rect 2179 33884 2774 33912
rect 2976 33912 3004 33943
rect 3142 33940 3148 33952
rect 3200 33940 3206 33992
rect 3252 33989 3280 34088
rect 3237 33983 3295 33989
rect 3237 33949 3249 33983
rect 3283 33949 3295 33983
rect 4062 33980 4068 33992
rect 4023 33952 4068 33980
rect 3237 33943 3295 33949
rect 4062 33940 4068 33952
rect 4120 33940 4126 33992
rect 4157 33983 4215 33989
rect 4157 33949 4169 33983
rect 4203 33949 4215 33983
rect 4157 33943 4215 33949
rect 4249 33983 4307 33989
rect 4249 33949 4261 33983
rect 4295 33980 4307 33983
rect 4338 33980 4344 33992
rect 4295 33952 4344 33980
rect 4295 33949 4307 33952
rect 4249 33943 4307 33949
rect 4172 33912 4200 33943
rect 4338 33940 4344 33952
rect 4396 33940 4402 33992
rect 4433 33983 4491 33989
rect 4433 33949 4445 33983
rect 4479 33980 4491 33983
rect 4724 33980 4752 34088
rect 7282 34076 7288 34128
rect 7340 34116 7346 34128
rect 7837 34119 7895 34125
rect 7837 34116 7849 34119
rect 7340 34088 7849 34116
rect 7340 34076 7346 34088
rect 7837 34085 7849 34088
rect 7883 34116 7895 34119
rect 7926 34116 7932 34128
rect 7883 34088 7932 34116
rect 7883 34085 7895 34088
rect 7837 34079 7895 34085
rect 7926 34076 7932 34088
rect 7984 34116 7990 34128
rect 29733 34119 29791 34125
rect 29733 34116 29745 34119
rect 7984 34088 29745 34116
rect 7984 34076 7990 34088
rect 29733 34085 29745 34088
rect 29779 34085 29791 34119
rect 29733 34079 29791 34085
rect 7558 34048 7564 34060
rect 7208 34020 7564 34048
rect 5166 33980 5172 33992
rect 4479 33952 5172 33980
rect 4479 33949 4491 33952
rect 4433 33943 4491 33949
rect 5166 33940 5172 33952
rect 5224 33940 5230 33992
rect 5534 33980 5540 33992
rect 5495 33952 5540 33980
rect 5534 33940 5540 33952
rect 5592 33940 5598 33992
rect 7208 33989 7236 34020
rect 7558 34008 7564 34020
rect 7616 34048 7622 34060
rect 14369 34051 14427 34057
rect 7616 34020 9352 34048
rect 7616 34008 7622 34020
rect 7193 33983 7251 33989
rect 7193 33949 7205 33983
rect 7239 33949 7251 33983
rect 8938 33980 8944 33992
rect 8899 33952 8944 33980
rect 7193 33943 7251 33949
rect 8938 33940 8944 33952
rect 8996 33940 9002 33992
rect 9030 33940 9036 33992
rect 9088 33980 9094 33992
rect 9324 33989 9352 34020
rect 14369 34017 14381 34051
rect 14415 34048 14427 34051
rect 15194 34048 15200 34060
rect 14415 34020 15200 34048
rect 14415 34017 14427 34020
rect 14369 34011 14427 34017
rect 15194 34008 15200 34020
rect 15252 34048 15258 34060
rect 16761 34051 16819 34057
rect 16761 34048 16773 34051
rect 15252 34020 16068 34048
rect 15252 34008 15258 34020
rect 9309 33983 9367 33989
rect 9088 33952 9133 33980
rect 9088 33940 9094 33952
rect 9309 33949 9321 33983
rect 9355 33949 9367 33983
rect 9309 33943 9367 33949
rect 9447 33983 9505 33989
rect 9447 33949 9459 33983
rect 9493 33980 9505 33983
rect 13630 33980 13636 33992
rect 9493 33952 13636 33980
rect 9493 33949 9505 33952
rect 9447 33943 9505 33949
rect 13630 33940 13636 33952
rect 13688 33940 13694 33992
rect 13814 33940 13820 33992
rect 13872 33980 13878 33992
rect 14093 33983 14151 33989
rect 14093 33980 14105 33983
rect 13872 33952 14105 33980
rect 13872 33940 13878 33952
rect 14093 33949 14105 33952
rect 14139 33949 14151 33983
rect 15930 33980 15936 33992
rect 15891 33952 15936 33980
rect 14093 33943 14151 33949
rect 15930 33940 15936 33952
rect 15988 33940 15994 33992
rect 16040 33989 16068 34020
rect 16132 34020 16773 34048
rect 16132 33989 16160 34020
rect 16761 34017 16773 34020
rect 16807 34017 16819 34051
rect 26234 34048 26240 34060
rect 16761 34011 16819 34017
rect 24872 34020 26240 34048
rect 16025 33983 16083 33989
rect 16025 33949 16037 33983
rect 16071 33949 16083 33983
rect 16025 33943 16083 33949
rect 16117 33983 16175 33989
rect 16117 33949 16129 33983
rect 16163 33949 16175 33983
rect 16117 33943 16175 33949
rect 16301 33983 16359 33989
rect 16301 33949 16313 33983
rect 16347 33949 16359 33983
rect 16301 33943 16359 33949
rect 5258 33912 5264 33924
rect 2976 33884 5264 33912
rect 2179 33881 2191 33884
rect 2133 33875 2191 33881
rect 2746 33844 2774 33884
rect 5258 33872 5264 33884
rect 5316 33872 5322 33924
rect 7009 33915 7067 33921
rect 7009 33881 7021 33915
rect 7055 33912 7067 33915
rect 7558 33912 7564 33924
rect 7055 33884 7564 33912
rect 7055 33881 7067 33884
rect 7009 33875 7067 33881
rect 7558 33872 7564 33884
rect 7616 33872 7622 33924
rect 9214 33912 9220 33924
rect 9175 33884 9220 33912
rect 9214 33872 9220 33884
rect 9272 33872 9278 33924
rect 15470 33872 15476 33924
rect 15528 33912 15534 33924
rect 16316 33912 16344 33943
rect 16574 33940 16580 33992
rect 16632 33980 16638 33992
rect 17129 33983 17187 33989
rect 17129 33980 17141 33983
rect 16632 33952 17141 33980
rect 16632 33940 16638 33952
rect 17129 33949 17141 33952
rect 17175 33980 17187 33983
rect 17678 33980 17684 33992
rect 17175 33952 17684 33980
rect 17175 33949 17187 33952
rect 17129 33943 17187 33949
rect 17678 33940 17684 33952
rect 17736 33940 17742 33992
rect 18693 33983 18751 33989
rect 18693 33949 18705 33983
rect 18739 33980 18751 33983
rect 19242 33980 19248 33992
rect 18739 33952 19248 33980
rect 18739 33949 18751 33952
rect 18693 33943 18751 33949
rect 19242 33940 19248 33952
rect 19300 33980 19306 33992
rect 19705 33983 19763 33989
rect 19705 33980 19717 33983
rect 19300 33952 19717 33980
rect 19300 33940 19306 33952
rect 19705 33949 19717 33952
rect 19751 33949 19763 33983
rect 19886 33980 19892 33992
rect 19847 33952 19892 33980
rect 19705 33943 19763 33949
rect 19886 33940 19892 33952
rect 19944 33940 19950 33992
rect 19978 33940 19984 33992
rect 20036 33980 20042 33992
rect 20119 33983 20177 33989
rect 20036 33952 20081 33980
rect 20036 33940 20042 33952
rect 20119 33949 20131 33983
rect 20165 33980 20177 33983
rect 20346 33980 20352 33992
rect 20165 33952 20352 33980
rect 20165 33949 20177 33952
rect 20119 33943 20177 33949
rect 20346 33940 20352 33952
rect 20404 33980 20410 33992
rect 20809 33983 20867 33989
rect 20809 33980 20821 33983
rect 20404 33952 20821 33980
rect 20404 33940 20410 33952
rect 20809 33949 20821 33952
rect 20855 33949 20867 33983
rect 20809 33943 20867 33949
rect 23753 33983 23811 33989
rect 23753 33949 23765 33983
rect 23799 33980 23811 33983
rect 24118 33980 24124 33992
rect 23799 33952 24124 33980
rect 23799 33949 23811 33952
rect 23753 33943 23811 33949
rect 24118 33940 24124 33952
rect 24176 33980 24182 33992
rect 24394 33980 24400 33992
rect 24176 33952 24400 33980
rect 24176 33940 24182 33952
rect 24394 33940 24400 33952
rect 24452 33980 24458 33992
rect 24627 33983 24685 33989
rect 24627 33980 24639 33983
rect 24452 33952 24639 33980
rect 24452 33940 24458 33952
rect 24627 33949 24639 33952
rect 24673 33949 24685 33983
rect 24762 33980 24768 33992
rect 24723 33952 24768 33980
rect 24627 33943 24685 33949
rect 24762 33940 24768 33952
rect 24820 33940 24826 33992
rect 24872 33989 24900 34020
rect 26234 34008 26240 34020
rect 26292 34008 26298 34060
rect 27062 34008 27068 34060
rect 27120 34048 27126 34060
rect 27120 34020 27936 34048
rect 27120 34008 27126 34020
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33949 24915 33983
rect 24857 33943 24915 33949
rect 25041 33983 25099 33989
rect 25041 33949 25053 33983
rect 25087 33980 25099 33983
rect 25130 33980 25136 33992
rect 25087 33952 25136 33980
rect 25087 33949 25099 33952
rect 25041 33943 25099 33949
rect 15528 33884 16344 33912
rect 15528 33872 15534 33884
rect 16132 33856 16160 33884
rect 16850 33872 16856 33924
rect 16908 33912 16914 33924
rect 16945 33915 17003 33921
rect 16945 33912 16957 33915
rect 16908 33884 16957 33912
rect 16908 33872 16914 33884
rect 16945 33881 16957 33884
rect 16991 33881 17003 33915
rect 16945 33875 17003 33881
rect 17957 33915 18015 33921
rect 17957 33881 17969 33915
rect 18003 33912 18015 33915
rect 18506 33912 18512 33924
rect 18003 33884 18512 33912
rect 18003 33881 18015 33884
rect 17957 33875 18015 33881
rect 18506 33872 18512 33884
rect 18564 33872 18570 33924
rect 23842 33872 23848 33924
rect 23900 33912 23906 33924
rect 25056 33912 25084 33943
rect 25130 33940 25136 33952
rect 25188 33940 25194 33992
rect 26694 33980 26700 33992
rect 26655 33952 26700 33980
rect 26694 33940 26700 33952
rect 26752 33980 26758 33992
rect 27338 33980 27344 33992
rect 26752 33952 27344 33980
rect 26752 33940 26758 33952
rect 27338 33940 27344 33952
rect 27396 33980 27402 33992
rect 27525 33983 27583 33989
rect 27525 33980 27537 33983
rect 27396 33952 27537 33980
rect 27396 33940 27402 33952
rect 27525 33949 27537 33952
rect 27571 33949 27583 33983
rect 27525 33943 27583 33949
rect 27614 33977 27672 33983
rect 27614 33943 27626 33977
rect 27660 33943 27672 33977
rect 27614 33937 27672 33943
rect 27706 33940 27712 33992
rect 27764 33989 27770 33992
rect 27908 33989 27936 34020
rect 27764 33980 27772 33989
rect 27893 33983 27951 33989
rect 27764 33952 27809 33980
rect 27764 33943 27772 33952
rect 27893 33949 27905 33983
rect 27939 33949 27951 33983
rect 29748 33980 29776 34079
rect 31757 34051 31815 34057
rect 31757 34048 31769 34051
rect 30760 34020 31769 34048
rect 30006 33980 30012 33992
rect 29748 33952 30012 33980
rect 27893 33943 27951 33949
rect 27764 33940 27770 33943
rect 30006 33940 30012 33952
rect 30064 33980 30070 33992
rect 30515 33983 30573 33989
rect 30515 33980 30527 33983
rect 30064 33952 30527 33980
rect 30064 33940 30070 33952
rect 30515 33949 30527 33952
rect 30561 33949 30573 33983
rect 30650 33980 30656 33992
rect 30611 33952 30656 33980
rect 30515 33943 30573 33949
rect 30650 33940 30656 33952
rect 30708 33940 30714 33992
rect 30760 33989 30788 34020
rect 31757 34017 31769 34020
rect 31803 34017 31815 34051
rect 31757 34011 31815 34017
rect 30745 33983 30803 33989
rect 30745 33949 30757 33983
rect 30791 33949 30803 33983
rect 30926 33980 30932 33992
rect 30887 33952 30932 33980
rect 30745 33943 30803 33949
rect 30926 33940 30932 33952
rect 30984 33940 30990 33992
rect 33318 33940 33324 33992
rect 33376 33980 33382 33992
rect 33505 33983 33563 33989
rect 33505 33980 33517 33983
rect 33376 33952 33517 33980
rect 33376 33940 33382 33952
rect 33505 33949 33517 33952
rect 33551 33949 33563 33983
rect 33686 33980 33692 33992
rect 33647 33952 33692 33980
rect 33505 33943 33563 33949
rect 33686 33940 33692 33952
rect 33744 33940 33750 33992
rect 33888 33989 33916 34156
rect 36262 34144 36268 34156
rect 36320 34144 36326 34196
rect 33781 33983 33839 33989
rect 33781 33949 33793 33983
rect 33827 33949 33839 33983
rect 33781 33943 33839 33949
rect 33873 33983 33931 33989
rect 33873 33949 33885 33983
rect 33919 33949 33931 33983
rect 34238 33980 34244 33992
rect 33873 33943 33931 33949
rect 33980 33952 34244 33980
rect 23900 33884 25084 33912
rect 23900 33872 23906 33884
rect 27632 33856 27660 33937
rect 29546 33872 29552 33924
rect 29604 33912 29610 33924
rect 31389 33915 31447 33921
rect 31389 33912 31401 33915
rect 29604 33884 31401 33912
rect 29604 33872 29610 33884
rect 31389 33881 31401 33884
rect 31435 33881 31447 33915
rect 31570 33912 31576 33924
rect 31531 33884 31576 33912
rect 31389 33875 31447 33881
rect 31570 33872 31576 33884
rect 31628 33872 31634 33924
rect 33226 33872 33232 33924
rect 33284 33912 33290 33924
rect 33796 33912 33824 33943
rect 33980 33912 34008 33952
rect 34238 33940 34244 33952
rect 34296 33940 34302 33992
rect 34422 33940 34428 33992
rect 34480 33980 34486 33992
rect 36081 33983 36139 33989
rect 34480 33952 36032 33980
rect 34480 33940 34486 33952
rect 33284 33884 34008 33912
rect 34149 33915 34207 33921
rect 33284 33872 33290 33884
rect 34149 33881 34161 33915
rect 34195 33912 34207 33915
rect 35814 33915 35872 33921
rect 35814 33912 35826 33915
rect 34195 33884 35826 33912
rect 34195 33881 34207 33884
rect 34149 33875 34207 33881
rect 35814 33881 35826 33884
rect 35860 33881 35872 33915
rect 36004 33912 36032 33952
rect 36081 33949 36093 33983
rect 36127 33980 36139 33983
rect 36170 33980 36176 33992
rect 36127 33952 36176 33980
rect 36127 33949 36139 33952
rect 36081 33943 36139 33949
rect 36170 33940 36176 33952
rect 36228 33980 36234 33992
rect 36722 33980 36728 33992
rect 36228 33952 36728 33980
rect 36228 33940 36234 33952
rect 36722 33940 36728 33952
rect 36780 33980 36786 33992
rect 38473 33983 38531 33989
rect 38473 33980 38485 33983
rect 36780 33952 38485 33980
rect 36780 33940 36786 33952
rect 38473 33949 38485 33952
rect 38519 33949 38531 33983
rect 38473 33943 38531 33949
rect 36909 33915 36967 33921
rect 36909 33912 36921 33915
rect 36004 33884 36921 33912
rect 35814 33875 35872 33881
rect 36909 33881 36921 33884
rect 36955 33912 36967 33915
rect 37274 33912 37280 33924
rect 36955 33884 37280 33912
rect 36955 33881 36967 33884
rect 36909 33875 36967 33881
rect 37274 33872 37280 33884
rect 37332 33872 37338 33924
rect 3234 33844 3240 33856
rect 2746 33816 3240 33844
rect 3234 33804 3240 33816
rect 3292 33804 3298 33856
rect 3786 33844 3792 33856
rect 3747 33816 3792 33844
rect 3786 33804 3792 33816
rect 3844 33804 3850 33856
rect 4985 33847 5043 33853
rect 4985 33813 4997 33847
rect 5031 33844 5043 33847
rect 5166 33844 5172 33856
rect 5031 33816 5172 33844
rect 5031 33813 5043 33816
rect 4985 33807 5043 33813
rect 5166 33804 5172 33816
rect 5224 33804 5230 33856
rect 8846 33804 8852 33856
rect 8904 33844 8910 33856
rect 9585 33847 9643 33853
rect 9585 33844 9597 33847
rect 8904 33816 9597 33844
rect 8904 33804 8910 33816
rect 9585 33813 9597 33816
rect 9631 33813 9643 33847
rect 11146 33844 11152 33856
rect 11107 33816 11152 33844
rect 9585 33807 9643 33813
rect 11146 33804 11152 33816
rect 11204 33804 11210 33856
rect 15654 33844 15660 33856
rect 15615 33816 15660 33844
rect 15654 33804 15660 33816
rect 15712 33804 15718 33856
rect 16114 33804 16120 33856
rect 16172 33804 16178 33856
rect 27246 33844 27252 33856
rect 27207 33816 27252 33844
rect 27246 33804 27252 33816
rect 27304 33804 27310 33856
rect 27614 33804 27620 33856
rect 27672 33804 27678 33856
rect 30282 33844 30288 33856
rect 30243 33816 30288 33844
rect 30282 33804 30288 33816
rect 30340 33804 30346 33856
rect 33962 33804 33968 33856
rect 34020 33844 34026 33856
rect 34701 33847 34759 33853
rect 34701 33844 34713 33847
rect 34020 33816 34713 33844
rect 34020 33804 34026 33816
rect 34701 33813 34713 33816
rect 34747 33813 34759 33847
rect 34701 33807 34759 33813
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 4338 33640 4344 33652
rect 4299 33612 4344 33640
rect 4338 33600 4344 33612
rect 4396 33600 4402 33652
rect 6730 33640 6736 33652
rect 6691 33612 6736 33640
rect 6730 33600 6736 33612
rect 6788 33600 6794 33652
rect 9214 33600 9220 33652
rect 9272 33640 9278 33652
rect 12618 33640 12624 33652
rect 9272 33612 12624 33640
rect 9272 33600 9278 33612
rect 12618 33600 12624 33612
rect 12676 33600 12682 33652
rect 13630 33600 13636 33652
rect 13688 33640 13694 33652
rect 15197 33643 15255 33649
rect 15197 33640 15209 33643
rect 13688 33612 15209 33640
rect 13688 33600 13694 33612
rect 15197 33609 15209 33612
rect 15243 33640 15255 33643
rect 19150 33640 19156 33652
rect 15243 33612 19156 33640
rect 15243 33609 15255 33612
rect 15197 33603 15255 33609
rect 19150 33600 19156 33612
rect 19208 33600 19214 33652
rect 19242 33600 19248 33652
rect 19300 33640 19306 33652
rect 19705 33643 19763 33649
rect 19705 33640 19717 33643
rect 19300 33612 19717 33640
rect 19300 33600 19306 33612
rect 19705 33609 19717 33612
rect 19751 33609 19763 33643
rect 29822 33640 29828 33652
rect 19705 33603 19763 33609
rect 22066 33612 29828 33640
rect 2768 33575 2826 33581
rect 2768 33541 2780 33575
rect 2814 33572 2826 33575
rect 3786 33572 3792 33584
rect 2814 33544 3792 33572
rect 2814 33541 2826 33544
rect 2768 33535 2826 33541
rect 3786 33532 3792 33544
rect 3844 33532 3850 33584
rect 5166 33532 5172 33584
rect 5224 33572 5230 33584
rect 6454 33572 6460 33584
rect 5224 33544 6460 33572
rect 5224 33532 5230 33544
rect 6454 33532 6460 33544
rect 6512 33572 6518 33584
rect 14458 33572 14464 33584
rect 6512 33544 14464 33572
rect 6512 33532 6518 33544
rect 14458 33532 14464 33544
rect 14516 33532 14522 33584
rect 17037 33575 17095 33581
rect 17037 33541 17049 33575
rect 17083 33572 17095 33575
rect 17083 33544 17356 33572
rect 17083 33541 17095 33544
rect 17037 33535 17095 33541
rect 4525 33507 4583 33513
rect 4525 33504 4537 33507
rect 3896 33476 4537 33504
rect 2406 33396 2412 33448
rect 2464 33436 2470 33448
rect 2501 33439 2559 33445
rect 2501 33436 2513 33439
rect 2464 33408 2513 33436
rect 2464 33396 2470 33408
rect 2501 33405 2513 33408
rect 2547 33405 2559 33439
rect 2501 33399 2559 33405
rect 3896 33377 3924 33476
rect 4525 33473 4537 33476
rect 4571 33504 4583 33507
rect 4614 33504 4620 33516
rect 4571 33476 4620 33504
rect 4571 33473 4583 33476
rect 4525 33467 4583 33473
rect 4614 33464 4620 33476
rect 4672 33464 4678 33516
rect 4706 33464 4712 33516
rect 4764 33504 4770 33516
rect 7558 33504 7564 33516
rect 4764 33476 7564 33504
rect 4764 33464 4770 33476
rect 7558 33464 7564 33476
rect 7616 33464 7622 33516
rect 12713 33507 12771 33513
rect 12713 33473 12725 33507
rect 12759 33473 12771 33507
rect 13262 33504 13268 33516
rect 13223 33476 13268 33504
rect 12713 33467 12771 33473
rect 3881 33371 3939 33377
rect 3881 33337 3893 33371
rect 3927 33337 3939 33371
rect 3881 33331 3939 33337
rect 7929 33303 7987 33309
rect 7929 33269 7941 33303
rect 7975 33300 7987 33303
rect 8110 33300 8116 33312
rect 7975 33272 8116 33300
rect 7975 33269 7987 33272
rect 7929 33263 7987 33269
rect 8110 33260 8116 33272
rect 8168 33260 8174 33312
rect 12728 33300 12756 33467
rect 13262 33464 13268 33476
rect 13320 33464 13326 33516
rect 13538 33513 13544 33516
rect 13532 33467 13544 33513
rect 13596 33504 13602 33516
rect 13596 33476 13632 33504
rect 13538 33464 13544 33467
rect 13596 33464 13602 33476
rect 15194 33464 15200 33516
rect 15252 33504 15258 33516
rect 15289 33507 15347 33513
rect 15289 33504 15301 33507
rect 15252 33476 15301 33504
rect 15252 33464 15258 33476
rect 15289 33473 15301 33476
rect 15335 33473 15347 33507
rect 16666 33504 16672 33516
rect 16627 33476 16672 33504
rect 15289 33467 15347 33473
rect 16666 33464 16672 33476
rect 16724 33464 16730 33516
rect 16850 33513 16856 33516
rect 16817 33507 16856 33513
rect 16817 33473 16829 33507
rect 16817 33467 16856 33473
rect 16850 33464 16856 33467
rect 16908 33464 16914 33516
rect 16945 33507 17003 33513
rect 16945 33473 16957 33507
rect 16991 33473 17003 33507
rect 17153 33507 17211 33513
rect 17153 33504 17165 33507
rect 16945 33467 17003 33473
rect 17144 33473 17165 33504
rect 17199 33473 17211 33507
rect 17328 33504 17356 33544
rect 17402 33532 17408 33584
rect 17460 33572 17466 33584
rect 22066 33572 22094 33612
rect 29822 33600 29828 33612
rect 29880 33640 29886 33652
rect 30193 33643 30251 33649
rect 30193 33640 30205 33643
rect 29880 33612 30205 33640
rect 29880 33600 29886 33612
rect 30193 33609 30205 33612
rect 30239 33609 30251 33643
rect 30193 33603 30251 33609
rect 33686 33600 33692 33652
rect 33744 33640 33750 33652
rect 34057 33643 34115 33649
rect 34057 33640 34069 33643
rect 33744 33612 34069 33640
rect 33744 33600 33750 33612
rect 34057 33609 34069 33612
rect 34103 33609 34115 33643
rect 34790 33640 34796 33652
rect 34751 33612 34796 33640
rect 34057 33603 34115 33609
rect 34790 33600 34796 33612
rect 34848 33600 34854 33652
rect 17460 33544 22094 33572
rect 17460 33532 17466 33544
rect 24762 33532 24768 33584
rect 24820 33572 24826 33584
rect 24820 33544 24992 33572
rect 24820 33532 24826 33544
rect 18509 33507 18567 33513
rect 18509 33504 18521 33507
rect 17328 33476 18521 33504
rect 17144 33467 17211 33473
rect 18509 33473 18521 33476
rect 18555 33473 18567 33507
rect 18690 33504 18696 33516
rect 18651 33476 18696 33504
rect 18509 33467 18567 33473
rect 16960 33436 16988 33467
rect 14292 33408 16988 33436
rect 14292 33300 14320 33408
rect 15194 33328 15200 33380
rect 15252 33368 15258 33380
rect 17144 33368 17172 33467
rect 18524 33436 18552 33467
rect 18690 33464 18696 33476
rect 18748 33464 18754 33516
rect 24578 33464 24584 33516
rect 24636 33504 24642 33516
rect 24673 33507 24731 33513
rect 24673 33504 24685 33507
rect 24636 33476 24685 33504
rect 24636 33464 24642 33476
rect 24673 33473 24685 33476
rect 24719 33473 24731 33507
rect 24854 33504 24860 33516
rect 24815 33476 24860 33504
rect 24673 33467 24731 33473
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 24964 33513 24992 33544
rect 27246 33532 27252 33584
rect 27304 33572 27310 33584
rect 27402 33575 27460 33581
rect 27402 33572 27414 33575
rect 27304 33544 27414 33572
rect 27304 33532 27310 33544
rect 27402 33541 27414 33544
rect 27448 33541 27460 33575
rect 27402 33535 27460 33541
rect 35894 33532 35900 33584
rect 35952 33581 35958 33584
rect 35952 33572 35964 33581
rect 35952 33544 35997 33572
rect 35952 33535 35964 33544
rect 35952 33532 35958 33535
rect 24949 33507 25007 33513
rect 24949 33473 24961 33507
rect 24995 33473 25007 33507
rect 24949 33467 25007 33473
rect 25041 33507 25099 33513
rect 25041 33473 25053 33507
rect 25087 33504 25099 33507
rect 25498 33504 25504 33516
rect 25087 33476 25504 33504
rect 25087 33473 25099 33476
rect 25041 33467 25099 33473
rect 20622 33436 20628 33448
rect 18524 33408 20628 33436
rect 20622 33396 20628 33408
rect 20680 33396 20686 33448
rect 25056 33436 25084 33467
rect 25498 33464 25504 33476
rect 25556 33464 25562 33516
rect 29638 33464 29644 33516
rect 29696 33504 29702 33516
rect 30009 33507 30067 33513
rect 30009 33504 30021 33507
rect 29696 33476 30021 33504
rect 29696 33464 29702 33476
rect 30009 33473 30021 33476
rect 30055 33473 30067 33507
rect 30009 33467 30067 33473
rect 33410 33464 33416 33516
rect 33468 33504 33474 33516
rect 33689 33507 33747 33513
rect 33689 33504 33701 33507
rect 33468 33476 33701 33504
rect 33468 33464 33474 33476
rect 33689 33473 33701 33476
rect 33735 33473 33747 33507
rect 33689 33467 33747 33473
rect 33873 33507 33931 33513
rect 33873 33473 33885 33507
rect 33919 33504 33931 33507
rect 33962 33504 33968 33516
rect 33919 33476 33968 33504
rect 33919 33473 33931 33476
rect 33873 33467 33931 33473
rect 33962 33464 33968 33476
rect 34020 33464 34026 33516
rect 27154 33436 27160 33448
rect 22066 33408 25084 33436
rect 27115 33408 27160 33436
rect 15252 33340 17172 33368
rect 15252 33328 15258 33340
rect 20346 33328 20352 33380
rect 20404 33368 20410 33380
rect 22066 33368 22094 33408
rect 27154 33396 27160 33408
rect 27212 33396 27218 33448
rect 30558 33396 30564 33448
rect 30616 33436 30622 33448
rect 32401 33439 32459 33445
rect 32401 33436 32413 33439
rect 30616 33408 32413 33436
rect 30616 33396 30622 33408
rect 32401 33405 32413 33408
rect 32447 33405 32459 33439
rect 32401 33399 32459 33405
rect 32677 33439 32735 33445
rect 32677 33405 32689 33439
rect 32723 33436 32735 33439
rect 33226 33436 33232 33448
rect 32723 33408 33232 33436
rect 32723 33405 32735 33408
rect 32677 33399 32735 33405
rect 20404 33340 22094 33368
rect 32416 33368 32444 33399
rect 33226 33396 33232 33408
rect 33284 33396 33290 33448
rect 36170 33436 36176 33448
rect 36131 33408 36176 33436
rect 36170 33396 36176 33408
rect 36228 33396 36234 33448
rect 32950 33368 32956 33380
rect 32416 33340 32956 33368
rect 20404 33328 20410 33340
rect 32950 33328 32956 33340
rect 33008 33328 33014 33380
rect 58158 33368 58164 33380
rect 58119 33340 58164 33368
rect 58158 33328 58164 33340
rect 58216 33328 58222 33380
rect 14366 33300 14372 33312
rect 12728 33272 14372 33300
rect 14366 33260 14372 33272
rect 14424 33260 14430 33312
rect 14642 33300 14648 33312
rect 14603 33272 14648 33300
rect 14642 33260 14648 33272
rect 14700 33260 14706 33312
rect 17310 33300 17316 33312
rect 17271 33272 17316 33300
rect 17310 33260 17316 33272
rect 17368 33260 17374 33312
rect 18230 33260 18236 33312
rect 18288 33300 18294 33312
rect 18325 33303 18383 33309
rect 18325 33300 18337 33303
rect 18288 33272 18337 33300
rect 18288 33260 18294 33272
rect 18325 33269 18337 33272
rect 18371 33269 18383 33303
rect 19242 33300 19248 33312
rect 19203 33272 19248 33300
rect 18325 33263 18383 33269
rect 19242 33260 19248 33272
rect 19300 33260 19306 33312
rect 23842 33260 23848 33312
rect 23900 33300 23906 33312
rect 24029 33303 24087 33309
rect 24029 33300 24041 33303
rect 23900 33272 24041 33300
rect 23900 33260 23906 33272
rect 24029 33269 24041 33272
rect 24075 33269 24087 33303
rect 25314 33300 25320 33312
rect 25275 33272 25320 33300
rect 24029 33263 24087 33269
rect 25314 33260 25320 33272
rect 25372 33260 25378 33312
rect 25498 33260 25504 33312
rect 25556 33300 25562 33312
rect 25777 33303 25835 33309
rect 25777 33300 25789 33303
rect 25556 33272 25789 33300
rect 25556 33260 25562 33272
rect 25777 33269 25789 33272
rect 25823 33269 25835 33303
rect 28534 33300 28540 33312
rect 28495 33272 28540 33300
rect 25777 33263 25835 33269
rect 28534 33260 28540 33272
rect 28592 33260 28598 33312
rect 29549 33303 29607 33309
rect 29549 33269 29561 33303
rect 29595 33300 29607 33303
rect 29638 33300 29644 33312
rect 29595 33272 29644 33300
rect 29595 33269 29607 33272
rect 29549 33263 29607 33269
rect 29638 33260 29644 33272
rect 29696 33260 29702 33312
rect 30926 33260 30932 33312
rect 30984 33300 30990 33312
rect 35986 33300 35992 33312
rect 30984 33272 35992 33300
rect 30984 33260 30990 33272
rect 35986 33260 35992 33272
rect 36044 33260 36050 33312
rect 37274 33300 37280 33312
rect 37235 33272 37280 33300
rect 37274 33260 37280 33272
rect 37332 33260 37338 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 3881 33099 3939 33105
rect 3881 33065 3893 33099
rect 3927 33096 3939 33099
rect 5166 33096 5172 33108
rect 3927 33068 5172 33096
rect 3927 33065 3939 33068
rect 3881 33059 3939 33065
rect 5166 33056 5172 33068
rect 5224 33056 5230 33108
rect 5258 33056 5264 33108
rect 5316 33096 5322 33108
rect 7190 33096 7196 33108
rect 5316 33068 7196 33096
rect 5316 33056 5322 33068
rect 7190 33056 7196 33068
rect 7248 33056 7254 33108
rect 8297 33099 8355 33105
rect 8297 33065 8309 33099
rect 8343 33096 8355 33099
rect 9950 33096 9956 33108
rect 8343 33068 9956 33096
rect 8343 33065 8355 33068
rect 8297 33059 8355 33065
rect 8110 32960 8116 32972
rect 7300 32932 8116 32960
rect 4893 32895 4951 32901
rect 4893 32861 4905 32895
rect 4939 32892 4951 32895
rect 6730 32892 6736 32904
rect 4939 32864 6736 32892
rect 4939 32861 4951 32864
rect 4893 32855 4951 32861
rect 6730 32852 6736 32864
rect 6788 32852 6794 32904
rect 7300 32892 7328 32932
rect 8110 32920 8116 32932
rect 8168 32920 8174 32972
rect 7374 32892 7380 32904
rect 7287 32864 7380 32892
rect 7374 32852 7380 32864
rect 7432 32852 7438 32904
rect 7469 32895 7527 32901
rect 7469 32861 7481 32895
rect 7515 32861 7527 32895
rect 7469 32855 7527 32861
rect 7561 32895 7619 32901
rect 7561 32861 7573 32895
rect 7607 32892 7619 32895
rect 7650 32892 7656 32904
rect 7607 32864 7656 32892
rect 7607 32861 7619 32864
rect 7561 32855 7619 32861
rect 6641 32827 6699 32833
rect 6641 32793 6653 32827
rect 6687 32824 6699 32827
rect 6822 32824 6828 32836
rect 6687 32796 6828 32824
rect 6687 32793 6699 32796
rect 6641 32787 6699 32793
rect 6822 32784 6828 32796
rect 6880 32784 6886 32836
rect 7484 32768 7512 32855
rect 7650 32852 7656 32864
rect 7708 32852 7714 32904
rect 7745 32895 7803 32901
rect 7745 32861 7757 32895
rect 7791 32892 7803 32895
rect 8312 32892 8340 33059
rect 9950 33056 9956 33068
rect 10008 33096 10014 33108
rect 10410 33096 10416 33108
rect 10008 33068 10416 33096
rect 10008 33056 10014 33068
rect 10410 33056 10416 33068
rect 10468 33056 10474 33108
rect 13538 33096 13544 33108
rect 13499 33068 13544 33096
rect 13538 33056 13544 33068
rect 13596 33056 13602 33108
rect 16574 33096 16580 33108
rect 14384 33068 16580 33096
rect 12710 32988 12716 33040
rect 12768 33028 12774 33040
rect 12768 33000 14320 33028
rect 12768 32988 12774 33000
rect 10410 32920 10416 32972
rect 10468 32960 10474 32972
rect 13814 32960 13820 32972
rect 10468 32932 13820 32960
rect 10468 32920 10474 32932
rect 10226 32892 10232 32904
rect 7791 32864 8340 32892
rect 10187 32864 10232 32892
rect 7791 32861 7803 32864
rect 7745 32855 7803 32861
rect 10226 32852 10232 32864
rect 10284 32892 10290 32904
rect 10870 32892 10876 32904
rect 10284 32864 10876 32892
rect 10284 32852 10290 32864
rect 10870 32852 10876 32864
rect 10928 32852 10934 32904
rect 12710 32852 12716 32904
rect 12768 32892 12774 32904
rect 12897 32895 12955 32901
rect 12897 32892 12909 32895
rect 12768 32864 12909 32892
rect 12768 32852 12774 32864
rect 12897 32861 12909 32864
rect 12943 32861 12955 32895
rect 13078 32892 13084 32904
rect 13039 32864 13084 32892
rect 12897 32855 12955 32861
rect 13078 32852 13084 32864
rect 13136 32852 13142 32904
rect 13188 32901 13216 32932
rect 13814 32920 13820 32932
rect 13872 32920 13878 32972
rect 13173 32895 13231 32901
rect 13173 32861 13185 32895
rect 13219 32861 13231 32895
rect 13173 32855 13231 32861
rect 13265 32895 13323 32901
rect 13265 32861 13277 32895
rect 13311 32861 13323 32895
rect 14090 32892 14096 32904
rect 14051 32864 14096 32892
rect 13265 32855 13323 32861
rect 12437 32827 12495 32833
rect 12437 32793 12449 32827
rect 12483 32824 12495 32827
rect 13280 32824 13308 32855
rect 14090 32852 14096 32864
rect 14148 32852 14154 32904
rect 14292 32892 14320 33000
rect 14384 32969 14412 33068
rect 16574 33056 16580 33068
rect 16632 33056 16638 33108
rect 16850 33056 16856 33108
rect 16908 33096 16914 33108
rect 16945 33099 17003 33105
rect 16945 33096 16957 33099
rect 16908 33068 16957 33096
rect 16908 33056 16914 33068
rect 16945 33065 16957 33068
rect 16991 33065 17003 33099
rect 16945 33059 17003 33065
rect 19242 33056 19248 33108
rect 19300 33096 19306 33108
rect 25222 33096 25228 33108
rect 19300 33068 25228 33096
rect 19300 33056 19306 33068
rect 25222 33056 25228 33068
rect 25280 33096 25286 33108
rect 25774 33096 25780 33108
rect 25280 33068 25780 33096
rect 25280 33056 25286 33068
rect 25774 33056 25780 33068
rect 25832 33056 25838 33108
rect 27706 33056 27712 33108
rect 27764 33096 27770 33108
rect 27801 33099 27859 33105
rect 27801 33096 27813 33099
rect 27764 33068 27813 33096
rect 27764 33056 27770 33068
rect 27801 33065 27813 33068
rect 27847 33065 27859 33099
rect 27801 33059 27859 33065
rect 31018 33056 31024 33108
rect 31076 33096 31082 33108
rect 31205 33099 31263 33105
rect 31205 33096 31217 33099
rect 31076 33068 31217 33096
rect 31076 33056 31082 33068
rect 31205 33065 31217 33068
rect 31251 33096 31263 33099
rect 31570 33096 31576 33108
rect 31251 33068 31576 33096
rect 31251 33065 31263 33068
rect 31205 33059 31263 33065
rect 31570 33056 31576 33068
rect 31628 33056 31634 33108
rect 14369 32963 14427 32969
rect 14369 32929 14381 32963
rect 14415 32929 14427 32963
rect 15470 32960 15476 32972
rect 14369 32923 14427 32929
rect 14660 32932 15476 32960
rect 14660 32892 14688 32932
rect 15470 32920 15476 32932
rect 15528 32920 15534 32972
rect 16666 32920 16672 32972
rect 16724 32960 16730 32972
rect 18138 32960 18144 32972
rect 16724 32932 18144 32960
rect 16724 32920 16730 32932
rect 14292 32864 14688 32892
rect 14734 32852 14740 32904
rect 14792 32892 14798 32904
rect 15565 32895 15623 32901
rect 15565 32892 15577 32895
rect 14792 32864 15577 32892
rect 14792 32852 14798 32864
rect 15565 32861 15577 32864
rect 15611 32892 15623 32895
rect 17126 32892 17132 32904
rect 15611 32864 17132 32892
rect 15611 32861 15623 32864
rect 15565 32855 15623 32861
rect 17126 32852 17132 32864
rect 17184 32892 17190 32904
rect 17954 32892 17960 32904
rect 17184 32864 17960 32892
rect 17184 32852 17190 32864
rect 17954 32852 17960 32864
rect 18012 32852 18018 32904
rect 18069 32901 18097 32932
rect 18138 32920 18144 32932
rect 18196 32920 18202 32972
rect 19260 32960 19288 33056
rect 20622 33028 20628 33040
rect 20583 33000 20628 33028
rect 20622 32988 20628 33000
rect 20680 32988 20686 33040
rect 18432 32932 19288 32960
rect 18055 32895 18113 32901
rect 18055 32861 18067 32895
rect 18101 32861 18113 32895
rect 18230 32892 18236 32904
rect 18191 32864 18236 32892
rect 18055 32855 18113 32861
rect 18230 32852 18236 32864
rect 18288 32852 18294 32904
rect 18432 32901 18460 32932
rect 24578 32920 24584 32972
rect 24636 32960 24642 32972
rect 24673 32963 24731 32969
rect 24673 32960 24685 32963
rect 24636 32932 24685 32960
rect 24636 32920 24642 32932
rect 24673 32929 24685 32932
rect 24719 32929 24731 32963
rect 24673 32923 24731 32929
rect 18325 32895 18383 32901
rect 18325 32861 18337 32895
rect 18371 32861 18383 32895
rect 18325 32855 18383 32861
rect 18417 32895 18475 32901
rect 18417 32861 18429 32895
rect 18463 32861 18475 32895
rect 19242 32892 19248 32904
rect 19203 32864 19248 32892
rect 18417 32855 18475 32861
rect 12483 32796 13308 32824
rect 12483 32793 12495 32796
rect 12437 32787 12495 32793
rect 12912 32768 12940 32796
rect 15654 32784 15660 32836
rect 15712 32824 15718 32836
rect 15810 32827 15868 32833
rect 15810 32824 15822 32827
rect 15712 32796 15822 32824
rect 15712 32784 15718 32796
rect 15810 32793 15822 32796
rect 15856 32793 15868 32827
rect 15810 32787 15868 32793
rect 7101 32759 7159 32765
rect 7101 32725 7113 32759
rect 7147 32756 7159 32759
rect 7190 32756 7196 32768
rect 7147 32728 7196 32756
rect 7147 32725 7159 32728
rect 7101 32719 7159 32725
rect 7190 32716 7196 32728
rect 7248 32716 7254 32768
rect 7466 32716 7472 32768
rect 7524 32716 7530 32768
rect 10134 32716 10140 32768
rect 10192 32756 10198 32768
rect 10321 32759 10379 32765
rect 10321 32756 10333 32759
rect 10192 32728 10333 32756
rect 10192 32716 10198 32728
rect 10321 32725 10333 32728
rect 10367 32725 10379 32759
rect 10321 32719 10379 32725
rect 12894 32716 12900 32768
rect 12952 32716 12958 32768
rect 17034 32716 17040 32768
rect 17092 32756 17098 32768
rect 18340 32756 18368 32855
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 24397 32895 24455 32901
rect 24397 32892 24409 32895
rect 24044 32864 24409 32892
rect 18693 32827 18751 32833
rect 18693 32793 18705 32827
rect 18739 32824 18751 32827
rect 19490 32827 19548 32833
rect 19490 32824 19502 32827
rect 18739 32796 19502 32824
rect 18739 32793 18751 32796
rect 18693 32787 18751 32793
rect 19490 32793 19502 32796
rect 19536 32793 19548 32827
rect 19490 32787 19548 32793
rect 24044 32768 24072 32864
rect 24397 32861 24409 32864
rect 24443 32861 24455 32895
rect 24397 32855 24455 32861
rect 27985 32895 28043 32901
rect 27985 32861 27997 32895
rect 28031 32892 28043 32895
rect 28534 32892 28540 32904
rect 28031 32864 28540 32892
rect 28031 32861 28043 32864
rect 27985 32855 28043 32861
rect 28534 32852 28540 32864
rect 28592 32852 28598 32904
rect 29825 32895 29883 32901
rect 29825 32861 29837 32895
rect 29871 32892 29883 32895
rect 33134 32892 33140 32904
rect 29871 32864 33140 32892
rect 29871 32861 29883 32864
rect 29825 32855 29883 32861
rect 33134 32852 33140 32864
rect 33192 32852 33198 32904
rect 28169 32827 28227 32833
rect 28169 32793 28181 32827
rect 28215 32824 28227 32827
rect 29546 32824 29552 32836
rect 28215 32796 29552 32824
rect 28215 32793 28227 32796
rect 28169 32787 28227 32793
rect 29546 32784 29552 32796
rect 29604 32824 29610 32836
rect 29914 32824 29920 32836
rect 29604 32796 29920 32824
rect 29604 32784 29610 32796
rect 29914 32784 29920 32796
rect 29972 32784 29978 32836
rect 30092 32827 30150 32833
rect 30092 32793 30104 32827
rect 30138 32824 30150 32827
rect 30282 32824 30288 32836
rect 30138 32796 30288 32824
rect 30138 32793 30150 32796
rect 30092 32787 30150 32793
rect 30282 32784 30288 32796
rect 30340 32784 30346 32836
rect 32122 32824 32128 32836
rect 32083 32796 32128 32824
rect 32122 32784 32128 32796
rect 32180 32784 32186 32836
rect 32309 32827 32367 32833
rect 32309 32793 32321 32827
rect 32355 32824 32367 32827
rect 33226 32824 33232 32836
rect 32355 32796 33232 32824
rect 32355 32793 32367 32796
rect 32309 32787 32367 32793
rect 33226 32784 33232 32796
rect 33284 32784 33290 32836
rect 19978 32756 19984 32768
rect 17092 32728 19984 32756
rect 17092 32716 17098 32728
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 21821 32759 21879 32765
rect 21821 32725 21833 32759
rect 21867 32756 21879 32759
rect 21910 32756 21916 32768
rect 21867 32728 21916 32756
rect 21867 32725 21879 32728
rect 21821 32719 21879 32725
rect 21910 32716 21916 32728
rect 21968 32716 21974 32768
rect 23845 32759 23903 32765
rect 23845 32725 23857 32759
rect 23891 32756 23903 32759
rect 24026 32756 24032 32768
rect 23891 32728 24032 32756
rect 23891 32725 23903 32728
rect 23845 32719 23903 32725
rect 24026 32716 24032 32728
rect 24084 32716 24090 32768
rect 32398 32716 32404 32768
rect 32456 32756 32462 32768
rect 32493 32759 32551 32765
rect 32493 32756 32505 32759
rect 32456 32728 32505 32756
rect 32456 32716 32462 32728
rect 32493 32725 32505 32728
rect 32539 32725 32551 32759
rect 32493 32719 32551 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 4890 32512 4896 32564
rect 4948 32552 4954 32564
rect 5169 32555 5227 32561
rect 5169 32552 5181 32555
rect 4948 32524 5181 32552
rect 4948 32512 4954 32524
rect 5169 32521 5181 32524
rect 5215 32552 5227 32555
rect 5350 32552 5356 32564
rect 5215 32524 5356 32552
rect 5215 32521 5227 32524
rect 5169 32515 5227 32521
rect 5350 32512 5356 32524
rect 5408 32512 5414 32564
rect 5813 32555 5871 32561
rect 5813 32521 5825 32555
rect 5859 32552 5871 32555
rect 6454 32552 6460 32564
rect 5859 32524 6460 32552
rect 5859 32521 5871 32524
rect 5813 32515 5871 32521
rect 6454 32512 6460 32524
rect 6512 32552 6518 32564
rect 6730 32552 6736 32564
rect 6512 32524 6736 32552
rect 6512 32512 6518 32524
rect 6730 32512 6736 32524
rect 6788 32512 6794 32564
rect 7650 32512 7656 32564
rect 7708 32552 7714 32564
rect 8757 32555 8815 32561
rect 8757 32552 8769 32555
rect 7708 32524 8769 32552
rect 7708 32512 7714 32524
rect 8757 32521 8769 32524
rect 8803 32521 8815 32555
rect 9122 32552 9128 32564
rect 8757 32515 8815 32521
rect 8864 32524 9128 32552
rect 5994 32444 6000 32496
rect 6052 32484 6058 32496
rect 8864 32484 8892 32524
rect 9122 32512 9128 32524
rect 9180 32552 9186 32564
rect 9180 32524 13041 32552
rect 9180 32512 9186 32524
rect 6052 32456 8892 32484
rect 8941 32487 8999 32493
rect 6052 32444 6058 32456
rect 8941 32453 8953 32487
rect 8987 32484 8999 32487
rect 9030 32484 9036 32496
rect 8987 32456 9036 32484
rect 8987 32453 8999 32456
rect 8941 32447 8999 32453
rect 7190 32425 7196 32428
rect 7184 32416 7196 32425
rect 7151 32388 7196 32416
rect 7184 32379 7196 32388
rect 7190 32376 7196 32379
rect 7248 32376 7254 32428
rect 6822 32308 6828 32360
rect 6880 32348 6886 32360
rect 6917 32351 6975 32357
rect 6917 32348 6929 32351
rect 6880 32320 6929 32348
rect 6880 32308 6886 32320
rect 6917 32317 6929 32320
rect 6963 32317 6975 32351
rect 6917 32311 6975 32317
rect 8297 32283 8355 32289
rect 8297 32249 8309 32283
rect 8343 32280 8355 32283
rect 8956 32280 8984 32447
rect 9030 32444 9036 32456
rect 9088 32444 9094 32496
rect 11882 32444 11888 32496
rect 11940 32484 11946 32496
rect 12897 32487 12955 32493
rect 12897 32484 12909 32487
rect 11940 32456 12909 32484
rect 11940 32444 11946 32456
rect 12897 32453 12909 32456
rect 12943 32453 12955 32487
rect 13013 32484 13041 32524
rect 13078 32512 13084 32564
rect 13136 32552 13142 32564
rect 13725 32555 13783 32561
rect 13725 32552 13737 32555
rect 13136 32524 13737 32552
rect 13136 32512 13142 32524
rect 13725 32521 13737 32524
rect 13771 32521 13783 32555
rect 13725 32515 13783 32521
rect 13832 32524 17632 32552
rect 13832 32484 13860 32524
rect 13013 32456 13860 32484
rect 13909 32487 13967 32493
rect 12897 32447 12955 32453
rect 13909 32453 13921 32487
rect 13955 32484 13967 32487
rect 14642 32484 14648 32496
rect 13955 32456 14648 32484
rect 13955 32453 13967 32456
rect 13909 32447 13967 32453
rect 14642 32444 14648 32456
rect 14700 32444 14706 32496
rect 17034 32484 17040 32496
rect 16995 32456 17040 32484
rect 17034 32444 17040 32456
rect 17092 32444 17098 32496
rect 9125 32419 9183 32425
rect 9125 32385 9137 32419
rect 9171 32416 9183 32419
rect 9674 32416 9680 32428
rect 9171 32388 9680 32416
rect 9171 32385 9183 32388
rect 9125 32379 9183 32385
rect 9674 32376 9680 32388
rect 9732 32376 9738 32428
rect 12526 32376 12532 32428
rect 12584 32416 12590 32428
rect 12713 32419 12771 32425
rect 12713 32416 12725 32419
rect 12584 32388 12725 32416
rect 12584 32376 12590 32388
rect 12713 32385 12725 32388
rect 12759 32416 12771 32419
rect 13262 32416 13268 32428
rect 12759 32388 13268 32416
rect 12759 32385 12771 32388
rect 12713 32379 12771 32385
rect 13262 32376 13268 32388
rect 13320 32376 13326 32428
rect 14090 32416 14096 32428
rect 14003 32388 14096 32416
rect 14090 32376 14096 32388
rect 14148 32376 14154 32428
rect 16850 32416 16856 32428
rect 16811 32388 16856 32416
rect 16850 32376 16856 32388
rect 16908 32376 16914 32428
rect 10505 32351 10563 32357
rect 10505 32317 10517 32351
rect 10551 32317 10563 32351
rect 10505 32311 10563 32317
rect 10781 32351 10839 32357
rect 10781 32317 10793 32351
rect 10827 32348 10839 32351
rect 13446 32348 13452 32360
rect 10827 32320 13452 32348
rect 10827 32317 10839 32320
rect 10781 32311 10839 32317
rect 8343 32252 8984 32280
rect 8343 32249 8355 32252
rect 8297 32243 8355 32249
rect 7558 32172 7564 32224
rect 7616 32212 7622 32224
rect 10520 32212 10548 32311
rect 13446 32308 13452 32320
rect 13504 32308 13510 32360
rect 12066 32240 12072 32292
rect 12124 32280 12130 32292
rect 14108 32280 14136 32376
rect 17126 32308 17132 32360
rect 17184 32348 17190 32360
rect 17497 32351 17555 32357
rect 17497 32348 17509 32351
rect 17184 32320 17509 32348
rect 17184 32308 17190 32320
rect 17497 32317 17509 32320
rect 17543 32317 17555 32351
rect 17604 32348 17632 32524
rect 18138 32512 18144 32564
rect 18196 32552 18202 32564
rect 18877 32555 18935 32561
rect 18877 32552 18889 32555
rect 18196 32524 18889 32552
rect 18196 32512 18202 32524
rect 18877 32521 18889 32524
rect 18923 32521 18935 32555
rect 21174 32552 21180 32564
rect 21135 32524 21180 32552
rect 18877 32515 18935 32521
rect 21174 32512 21180 32524
rect 21232 32552 21238 32564
rect 21634 32552 21640 32564
rect 21232 32524 21640 32552
rect 21232 32512 21238 32524
rect 21634 32512 21640 32524
rect 21692 32512 21698 32564
rect 22094 32512 22100 32564
rect 22152 32552 22158 32564
rect 24489 32555 24547 32561
rect 22152 32524 22197 32552
rect 22152 32512 22158 32524
rect 24489 32521 24501 32555
rect 24535 32552 24547 32555
rect 24854 32552 24860 32564
rect 24535 32524 24860 32552
rect 24535 32521 24547 32524
rect 24489 32515 24547 32521
rect 24854 32512 24860 32524
rect 24912 32512 24918 32564
rect 24949 32555 25007 32561
rect 24949 32521 24961 32555
rect 24995 32521 25007 32555
rect 24949 32515 25007 32521
rect 18506 32444 18512 32496
rect 18564 32484 18570 32496
rect 18969 32487 19027 32493
rect 18969 32484 18981 32487
rect 18564 32456 18981 32484
rect 18564 32444 18570 32456
rect 18969 32453 18981 32456
rect 19015 32484 19027 32487
rect 19613 32487 19671 32493
rect 19613 32484 19625 32487
rect 19015 32456 19625 32484
rect 19015 32453 19027 32456
rect 18969 32447 19027 32453
rect 19613 32453 19625 32456
rect 19659 32484 19671 32487
rect 22741 32487 22799 32493
rect 22741 32484 22753 32487
rect 19659 32456 22753 32484
rect 19659 32453 19671 32456
rect 19613 32447 19671 32453
rect 22741 32453 22753 32456
rect 22787 32484 22799 32487
rect 22787 32456 23428 32484
rect 22787 32453 22799 32456
rect 22741 32447 22799 32453
rect 17773 32419 17831 32425
rect 17773 32385 17785 32419
rect 17819 32416 17831 32419
rect 18690 32416 18696 32428
rect 17819 32388 18696 32416
rect 17819 32385 17831 32388
rect 17773 32379 17831 32385
rect 18690 32376 18696 32388
rect 18748 32376 18754 32428
rect 21910 32416 21916 32428
rect 21871 32388 21916 32416
rect 21910 32376 21916 32388
rect 21968 32416 21974 32428
rect 22830 32416 22836 32428
rect 21968 32388 22836 32416
rect 21968 32376 21974 32388
rect 22830 32376 22836 32388
rect 22888 32376 22894 32428
rect 23400 32425 23428 32456
rect 23750 32444 23756 32496
rect 23808 32484 23814 32496
rect 24305 32487 24363 32493
rect 24305 32484 24317 32487
rect 23808 32456 24317 32484
rect 23808 32444 23814 32456
rect 24305 32453 24317 32456
rect 24351 32484 24363 32487
rect 24964 32484 24992 32515
rect 25406 32512 25412 32564
rect 25464 32552 25470 32564
rect 28721 32555 28779 32561
rect 28721 32552 28733 32555
rect 25464 32524 28733 32552
rect 25464 32512 25470 32524
rect 28721 32521 28733 32524
rect 28767 32521 28779 32555
rect 28721 32515 28779 32521
rect 28810 32512 28816 32564
rect 28868 32552 28874 32564
rect 29730 32552 29736 32564
rect 28868 32524 29316 32552
rect 29691 32524 29736 32552
rect 28868 32512 28874 32524
rect 24351 32456 24992 32484
rect 24351 32453 24363 32456
rect 24305 32447 24363 32453
rect 25314 32444 25320 32496
rect 25372 32484 25378 32496
rect 26062 32487 26120 32493
rect 26062 32484 26074 32487
rect 25372 32456 26074 32484
rect 25372 32444 25378 32456
rect 26062 32453 26074 32456
rect 26108 32453 26120 32487
rect 26062 32447 26120 32453
rect 27985 32487 28043 32493
rect 27985 32453 27997 32487
rect 28031 32484 28043 32487
rect 28442 32484 28448 32496
rect 28031 32456 28448 32484
rect 28031 32453 28043 32456
rect 27985 32447 28043 32453
rect 28442 32444 28448 32456
rect 28500 32444 28506 32496
rect 28534 32444 28540 32496
rect 28592 32484 28598 32496
rect 28997 32487 29055 32493
rect 28997 32484 29009 32487
rect 28592 32456 29009 32484
rect 28592 32444 28598 32456
rect 28997 32453 29009 32456
rect 29043 32453 29055 32487
rect 28997 32447 29055 32453
rect 23385 32419 23443 32425
rect 23385 32385 23397 32419
rect 23431 32416 23443 32419
rect 24026 32416 24032 32428
rect 23431 32388 24032 32416
rect 23431 32385 23443 32388
rect 23385 32379 23443 32385
rect 24026 32376 24032 32388
rect 24084 32376 24090 32428
rect 24121 32419 24179 32425
rect 24121 32385 24133 32419
rect 24167 32416 24179 32419
rect 24210 32416 24216 32428
rect 24167 32388 24216 32416
rect 24167 32385 24179 32388
rect 24121 32379 24179 32385
rect 24210 32376 24216 32388
rect 24268 32376 24274 32428
rect 27893 32419 27951 32425
rect 27893 32385 27905 32419
rect 27939 32416 27951 32419
rect 28077 32419 28135 32425
rect 27939 32388 28028 32416
rect 27939 32385 27951 32388
rect 27893 32379 27951 32385
rect 20806 32348 20812 32360
rect 17604 32320 20812 32348
rect 17497 32311 17555 32317
rect 20806 32308 20812 32320
rect 20864 32308 20870 32360
rect 26329 32351 26387 32357
rect 26329 32317 26341 32351
rect 26375 32348 26387 32351
rect 27154 32348 27160 32360
rect 26375 32320 27160 32348
rect 26375 32317 26387 32320
rect 26329 32311 26387 32317
rect 27154 32308 27160 32320
rect 27212 32308 27218 32360
rect 12124 32252 14136 32280
rect 12124 32240 12130 32252
rect 21358 32240 21364 32292
rect 21416 32280 21422 32292
rect 23569 32283 23627 32289
rect 23569 32280 23581 32283
rect 21416 32252 23581 32280
rect 21416 32240 21422 32252
rect 23569 32249 23581 32252
rect 23615 32280 23627 32283
rect 23842 32280 23848 32292
rect 23615 32252 23848 32280
rect 23615 32249 23627 32252
rect 23569 32243 23627 32249
rect 23842 32240 23848 32252
rect 23900 32240 23906 32292
rect 7616 32184 10548 32212
rect 13081 32215 13139 32221
rect 7616 32172 7622 32184
rect 13081 32181 13093 32215
rect 13127 32212 13139 32215
rect 13630 32212 13636 32224
rect 13127 32184 13636 32212
rect 13127 32181 13139 32184
rect 13081 32175 13139 32181
rect 13630 32172 13636 32184
rect 13688 32172 13694 32224
rect 25038 32172 25044 32224
rect 25096 32212 25102 32224
rect 27709 32215 27767 32221
rect 27709 32212 27721 32215
rect 25096 32184 27721 32212
rect 25096 32172 25102 32184
rect 27709 32181 27721 32184
rect 27755 32181 27767 32215
rect 28000 32212 28028 32388
rect 28077 32385 28089 32419
rect 28123 32385 28135 32419
rect 28077 32379 28135 32385
rect 28092 32280 28120 32379
rect 28166 32376 28172 32428
rect 28224 32416 28230 32428
rect 29288 32425 29316 32524
rect 29730 32512 29736 32524
rect 29788 32512 29794 32564
rect 30558 32484 30564 32496
rect 30519 32456 30564 32484
rect 30558 32444 30564 32456
rect 30616 32484 30622 32496
rect 30742 32484 30748 32496
rect 30616 32456 30748 32484
rect 30616 32444 30622 32456
rect 30742 32444 30748 32456
rect 30800 32444 30806 32496
rect 33042 32444 33048 32496
rect 33100 32484 33106 32496
rect 33100 32456 33916 32484
rect 33100 32444 33106 32456
rect 28261 32419 28319 32425
rect 28261 32416 28273 32419
rect 28224 32388 28273 32416
rect 28224 32376 28230 32388
rect 28261 32385 28273 32388
rect 28307 32385 28319 32419
rect 28261 32379 28319 32385
rect 28905 32419 28963 32425
rect 28905 32385 28917 32419
rect 28951 32385 28963 32419
rect 28905 32379 28963 32385
rect 29089 32419 29147 32425
rect 29089 32385 29101 32419
rect 29135 32385 29147 32419
rect 29089 32379 29147 32385
rect 29273 32419 29331 32425
rect 29273 32385 29285 32419
rect 29319 32385 29331 32419
rect 29273 32379 29331 32385
rect 28920 32348 28948 32379
rect 28994 32348 29000 32360
rect 28920 32320 29000 32348
rect 28994 32308 29000 32320
rect 29052 32308 29058 32360
rect 29104 32280 29132 32379
rect 32858 32376 32864 32428
rect 32916 32416 32922 32428
rect 33698 32419 33756 32425
rect 33698 32416 33710 32419
rect 32916 32388 33710 32416
rect 32916 32376 32922 32388
rect 33698 32385 33710 32388
rect 33744 32385 33756 32419
rect 33698 32379 33756 32385
rect 33888 32348 33916 32456
rect 33965 32419 34023 32425
rect 33965 32385 33977 32419
rect 34011 32416 34023 32419
rect 36170 32416 36176 32428
rect 34011 32388 36176 32416
rect 34011 32385 34023 32388
rect 33965 32379 34023 32385
rect 36170 32376 36176 32388
rect 36228 32416 36234 32428
rect 37458 32416 37464 32428
rect 36228 32388 37464 32416
rect 36228 32376 36234 32388
rect 37458 32376 37464 32388
rect 37516 32376 37522 32428
rect 37550 32376 37556 32428
rect 37608 32416 37614 32428
rect 37717 32419 37775 32425
rect 37717 32416 37729 32419
rect 37608 32388 37729 32416
rect 37608 32376 37614 32388
rect 37717 32385 37729 32388
rect 37763 32385 37775 32419
rect 37717 32379 37775 32385
rect 33888 32320 35940 32348
rect 30558 32280 30564 32292
rect 28092 32252 30564 32280
rect 30558 32240 30564 32252
rect 30616 32240 30622 32292
rect 35912 32224 35940 32320
rect 28994 32212 29000 32224
rect 28000 32184 29000 32212
rect 27709 32175 27767 32181
rect 28994 32172 29000 32184
rect 29052 32212 29058 32224
rect 30098 32212 30104 32224
rect 29052 32184 30104 32212
rect 29052 32172 29058 32184
rect 30098 32172 30104 32184
rect 30156 32172 30162 32224
rect 30466 32212 30472 32224
rect 30427 32184 30472 32212
rect 30466 32172 30472 32184
rect 30524 32212 30530 32224
rect 30834 32212 30840 32224
rect 30524 32184 30840 32212
rect 30524 32172 30530 32184
rect 30834 32172 30840 32184
rect 30892 32172 30898 32224
rect 32585 32215 32643 32221
rect 32585 32181 32597 32215
rect 32631 32212 32643 32215
rect 33226 32212 33232 32224
rect 32631 32184 33232 32212
rect 32631 32181 32643 32184
rect 32585 32175 32643 32181
rect 33226 32172 33232 32184
rect 33284 32212 33290 32224
rect 33778 32212 33784 32224
rect 33284 32184 33784 32212
rect 33284 32172 33290 32184
rect 33778 32172 33784 32184
rect 33836 32172 33842 32224
rect 35894 32212 35900 32224
rect 35855 32184 35900 32212
rect 35894 32172 35900 32184
rect 35952 32172 35958 32224
rect 38654 32172 38660 32224
rect 38712 32212 38718 32224
rect 38841 32215 38899 32221
rect 38841 32212 38853 32215
rect 38712 32184 38853 32212
rect 38712 32172 38718 32184
rect 38841 32181 38853 32184
rect 38887 32181 38899 32215
rect 58158 32212 58164 32224
rect 58119 32184 58164 32212
rect 38841 32175 38899 32181
rect 58158 32172 58164 32184
rect 58216 32172 58222 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 6730 32008 6736 32020
rect 5000 31980 6736 32008
rect 1857 31807 1915 31813
rect 1857 31773 1869 31807
rect 1903 31804 1915 31807
rect 2406 31804 2412 31816
rect 1903 31776 2412 31804
rect 1903 31773 1915 31776
rect 1857 31767 1915 31773
rect 2406 31764 2412 31776
rect 2464 31764 2470 31816
rect 5000 31813 5028 31980
rect 6730 31968 6736 31980
rect 6788 31968 6794 32020
rect 13446 31968 13452 32020
rect 13504 32008 13510 32020
rect 16022 32008 16028 32020
rect 13504 31980 16028 32008
rect 13504 31968 13510 31980
rect 16022 31968 16028 31980
rect 16080 32008 16086 32020
rect 17126 32008 17132 32020
rect 16080 31980 17132 32008
rect 16080 31968 16086 31980
rect 17126 31968 17132 31980
rect 17184 31968 17190 32020
rect 22830 31968 22836 32020
rect 22888 32008 22894 32020
rect 22925 32011 22983 32017
rect 22925 32008 22937 32011
rect 22888 31980 22937 32008
rect 22888 31968 22894 31980
rect 22925 31977 22937 31980
rect 22971 31977 22983 32011
rect 23658 32008 23664 32020
rect 23619 31980 23664 32008
rect 22925 31971 22983 31977
rect 5258 31900 5264 31952
rect 5316 31940 5322 31952
rect 5316 31912 6132 31940
rect 5316 31900 5322 31912
rect 5368 31872 5396 31912
rect 5276 31844 5396 31872
rect 6104 31872 6132 31912
rect 6178 31900 6184 31952
rect 6236 31940 6242 31952
rect 6822 31940 6828 31952
rect 6236 31912 6828 31940
rect 6236 31900 6242 31912
rect 6822 31900 6828 31912
rect 6880 31940 6886 31952
rect 11882 31940 11888 31952
rect 6880 31912 9628 31940
rect 11843 31912 11888 31940
rect 6880 31900 6886 31912
rect 7190 31872 7196 31884
rect 6104 31844 6592 31872
rect 4985 31807 5043 31813
rect 4985 31773 4997 31807
rect 5031 31773 5043 31807
rect 5166 31804 5172 31816
rect 5127 31776 5172 31804
rect 4985 31767 5043 31773
rect 5166 31764 5172 31776
rect 5224 31764 5230 31816
rect 5276 31813 5304 31844
rect 5261 31807 5319 31813
rect 5261 31773 5273 31807
rect 5307 31773 5319 31807
rect 5261 31767 5319 31773
rect 5350 31764 5356 31816
rect 5408 31804 5414 31816
rect 5408 31776 5453 31804
rect 5408 31764 5414 31776
rect 5994 31764 6000 31816
rect 6052 31804 6058 31816
rect 6564 31813 6592 31844
rect 6656 31844 7196 31872
rect 6656 31813 6684 31844
rect 7190 31832 7196 31844
rect 7248 31832 7254 31884
rect 7282 31832 7288 31884
rect 7340 31872 7346 31884
rect 9600 31881 9628 31912
rect 11882 31900 11888 31912
rect 11940 31900 11946 31952
rect 22143 31943 22201 31949
rect 22143 31909 22155 31943
rect 22189 31940 22201 31943
rect 22554 31940 22560 31952
rect 22189 31912 22560 31940
rect 22189 31909 22201 31912
rect 22143 31903 22201 31909
rect 22554 31900 22560 31912
rect 22612 31900 22618 31952
rect 8113 31875 8171 31881
rect 8113 31872 8125 31875
rect 7340 31844 8125 31872
rect 7340 31832 7346 31844
rect 8113 31841 8125 31844
rect 8159 31841 8171 31875
rect 8113 31835 8171 31841
rect 9585 31875 9643 31881
rect 9585 31841 9597 31875
rect 9631 31841 9643 31875
rect 16393 31875 16451 31881
rect 16393 31872 16405 31875
rect 9585 31835 9643 31841
rect 13188 31844 16405 31872
rect 6457 31807 6515 31813
rect 6457 31804 6469 31807
rect 6052 31776 6469 31804
rect 6052 31764 6058 31776
rect 6457 31773 6469 31776
rect 6503 31773 6515 31807
rect 6457 31767 6515 31773
rect 6549 31807 6607 31813
rect 6549 31773 6561 31807
rect 6595 31773 6607 31807
rect 6549 31767 6607 31773
rect 6641 31807 6699 31813
rect 6641 31773 6653 31807
rect 6687 31773 6699 31807
rect 6641 31767 6699 31773
rect 6730 31764 6736 31816
rect 6788 31804 6794 31816
rect 6825 31807 6883 31813
rect 6825 31804 6837 31807
rect 6788 31776 6837 31804
rect 6788 31764 6794 31776
rect 6825 31773 6837 31776
rect 6871 31773 6883 31807
rect 6825 31767 6883 31773
rect 8389 31807 8447 31813
rect 8389 31773 8401 31807
rect 8435 31804 8447 31807
rect 8478 31804 8484 31816
rect 8435 31776 8484 31804
rect 8435 31773 8447 31776
rect 8389 31767 8447 31773
rect 8478 31764 8484 31776
rect 8536 31764 8542 31816
rect 9858 31813 9864 31816
rect 9852 31804 9864 31813
rect 9819 31776 9864 31804
rect 9852 31767 9864 31776
rect 9858 31764 9864 31767
rect 9916 31764 9922 31816
rect 11514 31764 11520 31816
rect 11572 31804 11578 31816
rect 13188 31804 13216 31844
rect 16393 31841 16405 31844
rect 16439 31872 16451 31875
rect 22373 31875 22431 31881
rect 22373 31872 22385 31875
rect 16439 31844 16988 31872
rect 16439 31841 16451 31844
rect 16393 31835 16451 31841
rect 11572 31776 13216 31804
rect 13265 31807 13323 31813
rect 11572 31764 11578 31776
rect 12360 31748 12388 31776
rect 13265 31773 13277 31807
rect 13311 31804 13323 31807
rect 14734 31804 14740 31816
rect 13311 31776 14740 31804
rect 13311 31773 13323 31776
rect 13265 31767 13323 31773
rect 14734 31764 14740 31776
rect 14792 31764 14798 31816
rect 16960 31813 16988 31844
rect 22066 31844 22385 31872
rect 16945 31807 17003 31813
rect 16945 31773 16957 31807
rect 16991 31773 17003 31807
rect 16945 31767 17003 31773
rect 18782 31764 18788 31816
rect 18840 31804 18846 31816
rect 20993 31807 21051 31813
rect 20993 31804 21005 31807
rect 18840 31776 21005 31804
rect 18840 31764 18846 31776
rect 20993 31773 21005 31776
rect 21039 31804 21051 31807
rect 22066 31804 22094 31844
rect 22373 31841 22385 31844
rect 22419 31841 22431 31875
rect 22373 31835 22431 31841
rect 22646 31832 22652 31884
rect 22704 31872 22710 31884
rect 22830 31872 22836 31884
rect 22704 31844 22836 31872
rect 22704 31832 22710 31844
rect 22830 31832 22836 31844
rect 22888 31832 22894 31884
rect 21039 31776 22094 31804
rect 22940 31804 22968 31971
rect 23658 31968 23664 31980
rect 23716 31968 23722 32020
rect 23842 31968 23848 32020
rect 23900 32008 23906 32020
rect 24118 32008 24124 32020
rect 23900 31980 24124 32008
rect 23900 31968 23906 31980
rect 24118 31968 24124 31980
rect 24176 31968 24182 32020
rect 29914 31968 29920 32020
rect 29972 32008 29978 32020
rect 30009 32011 30067 32017
rect 30009 32008 30021 32011
rect 29972 31980 30021 32008
rect 29972 31968 29978 31980
rect 30009 31977 30021 31980
rect 30055 31977 30067 32011
rect 32858 32008 32864 32020
rect 32819 31980 32864 32008
rect 30009 31971 30067 31977
rect 32858 31968 32864 31980
rect 32916 31968 32922 32020
rect 36633 32011 36691 32017
rect 36633 31977 36645 32011
rect 36679 32008 36691 32011
rect 37550 32008 37556 32020
rect 36679 31980 37556 32008
rect 36679 31977 36691 31980
rect 36633 31971 36691 31977
rect 37550 31968 37556 31980
rect 37608 31968 37614 32020
rect 30745 31943 30803 31949
rect 30745 31909 30757 31943
rect 30791 31940 30803 31943
rect 31662 31940 31668 31952
rect 30791 31912 31668 31940
rect 30791 31909 30803 31912
rect 30745 31903 30803 31909
rect 31662 31900 31668 31912
rect 31720 31900 31726 31952
rect 33318 31940 33324 31952
rect 32232 31912 33324 31940
rect 27154 31872 27160 31884
rect 27115 31844 27160 31872
rect 27154 31832 27160 31844
rect 27212 31832 27218 31884
rect 30282 31872 30288 31884
rect 29748 31844 30288 31872
rect 29748 31816 29776 31844
rect 30282 31832 30288 31844
rect 30340 31832 30346 31884
rect 23477 31807 23535 31813
rect 23477 31804 23489 31807
rect 22940 31776 23489 31804
rect 21039 31773 21051 31776
rect 20993 31767 21051 31773
rect 2130 31745 2136 31748
rect 2124 31699 2136 31745
rect 2188 31736 2194 31748
rect 2188 31708 2224 31736
rect 2130 31696 2136 31699
rect 2188 31696 2194 31708
rect 12342 31696 12348 31748
rect 12400 31696 12406 31748
rect 12986 31736 12992 31748
rect 13044 31745 13050 31748
rect 12956 31708 12992 31736
rect 12986 31696 12992 31708
rect 13044 31699 13056 31745
rect 23400 31736 23428 31776
rect 23477 31773 23489 31776
rect 23523 31773 23535 31807
rect 23477 31767 23535 31773
rect 28813 31807 28871 31813
rect 28813 31773 28825 31807
rect 28859 31804 28871 31807
rect 29730 31804 29736 31816
rect 28859 31776 29736 31804
rect 28859 31773 28871 31776
rect 28813 31767 28871 31773
rect 29730 31764 29736 31776
rect 29788 31764 29794 31816
rect 30193 31807 30251 31813
rect 30193 31773 30205 31807
rect 30239 31804 30251 31807
rect 30742 31804 30748 31816
rect 30239 31776 30748 31804
rect 30239 31773 30251 31776
rect 30193 31767 30251 31773
rect 30742 31764 30748 31776
rect 30800 31764 30806 31816
rect 30926 31804 30932 31816
rect 30887 31776 30932 31804
rect 30926 31764 30932 31776
rect 30984 31764 30990 31816
rect 31018 31764 31024 31816
rect 31076 31804 31082 31816
rect 31294 31804 31300 31816
rect 31076 31776 31121 31804
rect 31255 31776 31300 31804
rect 31076 31764 31082 31776
rect 31294 31764 31300 31776
rect 31352 31764 31358 31816
rect 32232 31813 32260 31912
rect 33318 31900 33324 31912
rect 33376 31900 33382 31952
rect 35894 31900 35900 31952
rect 35952 31940 35958 31952
rect 35952 31912 36492 31940
rect 35952 31900 35958 31912
rect 32950 31872 32956 31884
rect 32517 31844 32956 31872
rect 32217 31807 32275 31813
rect 32217 31773 32229 31807
rect 32263 31773 32275 31807
rect 32398 31804 32404 31816
rect 32359 31776 32404 31804
rect 32217 31767 32275 31773
rect 32398 31764 32404 31776
rect 32456 31764 32462 31816
rect 32517 31813 32545 31844
rect 32950 31832 32956 31844
rect 33008 31832 33014 31884
rect 35529 31875 35587 31881
rect 35529 31841 35541 31875
rect 35575 31872 35587 31875
rect 36078 31872 36084 31884
rect 35575 31844 36084 31872
rect 35575 31841 35587 31844
rect 35529 31835 35587 31841
rect 36078 31832 36084 31844
rect 36136 31832 36142 31884
rect 32512 31807 32570 31813
rect 32512 31773 32524 31807
rect 32558 31773 32570 31807
rect 32512 31767 32570 31773
rect 32605 31807 32663 31813
rect 32605 31773 32617 31807
rect 32651 31804 32663 31807
rect 32858 31804 32864 31816
rect 32651 31776 32864 31804
rect 32651 31773 32663 31776
rect 32605 31767 32663 31773
rect 32858 31764 32864 31776
rect 32916 31764 32922 31816
rect 35345 31807 35403 31813
rect 35345 31773 35357 31807
rect 35391 31804 35403 31807
rect 35434 31804 35440 31816
rect 35391 31776 35440 31804
rect 35391 31773 35403 31776
rect 35345 31767 35403 31773
rect 35434 31764 35440 31776
rect 35492 31764 35498 31816
rect 35986 31804 35992 31816
rect 35947 31776 35992 31804
rect 35986 31764 35992 31776
rect 36044 31764 36050 31816
rect 36170 31804 36176 31816
rect 36131 31776 36176 31804
rect 36170 31764 36176 31776
rect 36228 31764 36234 31816
rect 36265 31807 36323 31813
rect 36265 31773 36277 31807
rect 36311 31773 36323 31807
rect 36265 31767 36323 31773
rect 36377 31807 36435 31813
rect 36377 31773 36389 31807
rect 36423 31804 36435 31807
rect 36464 31804 36492 31912
rect 36423 31776 36492 31804
rect 36423 31773 36435 31776
rect 36377 31767 36435 31773
rect 28074 31736 28080 31748
rect 23400 31708 28080 31736
rect 13044 31696 13050 31699
rect 28074 31696 28080 31708
rect 28132 31696 28138 31748
rect 31113 31739 31171 31745
rect 31113 31705 31125 31739
rect 31159 31736 31171 31739
rect 31202 31736 31208 31748
rect 31159 31708 31208 31736
rect 31159 31705 31171 31708
rect 31113 31699 31171 31705
rect 31202 31696 31208 31708
rect 31260 31696 31266 31748
rect 35158 31736 35164 31748
rect 35119 31708 35164 31736
rect 35158 31696 35164 31708
rect 35216 31696 35222 31748
rect 3237 31671 3295 31677
rect 3237 31637 3249 31671
rect 3283 31668 3295 31671
rect 3418 31668 3424 31680
rect 3283 31640 3424 31668
rect 3283 31637 3295 31640
rect 3237 31631 3295 31637
rect 3418 31628 3424 31640
rect 3476 31628 3482 31680
rect 5626 31668 5632 31680
rect 5587 31640 5632 31668
rect 5626 31628 5632 31640
rect 5684 31628 5690 31680
rect 6178 31668 6184 31680
rect 6139 31640 6184 31668
rect 6178 31628 6184 31640
rect 6236 31628 6242 31680
rect 10962 31668 10968 31680
rect 10923 31640 10968 31668
rect 10962 31628 10968 31640
rect 11020 31628 11026 31680
rect 13354 31628 13360 31680
rect 13412 31668 13418 31680
rect 14185 31671 14243 31677
rect 14185 31668 14197 31671
rect 13412 31640 14197 31668
rect 13412 31628 13418 31640
rect 14185 31637 14197 31640
rect 14231 31668 14243 31671
rect 15010 31668 15016 31680
rect 14231 31640 15016 31668
rect 14231 31637 14243 31640
rect 14185 31631 14243 31637
rect 15010 31628 15016 31640
rect 15068 31628 15074 31680
rect 17954 31628 17960 31680
rect 18012 31668 18018 31680
rect 18233 31671 18291 31677
rect 18233 31668 18245 31671
rect 18012 31640 18245 31668
rect 18012 31628 18018 31640
rect 18233 31637 18245 31640
rect 18279 31637 18291 31671
rect 18233 31631 18291 31637
rect 24670 31628 24676 31680
rect 24728 31668 24734 31680
rect 34054 31668 34060 31680
rect 24728 31640 34060 31668
rect 24728 31628 24734 31640
rect 34054 31628 34060 31640
rect 34112 31628 34118 31680
rect 36280 31668 36308 31767
rect 36354 31668 36360 31680
rect 36280 31640 36360 31668
rect 36354 31628 36360 31640
rect 36412 31628 36418 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 2130 31464 2136 31476
rect 2091 31436 2136 31464
rect 2130 31424 2136 31436
rect 2188 31424 2194 31476
rect 5166 31424 5172 31476
rect 5224 31464 5230 31476
rect 5445 31467 5503 31473
rect 5445 31464 5457 31467
rect 5224 31436 5457 31464
rect 5224 31424 5230 31436
rect 5445 31433 5457 31436
rect 5491 31433 5503 31467
rect 6730 31464 6736 31476
rect 5445 31427 5503 31433
rect 5644 31436 6736 31464
rect 2682 31396 2688 31408
rect 2516 31368 2688 31396
rect 2516 31337 2544 31368
rect 2682 31356 2688 31368
rect 2740 31356 2746 31408
rect 5644 31405 5672 31436
rect 6730 31424 6736 31436
rect 6788 31424 6794 31476
rect 12986 31424 12992 31476
rect 13044 31464 13050 31476
rect 13081 31467 13139 31473
rect 13081 31464 13093 31467
rect 13044 31436 13093 31464
rect 13044 31424 13050 31436
rect 13081 31433 13093 31436
rect 13127 31433 13139 31467
rect 17681 31467 17739 31473
rect 17681 31464 17693 31467
rect 13081 31427 13139 31433
rect 13280 31436 17693 31464
rect 5629 31399 5687 31405
rect 5629 31365 5641 31399
rect 5675 31365 5687 31399
rect 5629 31359 5687 31365
rect 6178 31356 6184 31408
rect 6236 31396 6242 31408
rect 6610 31399 6668 31405
rect 6610 31396 6622 31399
rect 6236 31368 6622 31396
rect 6236 31356 6242 31368
rect 6610 31365 6622 31368
rect 6656 31365 6668 31399
rect 6610 31359 6668 31365
rect 11882 31356 11888 31408
rect 11940 31396 11946 31408
rect 12345 31399 12403 31405
rect 12345 31396 12357 31399
rect 11940 31368 12357 31396
rect 11940 31356 11946 31368
rect 12345 31365 12357 31368
rect 12391 31365 12403 31399
rect 12345 31359 12403 31365
rect 12894 31356 12900 31408
rect 12952 31396 12958 31408
rect 13280 31396 13308 31436
rect 17681 31433 17693 31436
rect 17727 31464 17739 31467
rect 18322 31464 18328 31476
rect 17727 31436 18328 31464
rect 17727 31433 17739 31436
rect 17681 31427 17739 31433
rect 18322 31424 18328 31436
rect 18380 31424 18386 31476
rect 24210 31464 24216 31476
rect 24171 31436 24216 31464
rect 24210 31424 24216 31436
rect 24268 31424 24274 31476
rect 32766 31464 32772 31476
rect 28184 31436 32772 31464
rect 12952 31368 13308 31396
rect 14921 31399 14979 31405
rect 12952 31356 12958 31368
rect 14921 31365 14933 31399
rect 14967 31396 14979 31399
rect 15838 31396 15844 31408
rect 14967 31368 15844 31396
rect 14967 31365 14979 31368
rect 14921 31359 14979 31365
rect 15838 31356 15844 31368
rect 15896 31356 15902 31408
rect 16022 31396 16028 31408
rect 15983 31368 16028 31396
rect 16022 31356 16028 31368
rect 16080 31356 16086 31408
rect 23014 31396 23020 31408
rect 22975 31368 23020 31396
rect 23014 31356 23020 31368
rect 23072 31356 23078 31408
rect 28184 31405 28212 31436
rect 32766 31424 32772 31436
rect 32824 31424 32830 31476
rect 35437 31467 35495 31473
rect 35437 31433 35449 31467
rect 35483 31464 35495 31467
rect 36170 31464 36176 31476
rect 35483 31436 36176 31464
rect 35483 31433 35495 31436
rect 35437 31427 35495 31433
rect 36170 31424 36176 31436
rect 36228 31424 36234 31476
rect 28169 31399 28227 31405
rect 28169 31365 28181 31399
rect 28215 31365 28227 31399
rect 29454 31396 29460 31408
rect 28169 31359 28227 31365
rect 28552 31368 29460 31396
rect 2389 31331 2447 31337
rect 2389 31297 2401 31331
rect 2435 31328 2447 31331
rect 2501 31331 2559 31337
rect 2435 31297 2452 31328
rect 2389 31291 2452 31297
rect 2501 31297 2513 31331
rect 2547 31297 2559 31331
rect 2501 31291 2559 31297
rect 2598 31334 2656 31340
rect 2598 31300 2610 31334
rect 2644 31328 2656 31334
rect 2777 31331 2835 31337
rect 2644 31300 2749 31328
rect 2598 31294 2656 31300
rect 2424 31192 2452 31291
rect 2721 31260 2749 31300
rect 2777 31297 2789 31331
rect 2823 31328 2835 31331
rect 2866 31328 2872 31340
rect 2823 31300 2872 31328
rect 2823 31297 2835 31300
rect 2777 31291 2835 31297
rect 2866 31288 2872 31300
rect 2924 31288 2930 31340
rect 3418 31328 3424 31340
rect 3379 31300 3424 31328
rect 3418 31288 3424 31300
rect 3476 31288 3482 31340
rect 3602 31328 3608 31340
rect 3563 31300 3608 31328
rect 3602 31288 3608 31300
rect 3660 31288 3666 31340
rect 5813 31331 5871 31337
rect 5813 31297 5825 31331
rect 5859 31328 5871 31331
rect 7558 31328 7564 31340
rect 5859 31300 7564 31328
rect 5859 31297 5871 31300
rect 5813 31291 5871 31297
rect 7558 31288 7564 31300
rect 7616 31288 7622 31340
rect 8202 31288 8208 31340
rect 8260 31328 8266 31340
rect 10413 31331 10471 31337
rect 10413 31328 10425 31331
rect 8260 31300 10425 31328
rect 8260 31288 8266 31300
rect 10413 31297 10425 31300
rect 10459 31297 10471 31331
rect 10413 31291 10471 31297
rect 10597 31331 10655 31337
rect 10597 31297 10609 31331
rect 10643 31328 10655 31331
rect 10962 31328 10968 31340
rect 10643 31300 10968 31328
rect 10643 31297 10655 31300
rect 10597 31291 10655 31297
rect 10962 31288 10968 31300
rect 11020 31328 11026 31340
rect 12069 31331 12127 31337
rect 12069 31328 12081 31331
rect 11020 31300 12081 31328
rect 11020 31288 11026 31300
rect 12069 31297 12081 31300
rect 12115 31297 12127 31331
rect 12069 31291 12127 31297
rect 12253 31331 12311 31337
rect 12253 31297 12265 31331
rect 12299 31297 12311 31331
rect 12253 31291 12311 31297
rect 12437 31331 12495 31337
rect 12437 31297 12449 31331
rect 12483 31328 12495 31331
rect 12618 31328 12624 31340
rect 12483 31300 12624 31328
rect 12483 31297 12495 31300
rect 12437 31291 12495 31297
rect 3237 31263 3295 31269
rect 3237 31260 3249 31263
rect 2721 31232 3249 31260
rect 3237 31229 3249 31232
rect 3283 31229 3295 31263
rect 6362 31260 6368 31272
rect 6323 31232 6368 31260
rect 3237 31223 3295 31229
rect 6362 31220 6368 31232
rect 6420 31220 6426 31272
rect 9674 31260 9680 31272
rect 9635 31232 9680 31260
rect 9674 31220 9680 31232
rect 9732 31220 9738 31272
rect 9953 31263 10011 31269
rect 9953 31229 9965 31263
rect 9999 31260 10011 31263
rect 11974 31260 11980 31272
rect 9999 31232 11980 31260
rect 9999 31229 10011 31232
rect 9953 31223 10011 31229
rect 11974 31220 11980 31232
rect 12032 31220 12038 31272
rect 2774 31192 2780 31204
rect 2424 31164 2780 31192
rect 2774 31152 2780 31164
rect 2832 31152 2838 31204
rect 7282 31084 7288 31136
rect 7340 31124 7346 31136
rect 7745 31127 7803 31133
rect 7745 31124 7757 31127
rect 7340 31096 7757 31124
rect 7340 31084 7346 31096
rect 7745 31093 7757 31096
rect 7791 31093 7803 31127
rect 7745 31087 7803 31093
rect 8297 31127 8355 31133
rect 8297 31093 8309 31127
rect 8343 31124 8355 31127
rect 8386 31124 8392 31136
rect 8343 31096 8392 31124
rect 8343 31093 8355 31096
rect 8297 31087 8355 31093
rect 8386 31084 8392 31096
rect 8444 31124 8450 31136
rect 9122 31124 9128 31136
rect 8444 31096 9128 31124
rect 8444 31084 8450 31096
rect 9122 31084 9128 31096
rect 9180 31084 9186 31136
rect 10318 31084 10324 31136
rect 10376 31124 10382 31136
rect 10781 31127 10839 31133
rect 10781 31124 10793 31127
rect 10376 31096 10793 31124
rect 10376 31084 10382 31096
rect 10781 31093 10793 31096
rect 10827 31093 10839 31127
rect 12268 31124 12296 31291
rect 12618 31288 12624 31300
rect 12676 31288 12682 31340
rect 13354 31328 13360 31340
rect 13315 31300 13360 31328
rect 13354 31288 13360 31300
rect 13412 31288 13418 31340
rect 13449 31331 13507 31337
rect 13449 31297 13461 31331
rect 13495 31297 13507 31331
rect 13449 31291 13507 31297
rect 13541 31331 13599 31337
rect 13541 31297 13553 31331
rect 13587 31328 13599 31331
rect 13630 31328 13636 31340
rect 13587 31300 13636 31328
rect 13587 31297 13599 31300
rect 13541 31291 13599 31297
rect 12986 31220 12992 31272
rect 13044 31260 13050 31272
rect 13464 31260 13492 31291
rect 13630 31288 13636 31300
rect 13688 31288 13694 31340
rect 13722 31288 13728 31340
rect 13780 31328 13786 31340
rect 14553 31331 14611 31337
rect 14553 31328 14565 31331
rect 13780 31300 13825 31328
rect 13924 31300 14565 31328
rect 13780 31288 13786 31300
rect 13044 31232 13492 31260
rect 13044 31220 13050 31232
rect 12434 31124 12440 31136
rect 12268 31096 12440 31124
rect 10781 31087 10839 31093
rect 12434 31084 12440 31096
rect 12492 31084 12498 31136
rect 12621 31127 12679 31133
rect 12621 31093 12633 31127
rect 12667 31124 12679 31127
rect 13924 31124 13952 31300
rect 14553 31297 14565 31300
rect 14599 31297 14611 31331
rect 14553 31291 14611 31297
rect 14642 31288 14648 31340
rect 14700 31328 14706 31340
rect 14700 31300 14745 31328
rect 14700 31288 14706 31300
rect 14826 31288 14832 31340
rect 14884 31328 14890 31340
rect 15059 31331 15117 31337
rect 14884 31300 14929 31328
rect 14884 31288 14890 31300
rect 15059 31297 15071 31331
rect 15105 31328 15117 31331
rect 15194 31328 15200 31340
rect 15105 31300 15200 31328
rect 15105 31297 15117 31300
rect 15059 31291 15117 31297
rect 15194 31288 15200 31300
rect 15252 31288 15258 31340
rect 19978 31288 19984 31340
rect 20036 31328 20042 31340
rect 21085 31331 21143 31337
rect 21085 31328 21097 31331
rect 20036 31300 21097 31328
rect 20036 31288 20042 31300
rect 21085 31297 21097 31300
rect 21131 31297 21143 31331
rect 21085 31291 21143 31297
rect 21634 31288 21640 31340
rect 21692 31328 21698 31340
rect 22189 31331 22247 31337
rect 22189 31328 22201 31331
rect 21692 31300 22201 31328
rect 21692 31288 21698 31300
rect 22189 31297 22201 31300
rect 22235 31297 22247 31331
rect 22189 31291 22247 31297
rect 22281 31331 22339 31337
rect 22281 31297 22293 31331
rect 22327 31297 22339 31331
rect 22281 31291 22339 31297
rect 22373 31331 22431 31337
rect 22373 31297 22385 31331
rect 22419 31297 22431 31331
rect 22554 31328 22560 31340
rect 22515 31300 22560 31328
rect 22373 31291 22431 31297
rect 14366 31220 14372 31272
rect 14424 31260 14430 31272
rect 14844 31260 14872 31288
rect 14424 31232 14872 31260
rect 20809 31263 20867 31269
rect 14424 31220 14430 31232
rect 20809 31229 20821 31263
rect 20855 31229 20867 31263
rect 20809 31223 20867 31229
rect 15197 31195 15255 31201
rect 15197 31161 15209 31195
rect 15243 31192 15255 31195
rect 15470 31192 15476 31204
rect 15243 31164 15476 31192
rect 15243 31161 15255 31164
rect 15197 31155 15255 31161
rect 15470 31152 15476 31164
rect 15528 31152 15534 31204
rect 20824 31192 20852 31223
rect 21174 31220 21180 31272
rect 21232 31260 21238 31272
rect 21818 31260 21824 31272
rect 21232 31232 21824 31260
rect 21232 31220 21238 31232
rect 21818 31220 21824 31232
rect 21876 31260 21882 31272
rect 22296 31260 22324 31291
rect 21876 31232 22324 31260
rect 22388 31260 22416 31291
rect 22554 31288 22560 31300
rect 22612 31288 22618 31340
rect 23198 31328 23204 31340
rect 23159 31300 23204 31328
rect 23198 31288 23204 31300
rect 23256 31288 23262 31340
rect 23658 31288 23664 31340
rect 23716 31328 23722 31340
rect 24029 31331 24087 31337
rect 24029 31328 24041 31331
rect 23716 31300 24041 31328
rect 23716 31288 23722 31300
rect 24029 31297 24041 31300
rect 24075 31297 24087 31331
rect 24029 31291 24087 31297
rect 27985 31331 28043 31337
rect 27985 31297 27997 31331
rect 28031 31328 28043 31331
rect 28552 31328 28580 31368
rect 29454 31356 29460 31368
rect 29512 31356 29518 31408
rect 30282 31396 30288 31408
rect 30243 31368 30288 31396
rect 30282 31356 30288 31368
rect 30340 31356 30346 31408
rect 31110 31396 31116 31408
rect 31071 31368 31116 31396
rect 31110 31356 31116 31368
rect 31168 31356 31174 31408
rect 31202 31356 31208 31408
rect 31260 31396 31266 31408
rect 35069 31399 35127 31405
rect 31260 31368 31305 31396
rect 31260 31356 31266 31368
rect 35069 31365 35081 31399
rect 35115 31396 35127 31399
rect 35158 31396 35164 31408
rect 35115 31368 35164 31396
rect 35115 31365 35127 31368
rect 35069 31359 35127 31365
rect 35158 31356 35164 31368
rect 35216 31396 35222 31408
rect 35526 31396 35532 31408
rect 35216 31368 35532 31396
rect 35216 31356 35222 31368
rect 35526 31356 35532 31368
rect 35584 31356 35590 31408
rect 35986 31396 35992 31408
rect 35912 31368 35992 31396
rect 28031 31300 28580 31328
rect 28629 31331 28687 31337
rect 28031 31297 28043 31300
rect 27985 31291 28043 31297
rect 28629 31297 28641 31331
rect 28675 31297 28687 31331
rect 28629 31291 28687 31297
rect 23385 31263 23443 31269
rect 23385 31260 23397 31263
rect 22388 31232 23397 31260
rect 21876 31220 21882 31232
rect 23385 31229 23397 31232
rect 23431 31229 23443 31263
rect 28644 31260 28672 31291
rect 30926 31288 30932 31340
rect 30984 31328 30990 31340
rect 31021 31331 31079 31337
rect 31021 31328 31033 31331
rect 30984 31300 31033 31328
rect 30984 31288 30990 31300
rect 31021 31297 31033 31300
rect 31067 31297 31079 31331
rect 31021 31291 31079 31297
rect 31389 31331 31447 31337
rect 31389 31297 31401 31331
rect 31435 31328 31447 31331
rect 31754 31328 31760 31340
rect 31435 31300 31760 31328
rect 31435 31297 31447 31300
rect 31389 31291 31447 31297
rect 23385 31223 23443 31229
rect 27264 31232 28672 31260
rect 31036 31260 31064 31291
rect 31754 31288 31760 31300
rect 31812 31288 31818 31340
rect 35912 31337 35940 31368
rect 35986 31356 35992 31368
rect 36044 31356 36050 31408
rect 36354 31396 36360 31408
rect 36188 31368 36360 31396
rect 35253 31331 35311 31337
rect 35253 31297 35265 31331
rect 35299 31297 35311 31331
rect 35253 31291 35311 31297
rect 35897 31331 35955 31337
rect 35897 31297 35909 31331
rect 35943 31297 35955 31331
rect 36078 31328 36084 31340
rect 36039 31300 36084 31328
rect 35897 31291 35955 31297
rect 33134 31260 33140 31272
rect 31036 31232 33140 31260
rect 20824 31164 22094 31192
rect 12667 31096 13952 31124
rect 12667 31093 12679 31096
rect 12621 31087 12679 31093
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 15657 31127 15715 31133
rect 15657 31124 15669 31127
rect 15344 31096 15669 31124
rect 15344 31084 15350 31096
rect 15657 31093 15669 31096
rect 15703 31093 15715 31127
rect 19150 31124 19156 31136
rect 19111 31096 19156 31124
rect 15657 31087 15715 31093
rect 19150 31084 19156 31096
rect 19208 31084 19214 31136
rect 19797 31127 19855 31133
rect 19797 31093 19809 31127
rect 19843 31124 19855 31127
rect 19978 31124 19984 31136
rect 19843 31096 19984 31124
rect 19843 31093 19855 31096
rect 19797 31087 19855 31093
rect 19978 31084 19984 31096
rect 20036 31084 20042 31136
rect 21910 31124 21916 31136
rect 21871 31096 21916 31124
rect 21910 31084 21916 31096
rect 21968 31084 21974 31136
rect 22066 31124 22094 31164
rect 22278 31152 22284 31204
rect 22336 31192 22342 31204
rect 27264 31201 27292 31232
rect 33134 31220 33140 31232
rect 33192 31220 33198 31272
rect 33226 31220 33232 31272
rect 33284 31260 33290 31272
rect 35268 31260 35296 31291
rect 36078 31288 36084 31300
rect 36136 31288 36142 31340
rect 36188 31337 36216 31368
rect 36354 31356 36360 31368
rect 36412 31356 36418 31408
rect 36541 31399 36599 31405
rect 36541 31365 36553 31399
rect 36587 31396 36599 31399
rect 38258 31399 38316 31405
rect 38258 31396 38270 31399
rect 36587 31368 38270 31396
rect 36587 31365 36599 31368
rect 36541 31359 36599 31365
rect 38258 31365 38270 31368
rect 38304 31365 38316 31399
rect 38258 31359 38316 31365
rect 36173 31331 36231 31337
rect 36173 31297 36185 31331
rect 36219 31297 36231 31331
rect 36173 31291 36231 31297
rect 36262 31288 36268 31340
rect 36320 31328 36326 31340
rect 37277 31331 37335 31337
rect 37277 31328 37289 31331
rect 36320 31300 37289 31328
rect 36320 31288 36326 31300
rect 37277 31297 37289 31300
rect 37323 31297 37335 31331
rect 37277 31291 37335 31297
rect 37458 31288 37464 31340
rect 37516 31328 37522 31340
rect 37918 31328 37924 31340
rect 37516 31300 37924 31328
rect 37516 31288 37522 31300
rect 37918 31288 37924 31300
rect 37976 31328 37982 31340
rect 38013 31331 38071 31337
rect 38013 31328 38025 31331
rect 37976 31300 38025 31328
rect 37976 31288 37982 31300
rect 38013 31297 38025 31300
rect 38059 31297 38071 31331
rect 38654 31328 38660 31340
rect 38013 31291 38071 31297
rect 38120 31300 38660 31328
rect 38120 31260 38148 31300
rect 38654 31288 38660 31300
rect 38712 31288 38718 31340
rect 33284 31232 38148 31260
rect 33284 31220 33290 31232
rect 27249 31195 27307 31201
rect 27249 31192 27261 31195
rect 22336 31164 27261 31192
rect 22336 31152 22342 31164
rect 27249 31161 27261 31164
rect 27295 31161 27307 31195
rect 27249 31155 27307 31161
rect 23014 31124 23020 31136
rect 22066 31096 23020 31124
rect 23014 31084 23020 31096
rect 23072 31084 23078 31136
rect 24765 31127 24823 31133
rect 24765 31093 24777 31127
rect 24811 31124 24823 31127
rect 24854 31124 24860 31136
rect 24811 31096 24860 31124
rect 24811 31093 24823 31096
rect 24765 31087 24823 31093
rect 24854 31084 24860 31096
rect 24912 31124 24918 31136
rect 25682 31124 25688 31136
rect 24912 31096 25688 31124
rect 24912 31084 24918 31096
rect 25682 31084 25688 31096
rect 25740 31084 25746 31136
rect 27801 31127 27859 31133
rect 27801 31093 27813 31127
rect 27847 31124 27859 31127
rect 28718 31124 28724 31136
rect 27847 31096 28724 31124
rect 27847 31093 27859 31096
rect 27801 31087 27859 31093
rect 28718 31084 28724 31096
rect 28776 31084 28782 31136
rect 30837 31127 30895 31133
rect 30837 31093 30849 31127
rect 30883 31124 30895 31127
rect 31018 31124 31024 31136
rect 30883 31096 31024 31124
rect 30883 31093 30895 31096
rect 30837 31087 30895 31093
rect 31018 31084 31024 31096
rect 31076 31084 31082 31136
rect 32217 31127 32275 31133
rect 32217 31093 32229 31127
rect 32263 31124 32275 31127
rect 32858 31124 32864 31136
rect 32263 31096 32864 31124
rect 32263 31093 32275 31096
rect 32217 31087 32275 31093
rect 32858 31084 32864 31096
rect 32916 31084 32922 31136
rect 35434 31084 35440 31136
rect 35492 31124 35498 31136
rect 39393 31127 39451 31133
rect 39393 31124 39405 31127
rect 35492 31096 39405 31124
rect 35492 31084 35498 31096
rect 39393 31093 39405 31096
rect 39439 31093 39451 31127
rect 39393 31087 39451 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 6362 30920 6368 30932
rect 5368 30892 6368 30920
rect 2406 30744 2412 30796
rect 2464 30784 2470 30796
rect 5368 30793 5396 30892
rect 6362 30880 6368 30892
rect 6420 30880 6426 30932
rect 7190 30920 7196 30932
rect 7151 30892 7196 30920
rect 7190 30880 7196 30892
rect 7248 30880 7254 30932
rect 10873 30923 10931 30929
rect 10873 30889 10885 30923
rect 10919 30920 10931 30923
rect 11514 30920 11520 30932
rect 10919 30892 11520 30920
rect 10919 30889 10931 30892
rect 10873 30883 10931 30889
rect 11514 30880 11520 30892
rect 11572 30880 11578 30932
rect 12713 30923 12771 30929
rect 12713 30920 12725 30923
rect 12406 30892 12725 30920
rect 5353 30787 5411 30793
rect 5353 30784 5365 30787
rect 2464 30756 5365 30784
rect 2464 30744 2470 30756
rect 5353 30753 5365 30756
rect 5399 30753 5411 30787
rect 5353 30747 5411 30753
rect 5626 30725 5632 30728
rect 5620 30716 5632 30725
rect 5587 30688 5632 30716
rect 5620 30679 5632 30688
rect 5626 30676 5632 30679
rect 5684 30676 5690 30728
rect 7558 30716 7564 30728
rect 7519 30688 7564 30716
rect 7558 30676 7564 30688
rect 7616 30676 7622 30728
rect 12161 30719 12219 30725
rect 12161 30685 12173 30719
rect 12207 30716 12219 30719
rect 12406 30716 12434 30892
rect 12713 30889 12725 30892
rect 12759 30920 12771 30923
rect 22925 30923 22983 30929
rect 12759 30892 20300 30920
rect 12759 30889 12771 30892
rect 12713 30883 12771 30889
rect 13722 30812 13728 30864
rect 13780 30852 13786 30864
rect 14093 30855 14151 30861
rect 14093 30852 14105 30855
rect 13780 30824 14105 30852
rect 13780 30812 13786 30824
rect 14093 30821 14105 30824
rect 14139 30821 14151 30855
rect 14093 30815 14151 30821
rect 15838 30812 15844 30864
rect 15896 30852 15902 30864
rect 16117 30855 16175 30861
rect 16117 30852 16129 30855
rect 15896 30824 16129 30852
rect 15896 30812 15902 30824
rect 16117 30821 16129 30824
rect 16163 30821 16175 30855
rect 16117 30815 16175 30821
rect 14734 30784 14740 30796
rect 14695 30756 14740 30784
rect 14734 30744 14740 30756
rect 14792 30744 14798 30796
rect 17954 30744 17960 30796
rect 18012 30784 18018 30796
rect 19242 30784 19248 30796
rect 18012 30756 19248 30784
rect 18012 30744 18018 30756
rect 19242 30744 19248 30756
rect 19300 30744 19306 30796
rect 20272 30784 20300 30892
rect 22925 30889 22937 30923
rect 22971 30920 22983 30923
rect 23198 30920 23204 30932
rect 22971 30892 23204 30920
rect 22971 30889 22983 30892
rect 22925 30883 22983 30889
rect 23198 30880 23204 30892
rect 23256 30880 23262 30932
rect 23661 30923 23719 30929
rect 23661 30889 23673 30923
rect 23707 30920 23719 30923
rect 23842 30920 23848 30932
rect 23707 30892 23848 30920
rect 23707 30889 23719 30892
rect 23661 30883 23719 30889
rect 23842 30880 23848 30892
rect 23900 30880 23906 30932
rect 27801 30923 27859 30929
rect 27801 30889 27813 30923
rect 27847 30920 27859 30923
rect 27890 30920 27896 30932
rect 27847 30892 27896 30920
rect 27847 30889 27859 30892
rect 27801 30883 27859 30889
rect 27890 30880 27896 30892
rect 27948 30880 27954 30932
rect 34054 30880 34060 30932
rect 34112 30920 34118 30932
rect 35253 30923 35311 30929
rect 35253 30920 35265 30923
rect 34112 30892 35265 30920
rect 34112 30880 34118 30892
rect 35253 30889 35265 30892
rect 35299 30889 35311 30923
rect 35253 30883 35311 30889
rect 30558 30812 30564 30864
rect 30616 30852 30622 30864
rect 30616 30824 31616 30852
rect 30616 30812 30622 30824
rect 24673 30787 24731 30793
rect 20272 30756 21680 30784
rect 18322 30716 18328 30728
rect 12207 30688 12434 30716
rect 18283 30688 18328 30716
rect 12207 30685 12219 30688
rect 12161 30679 12219 30685
rect 18322 30676 18328 30688
rect 18380 30676 18386 30728
rect 18417 30719 18475 30725
rect 18417 30685 18429 30719
rect 18463 30685 18475 30719
rect 18417 30679 18475 30685
rect 7282 30608 7288 30660
rect 7340 30648 7346 30660
rect 7377 30651 7435 30657
rect 7377 30648 7389 30651
rect 7340 30620 7389 30648
rect 7340 30608 7346 30620
rect 7377 30617 7389 30620
rect 7423 30617 7435 30651
rect 7377 30611 7435 30617
rect 14734 30608 14740 30660
rect 14792 30648 14798 30660
rect 14982 30651 15040 30657
rect 14982 30648 14994 30651
rect 14792 30620 14994 30648
rect 14792 30608 14798 30620
rect 14982 30617 14994 30620
rect 15028 30617 15040 30651
rect 18432 30648 18460 30679
rect 18506 30676 18512 30728
rect 18564 30716 18570 30728
rect 18693 30719 18751 30725
rect 18564 30688 18609 30716
rect 18564 30676 18570 30688
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 18874 30716 18880 30728
rect 18739 30688 18880 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 18874 30676 18880 30688
rect 18932 30676 18938 30728
rect 21542 30716 21548 30728
rect 21503 30688 21548 30716
rect 21542 30676 21548 30688
rect 21600 30676 21606 30728
rect 21652 30716 21680 30756
rect 24673 30753 24685 30787
rect 24719 30784 24731 30787
rect 24762 30784 24768 30796
rect 24719 30756 24768 30784
rect 24719 30753 24731 30756
rect 24673 30747 24731 30753
rect 24762 30744 24768 30756
rect 24820 30744 24826 30796
rect 30466 30784 30472 30796
rect 28644 30756 30472 30784
rect 22278 30716 22284 30728
rect 21652 30688 22284 30716
rect 22278 30676 22284 30688
rect 22336 30676 22342 30728
rect 23845 30719 23903 30725
rect 23845 30685 23857 30719
rect 23891 30685 23903 30719
rect 24394 30716 24400 30728
rect 24355 30688 24400 30716
rect 23845 30679 23903 30685
rect 14982 30611 15040 30617
rect 17512 30620 18460 30648
rect 19512 30651 19570 30657
rect 2774 30540 2780 30592
rect 2832 30580 2838 30592
rect 2869 30583 2927 30589
rect 2869 30580 2881 30583
rect 2832 30552 2881 30580
rect 2832 30540 2838 30552
rect 2869 30549 2881 30552
rect 2915 30549 2927 30583
rect 6730 30580 6736 30592
rect 6691 30552 6736 30580
rect 2869 30543 2927 30549
rect 6730 30540 6736 30552
rect 6788 30540 6794 30592
rect 16942 30540 16948 30592
rect 17000 30580 17006 30592
rect 17512 30589 17540 30620
rect 19512 30617 19524 30651
rect 19558 30617 19570 30651
rect 19512 30611 19570 30617
rect 21812 30651 21870 30657
rect 21812 30617 21824 30651
rect 21858 30648 21870 30651
rect 21910 30648 21916 30660
rect 21858 30620 21916 30648
rect 21858 30617 21870 30620
rect 21812 30611 21870 30617
rect 17497 30583 17555 30589
rect 17497 30580 17509 30583
rect 17000 30552 17509 30580
rect 17000 30540 17006 30552
rect 17497 30549 17509 30552
rect 17543 30549 17555 30583
rect 18046 30580 18052 30592
rect 18007 30552 18052 30580
rect 17497 30543 17555 30549
rect 18046 30540 18052 30552
rect 18104 30540 18110 30592
rect 19426 30540 19432 30592
rect 19484 30580 19490 30592
rect 19536 30580 19564 30611
rect 21910 30608 21916 30620
rect 21968 30608 21974 30660
rect 23860 30648 23888 30679
rect 24394 30676 24400 30688
rect 24452 30676 24458 30728
rect 27062 30716 27068 30728
rect 27023 30688 27068 30716
rect 27062 30676 27068 30688
rect 27120 30676 27126 30728
rect 27890 30676 27896 30728
rect 27948 30716 27954 30728
rect 28644 30725 28672 30756
rect 30466 30744 30472 30756
rect 30524 30744 30530 30796
rect 30650 30784 30656 30796
rect 30611 30756 30656 30784
rect 30650 30744 30656 30756
rect 30708 30744 30714 30796
rect 28537 30719 28595 30725
rect 28537 30716 28549 30719
rect 27948 30688 28549 30716
rect 27948 30676 27954 30688
rect 28537 30685 28549 30688
rect 28583 30685 28595 30719
rect 28537 30679 28595 30685
rect 28629 30719 28687 30725
rect 28629 30685 28641 30719
rect 28675 30685 28687 30719
rect 28629 30679 28687 30685
rect 28718 30676 28724 30728
rect 28776 30716 28782 30728
rect 28905 30719 28963 30725
rect 28776 30688 28821 30716
rect 28776 30676 28782 30688
rect 28905 30685 28917 30719
rect 28951 30716 28963 30719
rect 28994 30716 29000 30728
rect 28951 30688 29000 30716
rect 28951 30685 28963 30688
rect 28905 30679 28963 30685
rect 28994 30676 29000 30688
rect 29052 30676 29058 30728
rect 30929 30719 30987 30725
rect 30929 30685 30941 30719
rect 30975 30685 30987 30719
rect 31386 30716 31392 30728
rect 31347 30688 31392 30716
rect 30929 30679 30987 30685
rect 24854 30648 24860 30660
rect 23860 30620 24860 30648
rect 24854 30608 24860 30620
rect 24912 30608 24918 30660
rect 26234 30608 26240 30660
rect 26292 30648 26298 30660
rect 26798 30651 26856 30657
rect 26798 30648 26810 30651
rect 26292 30620 26810 30648
rect 26292 30608 26298 30620
rect 26798 30617 26810 30620
rect 26844 30617 26856 30651
rect 30944 30648 30972 30679
rect 31386 30676 31392 30688
rect 31444 30676 31450 30728
rect 31588 30725 31616 30824
rect 31573 30719 31631 30725
rect 31573 30685 31585 30719
rect 31619 30685 31631 30719
rect 33134 30716 33140 30728
rect 33095 30688 33140 30716
rect 31573 30679 31631 30685
rect 33134 30676 33140 30688
rect 33192 30676 33198 30728
rect 33226 30676 33232 30728
rect 33284 30716 33290 30728
rect 33502 30716 33508 30728
rect 33284 30688 33329 30716
rect 33463 30688 33508 30716
rect 33284 30676 33290 30688
rect 33502 30676 33508 30688
rect 33560 30676 33566 30728
rect 31846 30648 31852 30660
rect 30944 30620 31852 30648
rect 26798 30611 26856 30617
rect 31846 30608 31852 30620
rect 31904 30608 31910 30660
rect 32582 30608 32588 30660
rect 32640 30648 32646 30660
rect 33321 30651 33379 30657
rect 33321 30648 33333 30651
rect 32640 30620 33333 30648
rect 32640 30608 32646 30620
rect 33321 30617 33333 30620
rect 33367 30648 33379 30651
rect 33410 30648 33416 30660
rect 33367 30620 33416 30648
rect 33367 30617 33379 30620
rect 33321 30611 33379 30617
rect 33410 30608 33416 30620
rect 33468 30648 33474 30660
rect 33870 30648 33876 30660
rect 33468 30620 33876 30648
rect 33468 30608 33474 30620
rect 33870 30608 33876 30620
rect 33928 30608 33934 30660
rect 35268 30648 35296 30883
rect 35986 30812 35992 30864
rect 36044 30812 36050 30864
rect 36004 30784 36032 30812
rect 36354 30784 36360 30796
rect 35820 30756 36032 30784
rect 36096 30756 36360 30784
rect 35820 30725 35848 30756
rect 35805 30719 35863 30725
rect 35805 30685 35817 30719
rect 35851 30685 35863 30719
rect 35986 30716 35992 30728
rect 35947 30688 35992 30716
rect 35805 30679 35863 30685
rect 35986 30676 35992 30688
rect 36044 30676 36050 30728
rect 36096 30725 36124 30756
rect 36354 30744 36360 30756
rect 36412 30744 36418 30796
rect 37918 30784 37924 30796
rect 37879 30756 37924 30784
rect 37918 30744 37924 30756
rect 37976 30744 37982 30796
rect 36081 30719 36139 30725
rect 36081 30685 36093 30719
rect 36127 30685 36139 30719
rect 36081 30679 36139 30685
rect 36173 30719 36231 30725
rect 36173 30685 36185 30719
rect 36219 30685 36231 30719
rect 58158 30716 58164 30728
rect 58119 30688 58164 30716
rect 36173 30679 36231 30685
rect 36188 30648 36216 30679
rect 58158 30676 58164 30688
rect 58216 30676 58222 30728
rect 35268 30620 36216 30648
rect 36449 30651 36507 30657
rect 36449 30617 36461 30651
rect 36495 30648 36507 30651
rect 38166 30651 38224 30657
rect 38166 30648 38178 30651
rect 36495 30620 38178 30648
rect 36495 30617 36507 30620
rect 36449 30611 36507 30617
rect 38166 30617 38178 30620
rect 38212 30617 38224 30651
rect 38166 30611 38224 30617
rect 19484 30552 19564 30580
rect 19484 30540 19490 30552
rect 20070 30540 20076 30592
rect 20128 30580 20134 30592
rect 20625 30583 20683 30589
rect 20625 30580 20637 30583
rect 20128 30552 20637 30580
rect 20128 30540 20134 30552
rect 20625 30549 20637 30552
rect 20671 30549 20683 30583
rect 20625 30543 20683 30549
rect 22094 30540 22100 30592
rect 22152 30580 22158 30592
rect 23842 30580 23848 30592
rect 22152 30552 23848 30580
rect 22152 30540 22158 30552
rect 23842 30540 23848 30552
rect 23900 30540 23906 30592
rect 25130 30540 25136 30592
rect 25188 30580 25194 30592
rect 25685 30583 25743 30589
rect 25685 30580 25697 30583
rect 25188 30552 25697 30580
rect 25188 30540 25194 30552
rect 25685 30549 25697 30552
rect 25731 30549 25743 30583
rect 25685 30543 25743 30549
rect 28261 30583 28319 30589
rect 28261 30549 28273 30583
rect 28307 30580 28319 30583
rect 28350 30580 28356 30592
rect 28307 30552 28356 30580
rect 28307 30549 28319 30552
rect 28261 30543 28319 30549
rect 28350 30540 28356 30552
rect 28408 30540 28414 30592
rect 31757 30583 31815 30589
rect 31757 30549 31769 30583
rect 31803 30580 31815 30583
rect 32122 30580 32128 30592
rect 31803 30552 32128 30580
rect 31803 30549 31815 30552
rect 31757 30543 31815 30549
rect 32122 30540 32128 30552
rect 32180 30580 32186 30592
rect 32306 30580 32312 30592
rect 32180 30552 32312 30580
rect 32180 30540 32186 30552
rect 32306 30540 32312 30552
rect 32364 30540 32370 30592
rect 32950 30580 32956 30592
rect 32911 30552 32956 30580
rect 32950 30540 32956 30552
rect 33008 30540 33014 30592
rect 37366 30540 37372 30592
rect 37424 30580 37430 30592
rect 39301 30583 39359 30589
rect 39301 30580 39313 30583
rect 37424 30552 39313 30580
rect 37424 30540 37430 30552
rect 39301 30549 39313 30552
rect 39347 30549 39359 30583
rect 39301 30543 39359 30549
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 8478 30336 8484 30388
rect 8536 30376 8542 30388
rect 14734 30376 14740 30388
rect 8536 30348 14601 30376
rect 14695 30348 14740 30376
rect 8536 30336 8542 30348
rect 9858 30308 9864 30320
rect 9819 30280 9864 30308
rect 9858 30268 9864 30280
rect 9916 30268 9922 30320
rect 11517 30311 11575 30317
rect 11517 30308 11529 30311
rect 10152 30280 11529 30308
rect 2406 30240 2412 30252
rect 2367 30212 2412 30240
rect 2406 30200 2412 30212
rect 2464 30200 2470 30252
rect 2498 30200 2504 30252
rect 2556 30240 2562 30252
rect 10152 30249 10180 30280
rect 11517 30277 11529 30280
rect 11563 30308 11575 30311
rect 11698 30308 11704 30320
rect 11563 30280 11704 30308
rect 11563 30277 11575 30280
rect 11517 30271 11575 30277
rect 11698 30268 11704 30280
rect 11756 30268 11762 30320
rect 11974 30268 11980 30320
rect 12032 30308 12038 30320
rect 12069 30311 12127 30317
rect 12069 30308 12081 30311
rect 12032 30280 12081 30308
rect 12032 30268 12038 30280
rect 12069 30277 12081 30280
rect 12115 30277 12127 30311
rect 14573 30308 14601 30348
rect 14734 30336 14740 30348
rect 14792 30336 14798 30388
rect 15194 30336 15200 30388
rect 15252 30376 15258 30388
rect 15252 30348 16988 30376
rect 15252 30336 15258 30348
rect 14642 30308 14648 30320
rect 14555 30280 14648 30308
rect 12069 30271 12127 30277
rect 14642 30268 14648 30280
rect 14700 30308 14706 30320
rect 16850 30308 16856 30320
rect 14700 30280 16856 30308
rect 14700 30268 14706 30280
rect 2665 30243 2723 30249
rect 2665 30240 2677 30243
rect 2556 30212 2677 30240
rect 2556 30200 2562 30212
rect 2665 30209 2677 30212
rect 2711 30209 2723 30243
rect 2665 30203 2723 30209
rect 10137 30243 10195 30249
rect 10137 30209 10149 30243
rect 10183 30209 10195 30243
rect 10137 30203 10195 30209
rect 10229 30243 10287 30249
rect 10229 30209 10241 30243
rect 10275 30209 10287 30243
rect 10229 30203 10287 30209
rect 9306 30132 9312 30184
rect 9364 30172 9370 30184
rect 10244 30172 10272 30203
rect 10318 30200 10324 30252
rect 10376 30240 10382 30252
rect 10505 30243 10563 30249
rect 10376 30212 10421 30240
rect 10376 30200 10382 30212
rect 10505 30209 10517 30243
rect 10551 30209 10563 30243
rect 10505 30203 10563 30209
rect 9364 30144 10272 30172
rect 10520 30172 10548 30203
rect 10962 30200 10968 30252
rect 11020 30240 11026 30252
rect 12253 30243 12311 30249
rect 12253 30240 12265 30243
rect 11020 30212 12265 30240
rect 11020 30200 11026 30212
rect 12253 30209 12265 30212
rect 12299 30240 12311 30243
rect 14826 30240 14832 30252
rect 12299 30212 14832 30240
rect 12299 30209 12311 30212
rect 12253 30203 12311 30209
rect 14826 30200 14832 30212
rect 14884 30200 14890 30252
rect 15010 30240 15016 30252
rect 14971 30212 15016 30240
rect 15010 30200 15016 30212
rect 15068 30200 15074 30252
rect 15120 30249 15148 30280
rect 16850 30268 16856 30280
rect 16908 30268 16914 30320
rect 15105 30243 15163 30249
rect 15105 30209 15117 30243
rect 15151 30209 15163 30243
rect 15105 30203 15163 30209
rect 15197 30243 15255 30249
rect 15197 30209 15209 30243
rect 15243 30240 15255 30243
rect 15286 30240 15292 30252
rect 15243 30212 15292 30240
rect 15243 30209 15255 30212
rect 15197 30203 15255 30209
rect 15286 30200 15292 30212
rect 15344 30200 15350 30252
rect 15378 30200 15384 30252
rect 15436 30240 15442 30252
rect 16666 30240 16672 30252
rect 15436 30212 16672 30240
rect 15436 30200 15442 30212
rect 16666 30200 16672 30212
rect 16724 30200 16730 30252
rect 16960 30249 16988 30348
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 19797 30379 19855 30385
rect 19797 30376 19809 30379
rect 19484 30348 19809 30376
rect 19484 30336 19490 30348
rect 19797 30345 19809 30348
rect 19843 30345 19855 30379
rect 29454 30376 29460 30388
rect 29415 30348 29460 30376
rect 19797 30339 19855 30345
rect 29454 30336 29460 30348
rect 29512 30376 29518 30388
rect 35897 30379 35955 30385
rect 29512 30348 30512 30376
rect 29512 30336 29518 30348
rect 18046 30268 18052 30320
rect 18104 30308 18110 30320
rect 18202 30311 18260 30317
rect 18202 30308 18214 30311
rect 18104 30280 18214 30308
rect 18104 30268 18110 30280
rect 18202 30277 18214 30280
rect 18248 30277 18260 30311
rect 18202 30271 18260 30277
rect 18874 30268 18880 30320
rect 18932 30308 18938 30320
rect 21174 30308 21180 30320
rect 18932 30280 20484 30308
rect 21135 30280 21180 30308
rect 18932 30268 18938 30280
rect 16945 30243 17003 30249
rect 16945 30209 16957 30243
rect 16991 30209 17003 30243
rect 16945 30203 17003 30209
rect 19242 30200 19248 30252
rect 19300 30240 19306 30252
rect 20073 30243 20131 30249
rect 20073 30240 20085 30243
rect 19300 30212 20085 30240
rect 19300 30200 19306 30212
rect 20073 30209 20085 30212
rect 20119 30209 20131 30243
rect 20073 30203 20131 30209
rect 20165 30243 20223 30249
rect 20165 30209 20177 30243
rect 20211 30209 20223 30243
rect 20165 30203 20223 30209
rect 11054 30172 11060 30184
rect 10520 30144 11060 30172
rect 9364 30132 9370 30144
rect 11054 30132 11060 30144
rect 11112 30132 11118 30184
rect 12437 30175 12495 30181
rect 12437 30141 12449 30175
rect 12483 30172 12495 30175
rect 12989 30175 13047 30181
rect 12989 30172 13001 30175
rect 12483 30144 13001 30172
rect 12483 30141 12495 30144
rect 12437 30135 12495 30141
rect 12989 30141 13001 30144
rect 13035 30172 13047 30175
rect 15838 30172 15844 30184
rect 13035 30144 15844 30172
rect 13035 30141 13047 30144
rect 12989 30135 13047 30141
rect 12452 30104 12480 30135
rect 15838 30132 15844 30144
rect 15896 30132 15902 30184
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 16761 30175 16819 30181
rect 16761 30172 16773 30175
rect 16632 30144 16773 30172
rect 16632 30132 16638 30144
rect 16761 30141 16773 30144
rect 16807 30141 16819 30175
rect 17954 30172 17960 30184
rect 17915 30144 17960 30172
rect 16761 30135 16819 30141
rect 17954 30132 17960 30144
rect 18012 30132 18018 30184
rect 20180 30172 20208 30203
rect 20254 30200 20260 30252
rect 20312 30240 20318 30252
rect 20456 30249 20484 30280
rect 21174 30268 21180 30280
rect 21232 30268 21238 30320
rect 22465 30311 22523 30317
rect 22465 30277 22477 30311
rect 22511 30308 22523 30311
rect 23750 30308 23756 30320
rect 22511 30280 23756 30308
rect 22511 30277 22523 30280
rect 22465 30271 22523 30277
rect 23750 30268 23756 30280
rect 23808 30268 23814 30320
rect 23845 30311 23903 30317
rect 23845 30277 23857 30311
rect 23891 30308 23903 30311
rect 25130 30308 25136 30320
rect 23891 30280 25136 30308
rect 23891 30277 23903 30280
rect 23845 30271 23903 30277
rect 20441 30243 20499 30249
rect 20312 30212 20357 30240
rect 20312 30200 20318 30212
rect 20441 30209 20453 30243
rect 20487 30209 20499 30243
rect 20441 30203 20499 30209
rect 20993 30243 21051 30249
rect 20993 30209 21005 30243
rect 21039 30209 21051 30243
rect 20993 30203 21051 30209
rect 20346 30172 20352 30184
rect 20180 30144 20352 30172
rect 20346 30132 20352 30144
rect 20404 30172 20410 30184
rect 21008 30172 21036 30203
rect 22186 30200 22192 30252
rect 22244 30240 22250 30252
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 22244 30212 22385 30240
rect 22244 30200 22250 30212
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 22554 30200 22560 30252
rect 22612 30240 22618 30252
rect 22741 30243 22799 30249
rect 22612 30212 22657 30240
rect 22612 30200 22618 30212
rect 22741 30209 22753 30243
rect 22787 30240 22799 30243
rect 23198 30240 23204 30252
rect 22787 30212 23204 30240
rect 22787 30209 22799 30212
rect 22741 30203 22799 30209
rect 23198 30200 23204 30212
rect 23256 30200 23262 30252
rect 23658 30240 23664 30252
rect 23619 30212 23664 30240
rect 23658 30200 23664 30212
rect 23716 30200 23722 30252
rect 20404 30144 21036 30172
rect 20404 30132 20410 30144
rect 23474 30132 23480 30184
rect 23532 30172 23538 30184
rect 23860 30172 23888 30271
rect 25130 30268 25136 30280
rect 25188 30268 25194 30320
rect 25225 30311 25283 30317
rect 25225 30277 25237 30311
rect 25271 30308 25283 30311
rect 26234 30308 26240 30320
rect 25271 30280 26240 30308
rect 25271 30277 25283 30280
rect 25225 30271 25283 30277
rect 26234 30268 26240 30280
rect 26292 30268 26298 30320
rect 26973 30311 27031 30317
rect 26973 30277 26985 30311
rect 27019 30308 27031 30311
rect 29914 30308 29920 30320
rect 27019 30280 29920 30308
rect 27019 30277 27031 30280
rect 26973 30271 27031 30277
rect 24210 30200 24216 30252
rect 24268 30240 24274 30252
rect 24578 30240 24584 30252
rect 24268 30212 24584 30240
rect 24268 30200 24274 30212
rect 24578 30200 24584 30212
rect 24636 30200 24642 30252
rect 24765 30243 24823 30249
rect 24765 30209 24777 30243
rect 24811 30209 24823 30243
rect 24765 30203 24823 30209
rect 24857 30243 24915 30249
rect 24857 30209 24869 30243
rect 24903 30209 24915 30243
rect 24857 30203 24915 30209
rect 24995 30243 25053 30249
rect 24995 30209 25007 30243
rect 25041 30209 25053 30243
rect 25682 30240 25688 30252
rect 25595 30212 25688 30240
rect 24995 30203 25053 30209
rect 23532 30144 23888 30172
rect 24029 30175 24087 30181
rect 23532 30132 23538 30144
rect 24029 30141 24041 30175
rect 24075 30172 24087 30175
rect 24780 30172 24808 30203
rect 24075 30144 24808 30172
rect 24075 30141 24087 30144
rect 24029 30135 24087 30141
rect 11164 30076 12480 30104
rect 3694 29996 3700 30048
rect 3752 30036 3758 30048
rect 3789 30039 3847 30045
rect 3789 30036 3801 30039
rect 3752 30008 3801 30036
rect 3752 29996 3758 30008
rect 3789 30005 3801 30008
rect 3835 30005 3847 30039
rect 3789 29999 3847 30005
rect 9306 29996 9312 30048
rect 9364 30036 9370 30048
rect 9401 30039 9459 30045
rect 9401 30036 9413 30039
rect 9364 30008 9413 30036
rect 9364 29996 9370 30008
rect 9401 30005 9413 30008
rect 9447 30036 9459 30039
rect 11164 30036 11192 30076
rect 24394 30064 24400 30116
rect 24452 30104 24458 30116
rect 24872 30104 24900 30203
rect 25010 30172 25038 30203
rect 25682 30200 25688 30212
rect 25740 30240 25746 30252
rect 26988 30240 27016 30271
rect 29914 30268 29920 30280
rect 29972 30268 29978 30320
rect 30193 30311 30251 30317
rect 30193 30277 30205 30311
rect 30239 30308 30251 30311
rect 30374 30308 30380 30320
rect 30239 30280 30380 30308
rect 30239 30277 30251 30280
rect 30193 30271 30251 30277
rect 30374 30268 30380 30280
rect 30432 30268 30438 30320
rect 25740 30212 27016 30240
rect 25740 30200 25746 30212
rect 27062 30200 27068 30252
rect 27120 30240 27126 30252
rect 28350 30249 28356 30252
rect 28077 30243 28135 30249
rect 28077 30240 28089 30243
rect 27120 30212 28089 30240
rect 27120 30200 27126 30212
rect 28077 30209 28089 30212
rect 28123 30209 28135 30243
rect 28344 30240 28356 30249
rect 28311 30212 28356 30240
rect 28077 30203 28135 30209
rect 28344 30203 28356 30212
rect 28350 30200 28356 30203
rect 28408 30200 28414 30252
rect 30098 30240 30104 30252
rect 30059 30212 30104 30240
rect 30098 30200 30104 30212
rect 30156 30200 30162 30252
rect 30484 30249 30512 30348
rect 32692 30348 34514 30376
rect 31202 30268 31208 30320
rect 31260 30308 31266 30320
rect 32582 30308 32588 30320
rect 31260 30280 32588 30308
rect 31260 30268 31266 30280
rect 32582 30268 32588 30280
rect 32640 30268 32646 30320
rect 32692 30317 32720 30348
rect 32677 30311 32735 30317
rect 32677 30277 32689 30311
rect 32723 30277 32735 30311
rect 33686 30308 33692 30320
rect 33647 30280 33692 30308
rect 32677 30271 32735 30277
rect 33686 30268 33692 30280
rect 33744 30268 33750 30320
rect 34486 30308 34514 30348
rect 35897 30345 35909 30379
rect 35943 30376 35955 30379
rect 35986 30376 35992 30388
rect 35943 30348 35992 30376
rect 35943 30345 35955 30348
rect 35897 30339 35955 30345
rect 35986 30336 35992 30348
rect 36044 30336 36050 30388
rect 35713 30311 35771 30317
rect 35713 30308 35725 30311
rect 34486 30280 35725 30308
rect 35713 30277 35725 30280
rect 35759 30308 35771 30311
rect 37366 30308 37372 30320
rect 35759 30280 37372 30308
rect 35759 30277 35771 30280
rect 35713 30271 35771 30277
rect 37366 30268 37372 30280
rect 37424 30268 37430 30320
rect 30285 30243 30343 30249
rect 30285 30209 30297 30243
rect 30331 30209 30343 30243
rect 30285 30203 30343 30209
rect 30469 30243 30527 30249
rect 30469 30209 30481 30243
rect 30515 30209 30527 30243
rect 30469 30203 30527 30209
rect 32401 30243 32459 30249
rect 32401 30209 32413 30243
rect 32447 30209 32459 30243
rect 32401 30203 32459 30209
rect 32769 30243 32827 30249
rect 32769 30209 32781 30243
rect 32815 30240 32827 30243
rect 33134 30240 33140 30252
rect 32815 30212 33140 30240
rect 32815 30209 32827 30212
rect 32769 30203 32827 30209
rect 30300 30172 30328 30203
rect 30558 30172 30564 30184
rect 25010 30144 26004 30172
rect 30300 30144 30564 30172
rect 25010 30116 25038 30144
rect 24452 30076 24900 30104
rect 24452 30064 24458 30076
rect 24946 30064 24952 30116
rect 25004 30076 25038 30116
rect 25004 30064 25010 30076
rect 9447 30008 11192 30036
rect 9447 30005 9459 30008
rect 9401 29999 9459 30005
rect 11698 29996 11704 30048
rect 11756 30036 11762 30048
rect 12894 30036 12900 30048
rect 11756 30008 12900 30036
rect 11756 29996 11762 30008
rect 12894 29996 12900 30008
rect 12952 30036 12958 30048
rect 13170 30036 13176 30048
rect 12952 30008 13176 30036
rect 12952 29996 12958 30008
rect 13170 29996 13176 30008
rect 13228 29996 13234 30048
rect 15010 29996 15016 30048
rect 15068 30036 15074 30048
rect 15930 30036 15936 30048
rect 15068 30008 15936 30036
rect 15068 29996 15074 30008
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 17126 30036 17132 30048
rect 17087 30008 17132 30036
rect 17126 29996 17132 30008
rect 17184 29996 17190 30048
rect 19334 30036 19340 30048
rect 19295 30008 19340 30036
rect 19334 29996 19340 30008
rect 19392 29996 19398 30048
rect 22189 30039 22247 30045
rect 22189 30005 22201 30039
rect 22235 30036 22247 30039
rect 22370 30036 22376 30048
rect 22235 30008 22376 30036
rect 22235 30005 22247 30008
rect 22189 29999 22247 30005
rect 22370 29996 22376 30008
rect 22428 29996 22434 30048
rect 25866 30036 25872 30048
rect 25827 30008 25872 30036
rect 25866 29996 25872 30008
rect 25924 29996 25930 30048
rect 25976 30036 26004 30144
rect 30558 30132 30564 30144
rect 30616 30132 30622 30184
rect 32416 30172 32444 30203
rect 33134 30200 33140 30212
rect 33192 30240 33198 30252
rect 33502 30240 33508 30252
rect 33192 30212 33508 30240
rect 33192 30200 33198 30212
rect 33502 30200 33508 30212
rect 33560 30240 33566 30252
rect 33597 30243 33655 30249
rect 33597 30240 33609 30243
rect 33560 30212 33609 30240
rect 33560 30200 33566 30212
rect 33597 30209 33609 30212
rect 33643 30209 33655 30243
rect 33597 30203 33655 30209
rect 33781 30243 33839 30249
rect 33781 30209 33793 30243
rect 33827 30240 33839 30243
rect 33870 30240 33876 30252
rect 33827 30212 33876 30240
rect 33827 30209 33839 30212
rect 33781 30203 33839 30209
rect 33870 30200 33876 30212
rect 33928 30200 33934 30252
rect 33965 30243 34023 30249
rect 33965 30209 33977 30243
rect 34011 30240 34023 30243
rect 34054 30240 34060 30252
rect 34011 30212 34060 30240
rect 34011 30209 34023 30212
rect 33965 30203 34023 30209
rect 34054 30200 34060 30212
rect 34112 30200 34118 30252
rect 35526 30240 35532 30252
rect 35487 30212 35532 30240
rect 35526 30200 35532 30212
rect 35584 30200 35590 30252
rect 34790 30172 34796 30184
rect 32416 30144 34796 30172
rect 34790 30132 34796 30144
rect 34848 30132 34854 30184
rect 32858 30104 32864 30116
rect 29012 30076 32864 30104
rect 29012 30036 29040 30076
rect 32858 30064 32864 30076
rect 32916 30064 32922 30116
rect 33686 30064 33692 30116
rect 33744 30104 33750 30116
rect 35434 30104 35440 30116
rect 33744 30076 35440 30104
rect 33744 30064 33750 30076
rect 35434 30064 35440 30076
rect 35492 30064 35498 30116
rect 25976 30008 29040 30036
rect 29270 29996 29276 30048
rect 29328 30036 29334 30048
rect 29917 30039 29975 30045
rect 29917 30036 29929 30039
rect 29328 30008 29929 30036
rect 29328 29996 29334 30008
rect 29917 30005 29929 30008
rect 29963 30005 29975 30039
rect 29917 29999 29975 30005
rect 30650 29996 30656 30048
rect 30708 30036 30714 30048
rect 31205 30039 31263 30045
rect 31205 30036 31217 30039
rect 30708 30008 31217 30036
rect 30708 29996 30714 30008
rect 31205 30005 31217 30008
rect 31251 30036 31263 30039
rect 31386 30036 31392 30048
rect 31251 30008 31392 30036
rect 31251 30005 31263 30008
rect 31205 29999 31263 30005
rect 31386 29996 31392 30008
rect 31444 29996 31450 30048
rect 32953 30039 33011 30045
rect 32953 30005 32965 30039
rect 32999 30036 33011 30039
rect 33318 30036 33324 30048
rect 32999 30008 33324 30036
rect 32999 30005 33011 30008
rect 32953 29999 33011 30005
rect 33318 29996 33324 30008
rect 33376 29996 33382 30048
rect 33413 30039 33471 30045
rect 33413 30005 33425 30039
rect 33459 30036 33471 30039
rect 33870 30036 33876 30048
rect 33459 30008 33876 30036
rect 33459 30005 33471 30008
rect 33413 29999 33471 30005
rect 33870 29996 33876 30008
rect 33928 29996 33934 30048
rect 36630 30036 36636 30048
rect 36591 30008 36636 30036
rect 36630 29996 36636 30008
rect 36688 29996 36694 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 2225 29835 2283 29841
rect 2225 29801 2237 29835
rect 2271 29832 2283 29835
rect 2498 29832 2504 29844
rect 2271 29804 2504 29832
rect 2271 29801 2283 29804
rect 2225 29795 2283 29801
rect 2498 29792 2504 29804
rect 2556 29792 2562 29844
rect 8202 29792 8208 29844
rect 8260 29832 8266 29844
rect 8941 29835 8999 29841
rect 8941 29832 8953 29835
rect 8260 29804 8953 29832
rect 8260 29792 8266 29804
rect 8941 29801 8953 29804
rect 8987 29801 8999 29835
rect 12986 29832 12992 29844
rect 8941 29795 8999 29801
rect 9048 29804 12992 29832
rect 2958 29764 2964 29776
rect 2470 29736 2964 29764
rect 2470 29637 2498 29736
rect 2958 29724 2964 29736
rect 3016 29764 3022 29776
rect 3789 29767 3847 29773
rect 3789 29764 3801 29767
rect 3016 29736 3801 29764
rect 3016 29724 3022 29736
rect 3789 29733 3801 29736
rect 3835 29733 3847 29767
rect 3789 29727 3847 29733
rect 7466 29724 7472 29776
rect 7524 29764 7530 29776
rect 7742 29764 7748 29776
rect 7524 29736 7748 29764
rect 7524 29724 7530 29736
rect 7742 29724 7748 29736
rect 7800 29764 7806 29776
rect 9048 29764 9076 29804
rect 12986 29792 12992 29804
rect 13044 29792 13050 29844
rect 18506 29792 18512 29844
rect 18564 29832 18570 29844
rect 18693 29835 18751 29841
rect 18693 29832 18705 29835
rect 18564 29804 18705 29832
rect 18564 29792 18570 29804
rect 18693 29801 18705 29804
rect 18739 29801 18751 29835
rect 20254 29832 20260 29844
rect 20215 29804 20260 29832
rect 18693 29795 18751 29801
rect 20254 29792 20260 29804
rect 20312 29792 20318 29844
rect 23845 29835 23903 29841
rect 23845 29832 23857 29835
rect 23446 29804 23857 29832
rect 7800 29736 9076 29764
rect 7800 29724 7806 29736
rect 15930 29724 15936 29776
rect 15988 29764 15994 29776
rect 23446 29764 23474 29804
rect 23845 29801 23857 29804
rect 23891 29832 23903 29835
rect 24946 29832 24952 29844
rect 23891 29804 24952 29832
rect 23891 29801 23903 29804
rect 23845 29795 23903 29801
rect 24946 29792 24952 29804
rect 25004 29792 25010 29844
rect 26326 29832 26332 29844
rect 25056 29804 26332 29832
rect 15988 29736 23474 29764
rect 24489 29767 24547 29773
rect 15988 29724 15994 29736
rect 24489 29733 24501 29767
rect 24535 29764 24547 29767
rect 24670 29764 24676 29776
rect 24535 29736 24676 29764
rect 24535 29733 24547 29736
rect 24489 29727 24547 29733
rect 24670 29724 24676 29736
rect 24728 29724 24734 29776
rect 3326 29656 3332 29708
rect 3384 29696 3390 29708
rect 9306 29696 9312 29708
rect 3384 29668 4660 29696
rect 9267 29668 9312 29696
rect 3384 29656 3390 29668
rect 2455 29631 2513 29637
rect 2455 29597 2467 29631
rect 2501 29597 2513 29631
rect 2590 29628 2596 29640
rect 2551 29600 2596 29628
rect 2455 29591 2513 29597
rect 2590 29588 2596 29600
rect 2648 29588 2654 29640
rect 2685 29631 2743 29637
rect 2685 29597 2697 29631
rect 2731 29597 2743 29631
rect 2685 29591 2743 29597
rect 2700 29504 2728 29591
rect 2866 29588 2872 29640
rect 2924 29628 2930 29640
rect 2924 29600 2969 29628
rect 2924 29588 2930 29600
rect 3418 29588 3424 29640
rect 3476 29628 3482 29640
rect 4632 29637 4660 29668
rect 9306 29656 9312 29668
rect 9364 29656 9370 29708
rect 16574 29656 16580 29708
rect 16632 29696 16638 29708
rect 24118 29696 24124 29708
rect 16632 29668 24124 29696
rect 16632 29656 16638 29668
rect 24118 29656 24124 29668
rect 24176 29656 24182 29708
rect 25056 29696 25084 29804
rect 26326 29792 26332 29804
rect 26384 29792 26390 29844
rect 29822 29832 29828 29844
rect 29783 29804 29828 29832
rect 29822 29792 29828 29804
rect 29880 29792 29886 29844
rect 31478 29792 31484 29844
rect 31536 29832 31542 29844
rect 36630 29832 36636 29844
rect 31536 29804 36636 29832
rect 31536 29792 31542 29804
rect 36630 29792 36636 29804
rect 36688 29792 36694 29844
rect 30834 29724 30840 29776
rect 30892 29724 30898 29776
rect 36648 29764 36676 29792
rect 36648 29736 37228 29764
rect 24412 29668 25084 29696
rect 26605 29699 26663 29705
rect 4341 29631 4399 29637
rect 4341 29628 4353 29631
rect 3476 29600 4353 29628
rect 3476 29588 3482 29600
rect 4341 29597 4353 29600
rect 4387 29597 4399 29631
rect 4341 29591 4399 29597
rect 4617 29631 4675 29637
rect 4617 29597 4629 29631
rect 4663 29597 4675 29631
rect 4617 29591 4675 29597
rect 4709 29631 4767 29637
rect 4709 29597 4721 29631
rect 4755 29628 4767 29631
rect 5166 29628 5172 29640
rect 4755 29600 5172 29628
rect 4755 29597 4767 29600
rect 4709 29591 4767 29597
rect 5166 29588 5172 29600
rect 5224 29588 5230 29640
rect 9125 29631 9183 29637
rect 9125 29597 9137 29631
rect 9171 29628 9183 29631
rect 9490 29628 9496 29640
rect 9171 29600 9496 29628
rect 9171 29597 9183 29600
rect 9125 29591 9183 29597
rect 9490 29588 9496 29600
rect 9548 29588 9554 29640
rect 10502 29628 10508 29640
rect 10463 29600 10508 29628
rect 10502 29588 10508 29600
rect 10560 29588 10566 29640
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29628 18567 29631
rect 19334 29628 19340 29640
rect 18555 29600 19340 29628
rect 18555 29597 18567 29600
rect 18509 29591 18567 29597
rect 19334 29588 19340 29600
rect 19392 29588 19398 29640
rect 19978 29628 19984 29640
rect 19891 29600 19984 29628
rect 10778 29569 10784 29572
rect 4525 29563 4583 29569
rect 4525 29529 4537 29563
rect 4571 29529 4583 29563
rect 4525 29523 4583 29529
rect 10772 29523 10784 29569
rect 10836 29560 10842 29572
rect 10836 29532 10872 29560
rect 2682 29452 2688 29504
rect 2740 29452 2746 29504
rect 4540 29492 4568 29523
rect 10778 29520 10784 29523
rect 10836 29520 10842 29532
rect 15746 29520 15752 29572
rect 15804 29560 15810 29572
rect 19904 29569 19932 29600
rect 19978 29588 19984 29600
rect 20036 29628 20042 29640
rect 21269 29631 21327 29637
rect 21269 29628 21281 29631
rect 20036 29600 21281 29628
rect 20036 29588 20042 29600
rect 21269 29597 21281 29600
rect 21315 29597 21327 29631
rect 21269 29591 21327 29597
rect 22186 29588 22192 29640
rect 22244 29628 22250 29640
rect 22373 29631 22431 29637
rect 22373 29628 22385 29631
rect 22244 29600 22385 29628
rect 22244 29588 22250 29600
rect 22373 29597 22385 29600
rect 22419 29597 22431 29631
rect 22554 29628 22560 29640
rect 22515 29600 22560 29628
rect 22373 29591 22431 29597
rect 22554 29588 22560 29600
rect 22612 29588 22618 29640
rect 22738 29628 22744 29640
rect 22699 29600 22744 29628
rect 22738 29588 22744 29600
rect 22796 29588 22802 29640
rect 17773 29563 17831 29569
rect 17773 29560 17785 29563
rect 15804 29532 17785 29560
rect 15804 29520 15810 29532
rect 17773 29529 17785 29532
rect 17819 29560 17831 29563
rect 18325 29563 18383 29569
rect 18325 29560 18337 29563
rect 17819 29532 18337 29560
rect 17819 29529 17831 29532
rect 17773 29523 17831 29529
rect 18325 29529 18337 29532
rect 18371 29560 18383 29563
rect 19889 29563 19947 29569
rect 19889 29560 19901 29563
rect 18371 29532 19901 29560
rect 18371 29529 18383 29532
rect 18325 29523 18383 29529
rect 19889 29529 19901 29532
rect 19935 29529 19947 29563
rect 20070 29560 20076 29572
rect 20031 29532 20076 29560
rect 19889 29523 19947 29529
rect 20070 29520 20076 29532
rect 20128 29520 20134 29572
rect 22465 29563 22523 29569
rect 22465 29529 22477 29563
rect 22511 29560 22523 29563
rect 24412 29560 24440 29668
rect 26605 29665 26617 29699
rect 26651 29696 26663 29699
rect 27062 29696 27068 29708
rect 26651 29668 27068 29696
rect 26651 29665 26663 29668
rect 26605 29659 26663 29665
rect 27062 29656 27068 29668
rect 27120 29656 27126 29708
rect 30852 29696 30880 29724
rect 35805 29699 35863 29705
rect 30852 29668 31156 29696
rect 24673 29631 24731 29637
rect 24673 29597 24685 29631
rect 24719 29628 24731 29631
rect 24719 29600 25452 29628
rect 24719 29597 24731 29600
rect 24673 29591 24731 29597
rect 24688 29560 24716 29591
rect 22511 29532 24440 29560
rect 24504 29532 24716 29560
rect 22511 29529 22523 29532
rect 22465 29523 22523 29529
rect 4706 29492 4712 29504
rect 4540 29464 4712 29492
rect 4706 29452 4712 29464
rect 4764 29452 4770 29504
rect 4798 29452 4804 29504
rect 4856 29492 4862 29504
rect 4893 29495 4951 29501
rect 4893 29492 4905 29495
rect 4856 29464 4905 29492
rect 4856 29452 4862 29464
rect 4893 29461 4905 29464
rect 4939 29461 4951 29495
rect 4893 29455 4951 29461
rect 7742 29452 7748 29504
rect 7800 29492 7806 29504
rect 7837 29495 7895 29501
rect 7837 29492 7849 29495
rect 7800 29464 7849 29492
rect 7800 29452 7806 29464
rect 7837 29461 7849 29464
rect 7883 29461 7895 29495
rect 7837 29455 7895 29461
rect 9766 29452 9772 29504
rect 9824 29492 9830 29504
rect 10045 29495 10103 29501
rect 10045 29492 10057 29495
rect 9824 29464 10057 29492
rect 9824 29452 9830 29464
rect 10045 29461 10057 29464
rect 10091 29492 10103 29495
rect 11054 29492 11060 29504
rect 10091 29464 11060 29492
rect 10091 29461 10103 29464
rect 10045 29455 10103 29461
rect 11054 29452 11060 29464
rect 11112 29452 11118 29504
rect 11698 29452 11704 29504
rect 11756 29492 11762 29504
rect 11885 29495 11943 29501
rect 11885 29492 11897 29495
rect 11756 29464 11897 29492
rect 11756 29452 11762 29464
rect 11885 29461 11897 29464
rect 11931 29461 11943 29495
rect 16574 29492 16580 29504
rect 16535 29464 16580 29492
rect 11885 29455 11943 29461
rect 16574 29452 16580 29464
rect 16632 29452 16638 29504
rect 16942 29452 16948 29504
rect 17000 29492 17006 29504
rect 19337 29495 19395 29501
rect 19337 29492 19349 29495
rect 17000 29464 19349 29492
rect 17000 29452 17006 29464
rect 19337 29461 19349 29464
rect 19383 29492 19395 29495
rect 20346 29492 20352 29504
rect 19383 29464 20352 29492
rect 19383 29461 19395 29464
rect 19337 29455 19395 29461
rect 20346 29452 20352 29464
rect 20404 29492 20410 29504
rect 20717 29495 20775 29501
rect 20717 29492 20729 29495
rect 20404 29464 20729 29492
rect 20404 29452 20410 29464
rect 20717 29461 20729 29464
rect 20763 29461 20775 29495
rect 20717 29455 20775 29461
rect 22189 29495 22247 29501
rect 22189 29461 22201 29495
rect 22235 29492 22247 29495
rect 23014 29492 23020 29504
rect 22235 29464 23020 29492
rect 22235 29461 22247 29464
rect 22189 29455 22247 29461
rect 23014 29452 23020 29464
rect 23072 29452 23078 29504
rect 23293 29495 23351 29501
rect 23293 29461 23305 29495
rect 23339 29492 23351 29495
rect 24504 29492 24532 29532
rect 23339 29464 24532 29492
rect 23339 29461 23351 29464
rect 23293 29455 23351 29461
rect 24578 29452 24584 29504
rect 24636 29492 24642 29504
rect 25225 29495 25283 29501
rect 25225 29492 25237 29495
rect 24636 29464 25237 29492
rect 24636 29452 24642 29464
rect 25225 29461 25237 29464
rect 25271 29461 25283 29495
rect 25424 29492 25452 29600
rect 29822 29588 29828 29640
rect 29880 29628 29886 29640
rect 31128 29637 31156 29668
rect 31772 29668 32076 29696
rect 30837 29631 30895 29637
rect 30837 29628 30849 29631
rect 29880 29600 30849 29628
rect 29880 29588 29886 29600
rect 30837 29597 30849 29600
rect 30883 29597 30895 29631
rect 31000 29631 31058 29637
rect 31000 29628 31012 29631
rect 30837 29591 30895 29597
rect 30944 29600 31012 29628
rect 25590 29520 25596 29572
rect 25648 29560 25654 29572
rect 26338 29563 26396 29569
rect 26338 29560 26350 29563
rect 25648 29532 26350 29560
rect 25648 29520 25654 29532
rect 26338 29529 26350 29532
rect 26384 29529 26396 29563
rect 30944 29560 30972 29600
rect 31000 29597 31012 29600
rect 31046 29597 31058 29631
rect 31000 29591 31058 29597
rect 31113 29631 31171 29637
rect 31113 29597 31125 29631
rect 31159 29597 31171 29631
rect 31113 29591 31171 29597
rect 31202 29588 31208 29640
rect 31260 29628 31266 29640
rect 31772 29628 31800 29668
rect 31938 29628 31944 29640
rect 31260 29600 31305 29628
rect 31404 29600 31800 29628
rect 31899 29600 31944 29628
rect 31260 29588 31266 29600
rect 31404 29560 31432 29600
rect 31938 29588 31944 29600
rect 31996 29588 32002 29640
rect 32048 29628 32076 29668
rect 35805 29665 35817 29699
rect 35851 29696 35863 29699
rect 36354 29696 36360 29708
rect 35851 29668 36360 29696
rect 35851 29665 35863 29668
rect 35805 29659 35863 29665
rect 36354 29656 36360 29668
rect 36412 29696 36418 29708
rect 36412 29668 37136 29696
rect 36412 29656 36418 29668
rect 34149 29631 34207 29637
rect 34149 29628 34161 29631
rect 32048 29600 34161 29628
rect 34149 29597 34161 29600
rect 34195 29597 34207 29631
rect 34149 29591 34207 29597
rect 34606 29588 34612 29640
rect 34664 29628 34670 29640
rect 34701 29631 34759 29637
rect 34701 29628 34713 29631
rect 34664 29600 34713 29628
rect 34664 29588 34670 29600
rect 34701 29597 34713 29600
rect 34747 29597 34759 29631
rect 34701 29591 34759 29597
rect 35529 29631 35587 29637
rect 35529 29597 35541 29631
rect 35575 29628 35587 29631
rect 35618 29628 35624 29640
rect 35575 29600 35624 29628
rect 35575 29597 35587 29600
rect 35529 29591 35587 29597
rect 35618 29588 35624 29600
rect 35676 29588 35682 29640
rect 36078 29588 36084 29640
rect 36136 29628 36142 29640
rect 36817 29631 36875 29637
rect 36817 29628 36829 29631
rect 36136 29600 36829 29628
rect 36136 29588 36142 29600
rect 36817 29597 36829 29600
rect 36863 29597 36875 29631
rect 36998 29628 37004 29640
rect 36959 29600 37004 29628
rect 36817 29591 36875 29597
rect 36998 29588 37004 29600
rect 37056 29588 37062 29640
rect 37108 29637 37136 29668
rect 37200 29637 37228 29736
rect 37093 29631 37151 29637
rect 37093 29597 37105 29631
rect 37139 29597 37151 29631
rect 37093 29591 37151 29597
rect 37185 29631 37243 29637
rect 37185 29597 37197 29631
rect 37231 29597 37243 29631
rect 58158 29628 58164 29640
rect 58119 29600 58164 29628
rect 37185 29591 37243 29597
rect 58158 29588 58164 29600
rect 58216 29588 58222 29640
rect 30944 29532 31432 29560
rect 31481 29563 31539 29569
rect 26338 29523 26396 29529
rect 31481 29529 31493 29563
rect 31527 29560 31539 29563
rect 32186 29563 32244 29569
rect 32186 29560 32198 29563
rect 31527 29532 32198 29560
rect 31527 29529 31539 29532
rect 31481 29523 31539 29529
rect 32186 29529 32198 29532
rect 32232 29529 32244 29563
rect 32186 29523 32244 29529
rect 32306 29520 32312 29572
rect 32364 29560 32370 29572
rect 33781 29563 33839 29569
rect 33781 29560 33793 29563
rect 32364 29532 33793 29560
rect 32364 29520 32370 29532
rect 33781 29529 33793 29532
rect 33827 29529 33839 29563
rect 33781 29523 33839 29529
rect 33965 29563 34023 29569
rect 33965 29529 33977 29563
rect 34011 29529 34023 29563
rect 33965 29523 34023 29529
rect 26418 29492 26424 29504
rect 25424 29464 26424 29492
rect 25225 29455 25283 29461
rect 26418 29452 26424 29464
rect 26476 29452 26482 29504
rect 30006 29452 30012 29504
rect 30064 29492 30070 29504
rect 30285 29495 30343 29501
rect 30285 29492 30297 29495
rect 30064 29464 30297 29492
rect 30064 29452 30070 29464
rect 30285 29461 30297 29464
rect 30331 29492 30343 29495
rect 31202 29492 31208 29504
rect 30331 29464 31208 29492
rect 30331 29461 30343 29464
rect 30285 29455 30343 29461
rect 31202 29452 31208 29464
rect 31260 29452 31266 29504
rect 33226 29452 33232 29504
rect 33284 29492 33290 29504
rect 33321 29495 33379 29501
rect 33321 29492 33333 29495
rect 33284 29464 33333 29492
rect 33284 29452 33290 29464
rect 33321 29461 33333 29464
rect 33367 29492 33379 29495
rect 33980 29492 34008 29523
rect 33367 29464 34008 29492
rect 34885 29495 34943 29501
rect 33367 29461 33379 29464
rect 33321 29455 33379 29461
rect 34885 29461 34897 29495
rect 34931 29492 34943 29495
rect 35526 29492 35532 29504
rect 34931 29464 35532 29492
rect 34931 29461 34943 29464
rect 34885 29455 34943 29461
rect 35526 29452 35532 29464
rect 35584 29452 35590 29504
rect 37458 29492 37464 29504
rect 37419 29464 37464 29492
rect 37458 29452 37464 29464
rect 37516 29452 37522 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 2866 29248 2872 29300
rect 2924 29288 2930 29300
rect 10134 29288 10140 29300
rect 2924 29260 10140 29288
rect 2924 29248 2930 29260
rect 2590 29180 2596 29232
rect 2648 29220 2654 29232
rect 2648 29192 3188 29220
rect 2648 29180 2654 29192
rect 3160 29161 3188 29192
rect 3053 29155 3111 29161
rect 2976 29127 3065 29155
rect 2777 28951 2835 28957
rect 2777 28917 2789 28951
rect 2823 28948 2835 28951
rect 2866 28948 2872 28960
rect 2823 28920 2872 28948
rect 2823 28917 2835 28920
rect 2777 28911 2835 28917
rect 2866 28908 2872 28920
rect 2924 28908 2930 28960
rect 2976 28948 3004 29127
rect 3053 29121 3065 29127
rect 3099 29121 3111 29155
rect 3053 29115 3111 29121
rect 3145 29155 3203 29161
rect 3145 29121 3157 29155
rect 3191 29121 3203 29155
rect 3145 29115 3203 29121
rect 3242 29155 3300 29161
rect 3242 29121 3254 29155
rect 3288 29152 3300 29155
rect 3421 29155 3479 29161
rect 3288 29124 3372 29152
rect 3288 29121 3300 29124
rect 3242 29115 3300 29121
rect 3344 29084 3372 29124
rect 3421 29121 3433 29155
rect 3467 29152 3479 29155
rect 3620 29152 3648 29260
rect 10134 29248 10140 29260
rect 10192 29248 10198 29300
rect 10410 29248 10416 29300
rect 10468 29248 10474 29300
rect 10778 29288 10784 29300
rect 10739 29260 10784 29288
rect 10778 29248 10784 29260
rect 10836 29248 10842 29300
rect 13722 29248 13728 29300
rect 13780 29288 13786 29300
rect 14369 29291 14427 29297
rect 14369 29288 14381 29291
rect 13780 29260 14381 29288
rect 13780 29248 13786 29260
rect 14369 29257 14381 29260
rect 14415 29257 14427 29291
rect 23474 29288 23480 29300
rect 14369 29251 14427 29257
rect 19996 29260 23480 29288
rect 4801 29223 4859 29229
rect 4801 29189 4813 29223
rect 4847 29220 4859 29223
rect 5074 29220 5080 29232
rect 4847 29192 5080 29220
rect 4847 29189 4859 29192
rect 4801 29183 4859 29189
rect 5074 29180 5080 29192
rect 5132 29180 5138 29232
rect 8202 29220 8208 29232
rect 8163 29192 8208 29220
rect 8202 29180 8208 29192
rect 8260 29180 8266 29232
rect 8570 29220 8576 29232
rect 8531 29192 8576 29220
rect 8570 29180 8576 29192
rect 8628 29180 8634 29232
rect 3467 29124 3648 29152
rect 3467 29121 3479 29124
rect 3421 29115 3479 29121
rect 3694 29112 3700 29164
rect 3752 29152 3758 29164
rect 4525 29155 4583 29161
rect 4525 29152 4537 29155
rect 3752 29124 4537 29152
rect 3752 29112 3758 29124
rect 4525 29121 4537 29124
rect 4571 29121 4583 29155
rect 4706 29152 4712 29164
rect 4667 29124 4712 29152
rect 4525 29115 4583 29121
rect 4706 29112 4712 29124
rect 4764 29112 4770 29164
rect 4893 29155 4951 29161
rect 4893 29121 4905 29155
rect 4939 29152 4951 29155
rect 5166 29152 5172 29164
rect 4939 29124 5172 29152
rect 4939 29121 4951 29124
rect 4893 29115 4951 29121
rect 5166 29112 5172 29124
rect 5224 29152 5230 29164
rect 7469 29155 7527 29161
rect 7469 29152 7481 29155
rect 5224 29124 7481 29152
rect 5224 29112 5230 29124
rect 7469 29121 7481 29124
rect 7515 29152 7527 29155
rect 7653 29155 7711 29161
rect 7515 29124 7604 29152
rect 7515 29121 7527 29124
rect 7469 29115 7527 29121
rect 3786 29084 3792 29096
rect 3344 29056 3792 29084
rect 3786 29044 3792 29056
rect 3844 29044 3850 29096
rect 4890 28976 4896 29028
rect 4948 29016 4954 29028
rect 5077 29019 5135 29025
rect 5077 29016 5089 29019
rect 4948 28988 5089 29016
rect 4948 28976 4954 28988
rect 5077 28985 5089 28988
rect 5123 28985 5135 29019
rect 7466 29016 7472 29028
rect 7427 28988 7472 29016
rect 5077 28979 5135 28985
rect 7466 28976 7472 28988
rect 7524 28976 7530 29028
rect 7576 29016 7604 29124
rect 7653 29121 7665 29155
rect 7699 29152 7711 29155
rect 7742 29152 7748 29164
rect 7699 29124 7748 29152
rect 7699 29121 7711 29124
rect 7653 29115 7711 29121
rect 7742 29112 7748 29124
rect 7800 29112 7806 29164
rect 8389 29155 8447 29161
rect 8389 29121 8401 29155
rect 8435 29152 8447 29155
rect 9122 29152 9128 29164
rect 8435 29124 9128 29152
rect 8435 29121 8447 29124
rect 8389 29115 8447 29121
rect 9122 29112 9128 29124
rect 9180 29112 9186 29164
rect 9214 29112 9220 29164
rect 9272 29161 9278 29164
rect 9382 29161 9440 29167
rect 9272 29155 9321 29161
rect 9272 29121 9275 29155
rect 9309 29121 9321 29155
rect 9382 29127 9394 29161
rect 9428 29158 9440 29161
rect 9428 29127 9444 29158
rect 9382 29121 9444 29127
rect 9272 29115 9321 29121
rect 9272 29112 9278 29115
rect 9416 29084 9444 29121
rect 9493 29155 9551 29161
rect 9493 29121 9505 29155
rect 9539 29152 9551 29155
rect 9582 29152 9588 29164
rect 9539 29124 9588 29152
rect 9539 29121 9551 29124
rect 9493 29115 9551 29121
rect 9582 29112 9588 29124
rect 9640 29112 9646 29164
rect 9677 29155 9735 29161
rect 9677 29121 9689 29155
rect 9723 29152 9735 29155
rect 9766 29152 9772 29164
rect 9723 29124 9772 29152
rect 9723 29121 9735 29124
rect 9677 29115 9735 29121
rect 9766 29112 9772 29124
rect 9824 29112 9830 29164
rect 10134 29152 10140 29164
rect 10095 29124 10140 29152
rect 10134 29112 10140 29124
rect 10192 29112 10198 29164
rect 10428 29161 10456 29248
rect 11698 29220 11704 29232
rect 11659 29192 11704 29220
rect 11698 29180 11704 29192
rect 11756 29220 11762 29232
rect 14182 29220 14188 29232
rect 11756 29192 14188 29220
rect 11756 29180 11762 29192
rect 14182 29180 14188 29192
rect 14240 29180 14246 29232
rect 15473 29223 15531 29229
rect 15473 29189 15485 29223
rect 15519 29220 15531 29223
rect 17126 29220 17132 29232
rect 15519 29192 17132 29220
rect 15519 29189 15531 29192
rect 15473 29183 15531 29189
rect 17126 29180 17132 29192
rect 17184 29180 17190 29232
rect 18506 29220 18512 29232
rect 17926 29192 18512 29220
rect 10321 29155 10379 29161
rect 10321 29121 10333 29155
rect 10367 29121 10379 29155
rect 10321 29115 10379 29121
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29121 10471 29155
rect 10413 29115 10471 29121
rect 10505 29155 10563 29161
rect 10505 29121 10517 29155
rect 10551 29152 10563 29155
rect 10778 29152 10784 29164
rect 10551 29124 10784 29152
rect 10551 29121 10563 29124
rect 10505 29115 10563 29121
rect 10336 29084 10364 29115
rect 10778 29112 10784 29124
rect 10836 29152 10842 29164
rect 11885 29155 11943 29161
rect 10836 29124 11652 29152
rect 10836 29112 10842 29124
rect 11517 29087 11575 29093
rect 11517 29084 11529 29087
rect 9416 29056 9490 29084
rect 10336 29056 11529 29084
rect 9462 29028 9490 29056
rect 11517 29053 11529 29056
rect 11563 29053 11575 29087
rect 11624 29084 11652 29124
rect 11885 29121 11897 29155
rect 11931 29152 11943 29155
rect 11974 29152 11980 29164
rect 11931 29124 11980 29152
rect 11931 29121 11943 29124
rect 11885 29115 11943 29121
rect 11974 29112 11980 29124
rect 12032 29112 12038 29164
rect 15654 29152 15660 29164
rect 15615 29124 15660 29152
rect 15654 29112 15660 29124
rect 15712 29112 15718 29164
rect 17926 29152 17954 29192
rect 18506 29180 18512 29192
rect 18564 29220 18570 29232
rect 19242 29220 19248 29232
rect 18564 29192 19248 29220
rect 18564 29180 18570 29192
rect 19242 29180 19248 29192
rect 19300 29180 19306 29232
rect 19426 29180 19432 29232
rect 19484 29220 19490 29232
rect 19996 29229 20024 29260
rect 23474 29248 23480 29260
rect 23532 29248 23538 29300
rect 24578 29288 24584 29300
rect 23584 29260 24584 29288
rect 19889 29223 19947 29229
rect 19889 29220 19901 29223
rect 19484 29192 19901 29220
rect 19484 29180 19490 29192
rect 19889 29189 19901 29192
rect 19935 29189 19947 29223
rect 19889 29183 19947 29189
rect 19981 29223 20039 29229
rect 19981 29189 19993 29223
rect 20027 29189 20039 29223
rect 22554 29220 22560 29232
rect 19981 29183 20039 29189
rect 22066 29192 22560 29220
rect 15764 29124 17954 29152
rect 18049 29155 18107 29161
rect 15764 29084 15792 29124
rect 18049 29121 18061 29155
rect 18095 29152 18107 29155
rect 18138 29152 18144 29164
rect 18095 29124 18144 29152
rect 18095 29121 18107 29124
rect 18049 29115 18107 29121
rect 18138 29112 18144 29124
rect 18196 29152 18202 29164
rect 18601 29155 18659 29161
rect 18601 29152 18613 29155
rect 18196 29124 18613 29152
rect 18196 29112 18202 29124
rect 18601 29121 18613 29124
rect 18647 29152 18659 29155
rect 18782 29152 18788 29164
rect 18647 29124 18788 29152
rect 18647 29121 18659 29124
rect 18601 29115 18659 29121
rect 18782 29112 18788 29124
rect 18840 29112 18846 29164
rect 19334 29112 19340 29164
rect 19392 29152 19398 29164
rect 19705 29155 19763 29161
rect 19705 29152 19717 29155
rect 19392 29124 19717 29152
rect 19392 29112 19398 29124
rect 19705 29121 19717 29124
rect 19751 29121 19763 29155
rect 19705 29115 19763 29121
rect 20073 29155 20131 29161
rect 20073 29121 20085 29155
rect 20119 29121 20131 29155
rect 20073 29115 20131 29121
rect 11624 29056 15792 29084
rect 11517 29047 11575 29053
rect 17402 29044 17408 29096
rect 17460 29084 17466 29096
rect 17460 29056 19288 29084
rect 17460 29044 17466 29056
rect 9214 29016 9220 29028
rect 7576 28988 9220 29016
rect 9214 28976 9220 28988
rect 9272 28976 9278 29028
rect 9398 28976 9404 29028
rect 9456 28988 9490 29028
rect 9456 28976 9462 28988
rect 17310 28976 17316 29028
rect 17368 29016 17374 29028
rect 18046 29016 18052 29028
rect 17368 28988 18052 29016
rect 17368 28976 17374 28988
rect 18046 28976 18052 28988
rect 18104 28976 18110 29028
rect 18785 29019 18843 29025
rect 18785 28985 18797 29019
rect 18831 29016 18843 29019
rect 18874 29016 18880 29028
rect 18831 28988 18880 29016
rect 18831 28985 18843 28988
rect 18785 28979 18843 28985
rect 18874 28976 18880 28988
rect 18932 28976 18938 29028
rect 19260 29016 19288 29056
rect 19978 29044 19984 29096
rect 20036 29084 20042 29096
rect 20088 29084 20116 29115
rect 21450 29112 21456 29164
rect 21508 29152 21514 29164
rect 22066 29152 22094 29192
rect 22554 29180 22560 29192
rect 22612 29180 22618 29232
rect 23290 29180 23296 29232
rect 23348 29220 23354 29232
rect 23584 29229 23612 29260
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 25409 29291 25467 29297
rect 25409 29257 25421 29291
rect 25455 29288 25467 29291
rect 25498 29288 25504 29300
rect 25455 29260 25504 29288
rect 25455 29257 25467 29260
rect 25409 29251 25467 29257
rect 25498 29248 25504 29260
rect 25556 29248 25562 29300
rect 30377 29291 30435 29297
rect 30377 29257 30389 29291
rect 30423 29288 30435 29291
rect 30742 29288 30748 29300
rect 30423 29260 30748 29288
rect 30423 29257 30435 29260
rect 30377 29251 30435 29257
rect 30742 29248 30748 29260
rect 30800 29248 30806 29300
rect 30834 29248 30840 29300
rect 30892 29288 30898 29300
rect 34606 29288 34612 29300
rect 30892 29260 30937 29288
rect 31726 29260 34612 29288
rect 30892 29248 30898 29260
rect 23569 29223 23627 29229
rect 23569 29220 23581 29223
rect 23348 29192 23581 29220
rect 23348 29180 23354 29192
rect 23569 29189 23581 29192
rect 23615 29189 23627 29223
rect 23569 29183 23627 29189
rect 23753 29223 23811 29229
rect 23753 29189 23765 29223
rect 23799 29220 23811 29223
rect 24670 29220 24676 29232
rect 23799 29192 24419 29220
rect 23799 29189 23811 29192
rect 23753 29183 23811 29189
rect 24391 29164 24419 29192
rect 24596 29192 24676 29220
rect 21508 29124 22094 29152
rect 23385 29155 23443 29161
rect 21508 29112 21514 29124
rect 23385 29121 23397 29155
rect 23431 29152 23443 29155
rect 23658 29152 23664 29164
rect 23431 29124 23664 29152
rect 23431 29121 23443 29124
rect 23385 29115 23443 29121
rect 23400 29084 23428 29115
rect 23658 29112 23664 29124
rect 23716 29112 23722 29164
rect 24210 29152 24216 29164
rect 24171 29124 24216 29152
rect 24210 29112 24216 29124
rect 24268 29112 24274 29164
rect 24376 29158 24434 29164
rect 24376 29124 24388 29158
rect 24422 29124 24434 29158
rect 24376 29118 24434 29124
rect 24492 29158 24550 29164
rect 24596 29161 24624 29192
rect 24670 29180 24676 29192
rect 24728 29220 24734 29232
rect 30006 29220 30012 29232
rect 24728 29192 30012 29220
rect 24728 29180 24734 29192
rect 30006 29180 30012 29192
rect 30064 29180 30070 29232
rect 30558 29180 30564 29232
rect 30616 29220 30622 29232
rect 30616 29192 31064 29220
rect 30616 29180 30622 29192
rect 24492 29124 24504 29158
rect 24538 29124 24550 29158
rect 24492 29118 24550 29124
rect 24581 29155 24639 29161
rect 24581 29121 24593 29155
rect 24627 29121 24639 29155
rect 20036 29056 20116 29084
rect 20180 29056 23428 29084
rect 20036 29044 20042 29056
rect 20180 29016 20208 29056
rect 23750 29044 23756 29096
rect 23808 29084 23814 29096
rect 24504 29084 24532 29118
rect 24581 29115 24639 29121
rect 24946 29112 24952 29164
rect 25004 29152 25010 29164
rect 25593 29155 25651 29161
rect 25593 29152 25605 29155
rect 25004 29124 25605 29152
rect 25004 29112 25010 29124
rect 25593 29121 25605 29124
rect 25639 29152 25651 29155
rect 26142 29152 26148 29164
rect 25639 29124 26148 29152
rect 25639 29121 25651 29124
rect 25593 29115 25651 29121
rect 26142 29112 26148 29124
rect 26200 29112 26206 29164
rect 30098 29112 30104 29164
rect 30156 29152 30162 29164
rect 30193 29155 30251 29161
rect 30193 29152 30205 29155
rect 30156 29124 30205 29152
rect 30156 29112 30162 29124
rect 30193 29121 30205 29124
rect 30239 29121 30251 29155
rect 30834 29152 30840 29164
rect 30795 29124 30840 29152
rect 30193 29115 30251 29121
rect 30834 29112 30840 29124
rect 30892 29112 30898 29164
rect 31036 29161 31064 29192
rect 31021 29155 31079 29161
rect 31021 29121 31033 29155
rect 31067 29121 31079 29155
rect 31021 29115 31079 29121
rect 29457 29087 29515 29093
rect 29457 29084 29469 29087
rect 23808 29056 24532 29084
rect 24642 29056 29469 29084
rect 23808 29044 23814 29056
rect 19260 28988 20208 29016
rect 20257 29019 20315 29025
rect 20257 28985 20269 29019
rect 20303 29016 20315 29019
rect 20346 29016 20352 29028
rect 20303 28988 20352 29016
rect 20303 28985 20315 28988
rect 20257 28979 20315 28985
rect 20346 28976 20352 28988
rect 20404 28976 20410 29028
rect 22741 29019 22799 29025
rect 22741 28985 22753 29019
rect 22787 29016 22799 29019
rect 22830 29016 22836 29028
rect 22787 28988 22836 29016
rect 22787 28985 22799 28988
rect 22741 28979 22799 28985
rect 22830 28976 22836 28988
rect 22888 29016 22894 29028
rect 23198 29016 23204 29028
rect 22888 28988 23204 29016
rect 22888 28976 22894 28988
rect 23198 28976 23204 28988
rect 23256 28976 23262 29028
rect 24118 28976 24124 29028
rect 24176 29016 24182 29028
rect 24642 29016 24670 29056
rect 29457 29053 29469 29056
rect 29503 29084 29515 29087
rect 30009 29087 30067 29093
rect 30009 29084 30021 29087
rect 29503 29056 30021 29084
rect 29503 29053 29515 29056
rect 29457 29047 29515 29053
rect 30009 29053 30021 29056
rect 30055 29084 30067 29087
rect 30650 29084 30656 29096
rect 30055 29056 30656 29084
rect 30055 29053 30067 29056
rect 30009 29047 30067 29053
rect 30650 29044 30656 29056
rect 30708 29044 30714 29096
rect 30742 29044 30748 29096
rect 30800 29084 30806 29096
rect 31726 29084 31754 29260
rect 34606 29248 34612 29260
rect 34664 29248 34670 29300
rect 36262 29248 36268 29300
rect 36320 29288 36326 29300
rect 38105 29291 38163 29297
rect 38105 29288 38117 29291
rect 36320 29260 38117 29288
rect 36320 29248 36326 29260
rect 38105 29257 38117 29260
rect 38151 29257 38163 29291
rect 38105 29251 38163 29257
rect 35253 29223 35311 29229
rect 35253 29189 35265 29223
rect 35299 29220 35311 29223
rect 35526 29220 35532 29232
rect 35299 29192 35532 29220
rect 35299 29189 35311 29192
rect 35253 29183 35311 29189
rect 35526 29180 35532 29192
rect 35584 29180 35590 29232
rect 35621 29223 35679 29229
rect 35621 29189 35633 29223
rect 35667 29220 35679 29223
rect 35667 29192 36308 29220
rect 35667 29189 35679 29192
rect 35621 29183 35679 29189
rect 33410 29152 33416 29164
rect 33371 29124 33416 29152
rect 33410 29112 33416 29124
rect 33468 29112 33474 29164
rect 35434 29152 35440 29164
rect 35395 29124 35440 29152
rect 35434 29112 35440 29124
rect 35492 29112 35498 29164
rect 36078 29152 36084 29164
rect 36039 29124 36084 29152
rect 36078 29112 36084 29124
rect 36136 29112 36142 29164
rect 36280 29161 36308 29192
rect 37458 29180 37464 29232
rect 37516 29220 37522 29232
rect 39218 29223 39276 29229
rect 39218 29220 39230 29223
rect 37516 29192 39230 29220
rect 37516 29180 37522 29192
rect 39218 29189 39230 29192
rect 39264 29189 39276 29223
rect 39218 29183 39276 29189
rect 36538 29161 36544 29164
rect 36265 29155 36323 29161
rect 36265 29121 36277 29155
rect 36311 29121 36323 29155
rect 36265 29115 36323 29121
rect 36357 29155 36415 29161
rect 36357 29121 36369 29155
rect 36403 29121 36415 29155
rect 36357 29115 36415 29121
rect 36495 29155 36544 29161
rect 36495 29121 36507 29155
rect 36541 29121 36544 29155
rect 36495 29115 36544 29121
rect 30800 29056 31754 29084
rect 30800 29044 30806 29056
rect 33594 29044 33600 29096
rect 33652 29084 33658 29096
rect 33689 29087 33747 29093
rect 33689 29084 33701 29087
rect 33652 29056 33701 29084
rect 33652 29044 33658 29056
rect 33689 29053 33701 29056
rect 33735 29053 33747 29087
rect 33689 29047 33747 29053
rect 34238 29044 34244 29096
rect 34296 29084 34302 29096
rect 36096 29084 36124 29112
rect 34296 29056 36124 29084
rect 36372 29084 36400 29115
rect 36538 29112 36544 29115
rect 36596 29112 36602 29164
rect 39482 29084 39488 29096
rect 36372 29056 36492 29084
rect 39443 29056 39488 29084
rect 34296 29044 34302 29056
rect 36464 29028 36492 29056
rect 39482 29044 39488 29056
rect 39540 29044 39546 29096
rect 24176 28988 24670 29016
rect 24857 29019 24915 29025
rect 24176 28976 24182 28988
rect 24857 28985 24869 29019
rect 24903 29016 24915 29019
rect 25590 29016 25596 29028
rect 24903 28988 25596 29016
rect 24903 28985 24915 28988
rect 24857 28979 24915 28985
rect 25590 28976 25596 28988
rect 25648 28976 25654 29028
rect 26142 29016 26148 29028
rect 26103 28988 26148 29016
rect 26142 28976 26148 28988
rect 26200 28976 26206 29028
rect 36446 28976 36452 29028
rect 36504 28976 36510 29028
rect 36725 29019 36783 29025
rect 36725 28985 36737 29019
rect 36771 29016 36783 29019
rect 38378 29016 38384 29028
rect 36771 28988 38384 29016
rect 36771 28985 36783 28988
rect 36725 28979 36783 28985
rect 38378 28976 38384 28988
rect 38436 28976 38442 29028
rect 3973 28951 4031 28957
rect 3973 28948 3985 28951
rect 2976 28920 3985 28948
rect 3973 28917 3985 28920
rect 4019 28948 4031 28951
rect 7374 28948 7380 28960
rect 4019 28920 7380 28948
rect 4019 28917 4031 28920
rect 3973 28911 4031 28917
rect 7374 28908 7380 28920
rect 7432 28908 7438 28960
rect 9030 28948 9036 28960
rect 8991 28920 9036 28948
rect 9030 28908 9036 28920
rect 9088 28908 9094 28960
rect 9306 28908 9312 28960
rect 9364 28948 9370 28960
rect 10778 28948 10784 28960
rect 9364 28920 10784 28948
rect 9364 28908 9370 28920
rect 10778 28908 10784 28920
rect 10836 28908 10842 28960
rect 13630 28908 13636 28960
rect 13688 28948 13694 28960
rect 13817 28951 13875 28957
rect 13817 28948 13829 28951
rect 13688 28920 13829 28948
rect 13688 28908 13694 28920
rect 13817 28917 13829 28920
rect 13863 28917 13875 28951
rect 13817 28911 13875 28917
rect 15562 28908 15568 28960
rect 15620 28948 15626 28960
rect 15841 28951 15899 28957
rect 15841 28948 15853 28951
rect 15620 28920 15853 28948
rect 15620 28908 15626 28920
rect 15841 28917 15853 28920
rect 15887 28917 15899 28951
rect 15841 28911 15899 28917
rect 16945 28951 17003 28957
rect 16945 28917 16957 28951
rect 16991 28948 17003 28951
rect 17126 28948 17132 28960
rect 16991 28920 17132 28948
rect 16991 28917 17003 28920
rect 16945 28911 17003 28917
rect 17126 28908 17132 28920
rect 17184 28908 17190 28960
rect 20530 28908 20536 28960
rect 20588 28948 20594 28960
rect 25866 28948 25872 28960
rect 20588 28920 25872 28948
rect 20588 28908 20594 28920
rect 25866 28908 25872 28920
rect 25924 28908 25930 28960
rect 30834 28908 30840 28960
rect 30892 28948 30898 28960
rect 31386 28948 31392 28960
rect 30892 28920 31392 28948
rect 30892 28908 30898 28920
rect 31386 28908 31392 28920
rect 31444 28948 31450 28960
rect 31481 28951 31539 28957
rect 31481 28948 31493 28951
rect 31444 28920 31493 28948
rect 31444 28908 31450 28920
rect 31481 28917 31493 28920
rect 31527 28917 31539 28951
rect 31481 28911 31539 28917
rect 36354 28908 36360 28960
rect 36412 28948 36418 28960
rect 36538 28948 36544 28960
rect 36412 28920 36544 28948
rect 36412 28908 36418 28920
rect 36538 28908 36544 28920
rect 36596 28948 36602 28960
rect 37277 28951 37335 28957
rect 37277 28948 37289 28951
rect 36596 28920 37289 28948
rect 36596 28908 36602 28920
rect 37277 28917 37289 28920
rect 37323 28917 37335 28951
rect 37277 28911 37335 28917
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 2593 28747 2651 28753
rect 2593 28713 2605 28747
rect 2639 28744 2651 28747
rect 2682 28744 2688 28756
rect 2639 28716 2688 28744
rect 2639 28713 2651 28716
rect 2593 28707 2651 28713
rect 2682 28704 2688 28716
rect 2740 28704 2746 28756
rect 3786 28744 3792 28756
rect 3747 28716 3792 28744
rect 3786 28704 3792 28716
rect 3844 28704 3850 28756
rect 7558 28744 7564 28756
rect 7519 28716 7564 28744
rect 7558 28704 7564 28716
rect 7616 28704 7622 28756
rect 9122 28704 9128 28756
rect 9180 28744 9186 28756
rect 10321 28747 10379 28753
rect 10321 28744 10333 28747
rect 9180 28716 10333 28744
rect 9180 28704 9186 28716
rect 10321 28713 10333 28716
rect 10367 28713 10379 28747
rect 10778 28744 10784 28756
rect 10739 28716 10784 28744
rect 10321 28707 10379 28713
rect 10336 28676 10364 28707
rect 10778 28704 10784 28716
rect 10836 28704 10842 28756
rect 13078 28704 13084 28756
rect 13136 28744 13142 28756
rect 15197 28747 15255 28753
rect 13136 28716 14136 28744
rect 13136 28704 13142 28716
rect 12526 28676 12532 28688
rect 10336 28648 12532 28676
rect 12526 28636 12532 28648
rect 12584 28636 12590 28688
rect 12986 28636 12992 28688
rect 13044 28676 13050 28688
rect 13044 28648 13308 28676
rect 13044 28636 13050 28648
rect 2777 28543 2835 28549
rect 2777 28509 2789 28543
rect 2823 28540 2835 28543
rect 3694 28540 3700 28552
rect 2823 28512 3700 28540
rect 2823 28509 2835 28512
rect 2777 28503 2835 28509
rect 3694 28500 3700 28512
rect 3752 28500 3758 28552
rect 3970 28540 3976 28552
rect 3883 28512 3976 28540
rect 3970 28500 3976 28512
rect 4028 28540 4034 28552
rect 4709 28543 4767 28549
rect 4709 28540 4721 28543
rect 4028 28512 4721 28540
rect 4028 28500 4034 28512
rect 4709 28509 4721 28512
rect 4755 28509 4767 28543
rect 4982 28540 4988 28552
rect 4943 28512 4988 28540
rect 4709 28503 4767 28509
rect 4982 28500 4988 28512
rect 5040 28500 5046 28552
rect 5077 28543 5135 28549
rect 5077 28509 5089 28543
rect 5123 28540 5135 28543
rect 5166 28540 5172 28552
rect 5123 28512 5172 28540
rect 5123 28509 5135 28512
rect 5077 28503 5135 28509
rect 5166 28500 5172 28512
rect 5224 28500 5230 28552
rect 8941 28543 8999 28549
rect 7116 28512 7788 28540
rect 2961 28475 3019 28481
rect 2961 28441 2973 28475
rect 3007 28472 3019 28475
rect 3602 28472 3608 28484
rect 3007 28444 3608 28472
rect 3007 28441 3019 28444
rect 2961 28435 3019 28441
rect 3602 28432 3608 28444
rect 3660 28472 3666 28484
rect 4157 28475 4215 28481
rect 4157 28472 4169 28475
rect 3660 28444 4169 28472
rect 3660 28432 3666 28444
rect 4157 28441 4169 28444
rect 4203 28441 4215 28475
rect 4157 28435 4215 28441
rect 4893 28475 4951 28481
rect 4893 28441 4905 28475
rect 4939 28472 4951 28475
rect 7116 28472 7144 28512
rect 7650 28472 7656 28484
rect 4939 28444 7144 28472
rect 7611 28444 7656 28472
rect 4939 28441 4951 28444
rect 4893 28435 4951 28441
rect 4706 28364 4712 28416
rect 4764 28404 4770 28416
rect 4908 28404 4936 28435
rect 7650 28432 7656 28444
rect 7708 28432 7714 28484
rect 4764 28376 4936 28404
rect 5261 28407 5319 28413
rect 4764 28364 4770 28376
rect 5261 28373 5273 28407
rect 5307 28404 5319 28407
rect 6362 28404 6368 28416
rect 5307 28376 6368 28404
rect 5307 28373 5319 28376
rect 5261 28367 5319 28373
rect 6362 28364 6368 28376
rect 6420 28364 6426 28416
rect 7760 28404 7788 28512
rect 8941 28509 8953 28543
rect 8987 28540 8999 28543
rect 9766 28540 9772 28552
rect 8987 28512 9772 28540
rect 8987 28509 8999 28512
rect 8941 28503 8999 28509
rect 9766 28500 9772 28512
rect 9824 28540 9830 28552
rect 10502 28540 10508 28552
rect 9824 28512 10508 28540
rect 9824 28500 9830 28512
rect 10502 28500 10508 28512
rect 10560 28500 10566 28552
rect 13280 28549 13308 28648
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28509 13231 28543
rect 13173 28503 13231 28509
rect 13265 28543 13323 28549
rect 13265 28509 13277 28543
rect 13311 28509 13323 28543
rect 13265 28503 13323 28509
rect 9030 28432 9036 28484
rect 9088 28472 9094 28484
rect 9186 28475 9244 28481
rect 9186 28472 9198 28475
rect 9088 28444 9198 28472
rect 9088 28432 9094 28444
rect 9186 28441 9198 28444
rect 9232 28441 9244 28475
rect 9186 28435 9244 28441
rect 9490 28404 9496 28416
rect 7760 28376 9496 28404
rect 9490 28364 9496 28376
rect 9548 28364 9554 28416
rect 11882 28364 11888 28416
rect 11940 28404 11946 28416
rect 11977 28407 12035 28413
rect 11977 28404 11989 28407
rect 11940 28376 11989 28404
rect 11940 28364 11946 28376
rect 11977 28373 11989 28376
rect 12023 28373 12035 28407
rect 12894 28404 12900 28416
rect 12855 28376 12900 28404
rect 11977 28367 12035 28373
rect 12894 28364 12900 28376
rect 12952 28364 12958 28416
rect 13188 28404 13216 28503
rect 13354 28500 13360 28552
rect 13412 28540 13418 28552
rect 13541 28543 13599 28549
rect 13412 28512 13457 28540
rect 13412 28500 13418 28512
rect 13541 28509 13553 28543
rect 13587 28540 13599 28543
rect 13722 28540 13728 28552
rect 13587 28512 13728 28540
rect 13587 28509 13599 28512
rect 13541 28503 13599 28509
rect 13722 28500 13728 28512
rect 13780 28500 13786 28552
rect 14108 28549 14136 28716
rect 15197 28713 15209 28747
rect 15243 28744 15255 28747
rect 15654 28744 15660 28756
rect 15243 28716 15660 28744
rect 15243 28713 15255 28716
rect 15197 28707 15255 28713
rect 15212 28608 15240 28707
rect 15654 28704 15660 28716
rect 15712 28704 15718 28756
rect 17218 28704 17224 28756
rect 17276 28744 17282 28756
rect 24946 28744 24952 28756
rect 17276 28716 24952 28744
rect 17276 28704 17282 28716
rect 24946 28704 24952 28716
rect 25004 28704 25010 28756
rect 25041 28747 25099 28753
rect 25041 28713 25053 28747
rect 25087 28744 25099 28747
rect 25774 28744 25780 28756
rect 25087 28716 25780 28744
rect 25087 28713 25099 28716
rect 25041 28707 25099 28713
rect 25774 28704 25780 28716
rect 25832 28744 25838 28756
rect 34330 28744 34336 28756
rect 25832 28716 34336 28744
rect 25832 28704 25838 28716
rect 34330 28704 34336 28716
rect 34388 28744 34394 28756
rect 36354 28744 36360 28756
rect 34388 28716 36360 28744
rect 34388 28704 34394 28716
rect 36354 28704 36360 28716
rect 36412 28704 36418 28756
rect 36449 28747 36507 28753
rect 36449 28713 36461 28747
rect 36495 28744 36507 28747
rect 36998 28744 37004 28756
rect 36495 28716 37004 28744
rect 36495 28713 36507 28716
rect 36449 28707 36507 28713
rect 36998 28704 37004 28716
rect 37056 28704 37062 28756
rect 19426 28636 19432 28688
rect 19484 28676 19490 28688
rect 21450 28676 21456 28688
rect 19484 28648 21456 28676
rect 19484 28636 19490 28648
rect 21450 28636 21456 28648
rect 21508 28636 21514 28688
rect 14476 28580 15240 28608
rect 16577 28611 16635 28617
rect 14093 28543 14151 28549
rect 14093 28509 14105 28543
rect 14139 28509 14151 28543
rect 14093 28503 14151 28509
rect 14182 28500 14188 28552
rect 14240 28540 14246 28552
rect 14476 28549 14504 28580
rect 16577 28577 16589 28611
rect 16623 28608 16635 28611
rect 17954 28608 17960 28620
rect 16623 28580 17960 28608
rect 16623 28577 16635 28580
rect 16577 28571 16635 28577
rect 17954 28568 17960 28580
rect 18012 28568 18018 28620
rect 20070 28568 20076 28620
rect 20128 28608 20134 28620
rect 20128 28580 21680 28608
rect 20128 28568 20134 28580
rect 14461 28543 14519 28549
rect 14240 28512 14285 28540
rect 14240 28500 14246 28512
rect 14461 28509 14473 28543
rect 14507 28509 14519 28543
rect 14461 28503 14519 28509
rect 14550 28500 14556 28552
rect 14608 28549 14614 28552
rect 14608 28540 14616 28549
rect 15194 28540 15200 28552
rect 14608 28512 15200 28540
rect 14608 28503 14616 28512
rect 14608 28500 14614 28503
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 17037 28543 17095 28549
rect 17037 28509 17049 28543
rect 17083 28540 17095 28543
rect 17126 28540 17132 28552
rect 17083 28512 17132 28540
rect 17083 28509 17095 28512
rect 17037 28503 17095 28509
rect 17126 28500 17132 28512
rect 17184 28500 17190 28552
rect 19978 28500 19984 28552
rect 20036 28540 20042 28552
rect 21652 28549 21680 28580
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 22738 28608 22744 28620
rect 22152 28580 22744 28608
rect 22152 28568 22158 28580
rect 22738 28568 22744 28580
rect 22796 28568 22802 28620
rect 30469 28611 30527 28617
rect 30469 28577 30481 28611
rect 30515 28608 30527 28611
rect 30558 28608 30564 28620
rect 30515 28580 30564 28608
rect 30515 28577 30527 28580
rect 30469 28571 30527 28577
rect 30558 28568 30564 28580
rect 30616 28568 30622 28620
rect 33502 28608 33508 28620
rect 33463 28580 33508 28608
rect 33502 28568 33508 28580
rect 33560 28568 33566 28620
rect 34992 28580 36308 28608
rect 21269 28543 21327 28549
rect 21269 28540 21281 28543
rect 20036 28512 21281 28540
rect 20036 28500 20042 28512
rect 14369 28475 14427 28481
rect 14369 28441 14381 28475
rect 14415 28472 14427 28475
rect 14826 28472 14832 28484
rect 14415 28444 14832 28472
rect 14415 28441 14427 28444
rect 14369 28435 14427 28441
rect 14826 28432 14832 28444
rect 14884 28432 14890 28484
rect 16022 28432 16028 28484
rect 16080 28472 16086 28484
rect 16310 28475 16368 28481
rect 16310 28472 16322 28475
rect 16080 28444 16322 28472
rect 16080 28432 16086 28444
rect 16310 28441 16322 28444
rect 16356 28441 16368 28475
rect 16310 28435 16368 28441
rect 13630 28404 13636 28416
rect 13188 28376 13636 28404
rect 13630 28364 13636 28376
rect 13688 28364 13694 28416
rect 14737 28407 14795 28413
rect 14737 28373 14749 28407
rect 14783 28404 14795 28407
rect 15194 28404 15200 28416
rect 14783 28376 15200 28404
rect 14783 28373 14795 28376
rect 14737 28367 14795 28373
rect 15194 28364 15200 28376
rect 15252 28364 15258 28416
rect 17221 28407 17279 28413
rect 17221 28373 17233 28407
rect 17267 28404 17279 28407
rect 17310 28404 17316 28416
rect 17267 28376 17316 28404
rect 17267 28373 17279 28376
rect 17221 28367 17279 28373
rect 17310 28364 17316 28376
rect 17368 28404 17374 28416
rect 17494 28404 17500 28416
rect 17368 28376 17500 28404
rect 17368 28364 17374 28376
rect 17494 28364 17500 28376
rect 17552 28364 17558 28416
rect 21082 28404 21088 28416
rect 21043 28376 21088 28404
rect 21082 28364 21088 28376
rect 21140 28364 21146 28416
rect 21192 28404 21220 28512
rect 21269 28509 21281 28512
rect 21315 28509 21327 28543
rect 21269 28503 21327 28509
rect 21361 28543 21419 28549
rect 21361 28509 21373 28543
rect 21407 28540 21419 28543
rect 21637 28543 21695 28549
rect 21407 28512 21588 28540
rect 21407 28509 21419 28512
rect 21361 28503 21419 28509
rect 21450 28472 21456 28484
rect 21411 28444 21456 28472
rect 21450 28432 21456 28444
rect 21508 28432 21514 28484
rect 21560 28472 21588 28512
rect 21637 28509 21649 28543
rect 21683 28509 21695 28543
rect 23290 28540 23296 28552
rect 21637 28503 21695 28509
rect 22066 28512 23296 28540
rect 22066 28472 22094 28512
rect 23290 28500 23296 28512
rect 23348 28500 23354 28552
rect 24118 28500 24124 28552
rect 24176 28540 24182 28552
rect 28997 28543 29055 28549
rect 28997 28540 29009 28543
rect 24176 28512 29009 28540
rect 24176 28500 24182 28512
rect 28997 28509 29009 28512
rect 29043 28540 29055 28543
rect 30742 28540 30748 28552
rect 29043 28512 30748 28540
rect 29043 28509 29055 28512
rect 28997 28503 29055 28509
rect 30742 28500 30748 28512
rect 30800 28500 30806 28552
rect 31205 28543 31263 28549
rect 31205 28509 31217 28543
rect 31251 28509 31263 28543
rect 31386 28540 31392 28552
rect 31347 28512 31392 28540
rect 31205 28503 31263 28509
rect 21560 28444 22094 28472
rect 22649 28475 22707 28481
rect 22649 28441 22661 28475
rect 22695 28441 22707 28475
rect 25130 28472 25136 28484
rect 25091 28444 25136 28472
rect 22649 28435 22707 28441
rect 22186 28404 22192 28416
rect 21192 28376 22192 28404
rect 22186 28364 22192 28376
rect 22244 28404 22250 28416
rect 22664 28404 22692 28435
rect 25130 28432 25136 28444
rect 25188 28432 25194 28484
rect 30098 28432 30104 28484
rect 30156 28472 30162 28484
rect 31220 28472 31248 28503
rect 31386 28500 31392 28512
rect 31444 28540 31450 28552
rect 31849 28543 31907 28549
rect 31849 28540 31861 28543
rect 31444 28512 31861 28540
rect 31444 28500 31450 28512
rect 31849 28509 31861 28512
rect 31895 28509 31907 28543
rect 31849 28503 31907 28509
rect 33410 28500 33416 28552
rect 33468 28540 33474 28552
rect 34992 28549 35020 28580
rect 36280 28552 36308 28580
rect 33781 28543 33839 28549
rect 33781 28540 33793 28543
rect 33468 28512 33793 28540
rect 33468 28500 33474 28512
rect 33781 28509 33793 28512
rect 33827 28540 33839 28543
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 33827 28512 34897 28540
rect 33827 28509 33839 28512
rect 33781 28503 33839 28509
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 34977 28543 35035 28549
rect 34977 28509 34989 28543
rect 35023 28509 35035 28543
rect 34977 28503 35035 28509
rect 35253 28543 35311 28549
rect 35253 28509 35265 28543
rect 35299 28540 35311 28543
rect 35342 28540 35348 28552
rect 35299 28512 35348 28540
rect 35299 28509 35311 28512
rect 35253 28503 35311 28509
rect 35342 28500 35348 28512
rect 35400 28500 35406 28552
rect 35526 28500 35532 28552
rect 35584 28540 35590 28552
rect 36081 28543 36139 28549
rect 36081 28540 36093 28543
rect 35584 28512 36093 28540
rect 35584 28500 35590 28512
rect 36081 28509 36093 28512
rect 36127 28509 36139 28543
rect 36262 28540 36268 28552
rect 36223 28512 36268 28540
rect 36081 28503 36139 28509
rect 36262 28500 36268 28512
rect 36320 28500 36326 28552
rect 38378 28500 38384 28552
rect 38436 28549 38442 28552
rect 38436 28540 38448 28549
rect 38657 28543 38715 28549
rect 38436 28512 38481 28540
rect 38436 28503 38448 28512
rect 38657 28509 38669 28543
rect 38703 28540 38715 28543
rect 39482 28540 39488 28552
rect 38703 28512 39488 28540
rect 38703 28509 38715 28512
rect 38657 28503 38715 28509
rect 38436 28500 38442 28503
rect 39482 28500 39488 28512
rect 39540 28540 39546 28552
rect 39942 28540 39948 28552
rect 39540 28512 39948 28540
rect 39540 28500 39546 28512
rect 39942 28500 39948 28512
rect 40000 28500 40006 28552
rect 30156 28444 31248 28472
rect 30156 28432 30162 28444
rect 33594 28432 33600 28484
rect 33652 28472 33658 28484
rect 35069 28475 35127 28481
rect 35069 28472 35081 28475
rect 33652 28444 35081 28472
rect 33652 28432 33658 28444
rect 35069 28441 35081 28444
rect 35115 28441 35127 28475
rect 35069 28435 35127 28441
rect 22244 28376 22692 28404
rect 22244 28364 22250 28376
rect 22738 28364 22744 28416
rect 22796 28404 22802 28416
rect 23750 28404 23756 28416
rect 22796 28376 22841 28404
rect 23711 28376 23756 28404
rect 22796 28364 22802 28376
rect 23750 28364 23756 28376
rect 23808 28404 23814 28416
rect 24578 28404 24584 28416
rect 23808 28376 24584 28404
rect 23808 28364 23814 28376
rect 24578 28364 24584 28376
rect 24636 28364 24642 28416
rect 31389 28407 31447 28413
rect 31389 28373 31401 28407
rect 31435 28404 31447 28407
rect 31846 28404 31852 28416
rect 31435 28376 31852 28404
rect 31435 28373 31447 28376
rect 31389 28367 31447 28373
rect 31846 28364 31852 28376
rect 31904 28364 31910 28416
rect 34701 28407 34759 28413
rect 34701 28373 34713 28407
rect 34747 28404 34759 28407
rect 34790 28404 34796 28416
rect 34747 28376 34796 28404
rect 34747 28373 34759 28376
rect 34701 28367 34759 28373
rect 34790 28364 34796 28376
rect 34848 28364 34854 28416
rect 35434 28364 35440 28416
rect 35492 28404 35498 28416
rect 37277 28407 37335 28413
rect 37277 28404 37289 28407
rect 35492 28376 37289 28404
rect 35492 28364 35498 28376
rect 37277 28373 37289 28376
rect 37323 28373 37335 28407
rect 37277 28367 37335 28373
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 3970 28200 3976 28212
rect 3931 28172 3976 28200
rect 3970 28160 3976 28172
rect 4028 28160 4034 28212
rect 9398 28200 9404 28212
rect 9359 28172 9404 28200
rect 9398 28160 9404 28172
rect 9456 28160 9462 28212
rect 10042 28200 10048 28212
rect 9955 28172 10048 28200
rect 10042 28160 10048 28172
rect 10100 28200 10106 28212
rect 10778 28200 10784 28212
rect 10100 28172 10784 28200
rect 10100 28160 10106 28172
rect 10778 28160 10784 28172
rect 10836 28160 10842 28212
rect 12434 28160 12440 28212
rect 12492 28200 12498 28212
rect 13078 28200 13084 28212
rect 12492 28172 12756 28200
rect 13039 28172 13084 28200
rect 12492 28160 12498 28172
rect 6730 28132 6736 28144
rect 6691 28104 6736 28132
rect 6730 28092 6736 28104
rect 6788 28092 6794 28144
rect 9214 28092 9220 28144
rect 9272 28132 9278 28144
rect 12728 28141 12756 28172
rect 13078 28160 13084 28172
rect 13136 28160 13142 28212
rect 13354 28160 13360 28212
rect 13412 28200 13418 28212
rect 13909 28203 13967 28209
rect 13909 28200 13921 28203
rect 13412 28172 13921 28200
rect 13412 28160 13418 28172
rect 13909 28169 13921 28172
rect 13955 28169 13967 28203
rect 16022 28200 16028 28212
rect 15983 28172 16028 28200
rect 13909 28163 13967 28169
rect 16022 28160 16028 28172
rect 16080 28160 16086 28212
rect 17126 28160 17132 28212
rect 17184 28200 17190 28212
rect 17184 28172 24716 28200
rect 17184 28160 17190 28172
rect 12713 28135 12771 28141
rect 9272 28104 11744 28132
rect 9272 28092 9278 28104
rect 11716 28076 11744 28104
rect 12713 28101 12725 28135
rect 12759 28101 12771 28135
rect 12713 28095 12771 28101
rect 12805 28135 12863 28141
rect 12805 28101 12817 28135
rect 12851 28132 12863 28135
rect 13446 28132 13452 28144
rect 12851 28104 13452 28132
rect 12851 28101 12863 28104
rect 12805 28095 12863 28101
rect 13446 28092 13452 28104
rect 13504 28132 13510 28144
rect 13725 28135 13783 28141
rect 13725 28132 13737 28135
rect 13504 28104 13737 28132
rect 13504 28092 13510 28104
rect 13725 28101 13737 28104
rect 13771 28101 13783 28135
rect 13725 28095 13783 28101
rect 14642 28092 14648 28144
rect 14700 28132 14706 28144
rect 23750 28132 23756 28144
rect 14700 28104 15700 28132
rect 14700 28092 14706 28104
rect 2866 28073 2872 28076
rect 2860 28064 2872 28073
rect 2827 28036 2872 28064
rect 2860 28027 2872 28036
rect 2866 28024 2872 28027
rect 2924 28024 2930 28076
rect 6362 28064 6368 28076
rect 6323 28036 6368 28064
rect 6362 28024 6368 28036
rect 6420 28024 6426 28076
rect 6454 28024 6460 28076
rect 6512 28064 6518 28076
rect 6512 28036 6557 28064
rect 6512 28024 6518 28036
rect 6638 28024 6644 28076
rect 6696 28064 6702 28076
rect 6696 28036 6741 28064
rect 6696 28024 6702 28036
rect 6822 28024 6828 28076
rect 6880 28073 6886 28076
rect 6880 28064 6888 28073
rect 6880 28036 6925 28064
rect 6880 28027 6888 28036
rect 6880 28024 6886 28027
rect 8938 28024 8944 28076
rect 8996 28064 9002 28076
rect 9309 28067 9367 28073
rect 9309 28064 9321 28067
rect 8996 28036 9321 28064
rect 8996 28024 9002 28036
rect 9309 28033 9321 28036
rect 9355 28033 9367 28067
rect 9490 28064 9496 28076
rect 9451 28036 9496 28064
rect 9309 28027 9367 28033
rect 9490 28024 9496 28036
rect 9548 28024 9554 28076
rect 11698 28064 11704 28076
rect 11611 28036 11704 28064
rect 11698 28024 11704 28036
rect 11756 28024 11762 28076
rect 11882 28064 11888 28076
rect 11843 28036 11888 28064
rect 11882 28024 11888 28036
rect 11940 28024 11946 28076
rect 12526 28064 12532 28076
rect 12487 28036 12532 28064
rect 12526 28024 12532 28036
rect 12584 28024 12590 28076
rect 12618 28024 12624 28076
rect 12676 28064 12682 28076
rect 12897 28067 12955 28073
rect 12897 28064 12909 28067
rect 12676 28036 12909 28064
rect 12676 28024 12682 28036
rect 12897 28033 12909 28036
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 13262 28024 13268 28076
rect 13320 28064 13326 28076
rect 13541 28067 13599 28073
rect 13541 28064 13553 28067
rect 13320 28036 13553 28064
rect 13320 28024 13326 28036
rect 13541 28033 13553 28036
rect 13587 28033 13599 28067
rect 15378 28064 15384 28076
rect 15339 28036 15384 28064
rect 13541 28027 13599 28033
rect 15378 28024 15384 28036
rect 15436 28024 15442 28076
rect 15562 28064 15568 28076
rect 15523 28036 15568 28064
rect 15562 28024 15568 28036
rect 15620 28024 15626 28076
rect 15672 28073 15700 28104
rect 17696 28104 23756 28132
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28033 15715 28067
rect 15657 28027 15715 28033
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28033 15807 28067
rect 15749 28027 15807 28033
rect 17129 28067 17187 28073
rect 17129 28033 17141 28067
rect 17175 28064 17187 28067
rect 17218 28064 17224 28076
rect 17175 28036 17224 28064
rect 17175 28033 17187 28036
rect 17129 28027 17187 28033
rect 2590 27996 2596 28008
rect 2551 27968 2596 27996
rect 2590 27956 2596 27968
rect 2648 27956 2654 28008
rect 11900 27928 11928 28024
rect 13630 27956 13636 28008
rect 13688 27996 13694 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 13688 27968 14933 27996
rect 13688 27956 13694 27968
rect 14921 27965 14933 27968
rect 14967 27996 14979 27999
rect 15764 27996 15792 28027
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 17696 28064 17724 28104
rect 23750 28092 23756 28104
rect 23808 28092 23814 28144
rect 17328 28036 17724 28064
rect 18049 28067 18107 28073
rect 17328 27996 17356 28036
rect 18049 28033 18061 28067
rect 18095 28064 18107 28067
rect 19426 28064 19432 28076
rect 18095 28036 19432 28064
rect 18095 28033 18107 28036
rect 18049 28027 18107 28033
rect 19426 28024 19432 28036
rect 19484 28024 19490 28076
rect 19978 28064 19984 28076
rect 19939 28036 19984 28064
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 14967 27968 17356 27996
rect 14967 27965 14979 27968
rect 14921 27959 14979 27965
rect 17678 27956 17684 28008
rect 17736 27996 17742 28008
rect 17773 27999 17831 28005
rect 17773 27996 17785 27999
rect 17736 27968 17785 27996
rect 17736 27956 17742 27968
rect 17773 27965 17785 27968
rect 17819 27965 17831 27999
rect 17773 27959 17831 27965
rect 19334 27956 19340 28008
rect 19392 27996 19398 28008
rect 19705 27999 19763 28005
rect 19705 27996 19717 27999
rect 19392 27968 19717 27996
rect 19392 27956 19398 27968
rect 19705 27965 19717 27968
rect 19751 27965 19763 27999
rect 19705 27959 19763 27965
rect 17954 27928 17960 27940
rect 11900 27900 17960 27928
rect 17954 27888 17960 27900
rect 18012 27888 18018 27940
rect 21174 27928 21180 27940
rect 18984 27900 21180 27928
rect 7006 27860 7012 27872
rect 6967 27832 7012 27860
rect 7006 27820 7012 27832
rect 7064 27820 7070 27872
rect 8849 27863 8907 27869
rect 8849 27829 8861 27863
rect 8895 27860 8907 27863
rect 8938 27860 8944 27872
rect 8895 27832 8944 27860
rect 8895 27829 8907 27832
rect 8849 27823 8907 27829
rect 8938 27820 8944 27832
rect 8996 27820 9002 27872
rect 10597 27863 10655 27869
rect 10597 27829 10609 27863
rect 10643 27860 10655 27863
rect 11054 27860 11060 27872
rect 10643 27832 11060 27860
rect 10643 27829 10655 27832
rect 10597 27823 10655 27829
rect 11054 27820 11060 27832
rect 11112 27820 11118 27872
rect 11517 27863 11575 27869
rect 11517 27829 11529 27863
rect 11563 27860 11575 27863
rect 13262 27860 13268 27872
rect 11563 27832 13268 27860
rect 11563 27829 11575 27832
rect 11517 27823 11575 27829
rect 13262 27820 13268 27832
rect 13320 27820 13326 27872
rect 17221 27863 17279 27869
rect 17221 27829 17233 27863
rect 17267 27860 17279 27863
rect 18984 27860 19012 27900
rect 21174 27888 21180 27900
rect 21232 27928 21238 27940
rect 21634 27928 21640 27940
rect 21232 27900 21640 27928
rect 21232 27888 21238 27900
rect 21634 27888 21640 27900
rect 21692 27888 21698 27940
rect 24688 27937 24716 28172
rect 34241 28135 34299 28141
rect 34241 28101 34253 28135
rect 34287 28132 34299 28135
rect 35434 28132 35440 28144
rect 34287 28104 35440 28132
rect 34287 28101 34299 28104
rect 34241 28095 34299 28101
rect 35434 28092 35440 28104
rect 35492 28092 35498 28144
rect 26418 28064 26424 28076
rect 26331 28036 26424 28064
rect 26418 28024 26424 28036
rect 26476 28064 26482 28076
rect 27249 28067 27307 28073
rect 27249 28064 27261 28067
rect 26476 28036 27261 28064
rect 26476 28024 26482 28036
rect 27249 28033 27261 28036
rect 27295 28064 27307 28067
rect 29362 28064 29368 28076
rect 27295 28036 29368 28064
rect 27295 28033 27307 28036
rect 27249 28027 27307 28033
rect 29362 28024 29368 28036
rect 29420 28024 29426 28076
rect 30009 28067 30067 28073
rect 30009 28033 30021 28067
rect 30055 28064 30067 28067
rect 30098 28064 30104 28076
rect 30055 28036 30104 28064
rect 30055 28033 30067 28036
rect 30009 28027 30067 28033
rect 30098 28024 30104 28036
rect 30156 28024 30162 28076
rect 30742 28024 30748 28076
rect 30800 28064 30806 28076
rect 31573 28067 31631 28073
rect 31573 28064 31585 28067
rect 30800 28036 31585 28064
rect 30800 28024 30806 28036
rect 31573 28033 31585 28036
rect 31619 28064 31631 28067
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 31619 28036 32137 28064
rect 31619 28033 31631 28036
rect 31573 28027 31631 28033
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 33410 28024 33416 28076
rect 33468 28064 33474 28076
rect 34149 28067 34207 28073
rect 34149 28064 34161 28067
rect 33468 28036 34161 28064
rect 33468 28024 33474 28036
rect 34149 28033 34161 28036
rect 34195 28033 34207 28067
rect 34149 28027 34207 28033
rect 34333 28067 34391 28073
rect 34333 28033 34345 28067
rect 34379 28033 34391 28067
rect 34514 28064 34520 28076
rect 34475 28036 34520 28064
rect 34333 28027 34391 28033
rect 30285 27999 30343 28005
rect 30285 27996 30297 27999
rect 29012 27968 30297 27996
rect 24673 27931 24731 27937
rect 24673 27897 24685 27931
rect 24719 27928 24731 27931
rect 25130 27928 25136 27940
rect 24719 27900 25136 27928
rect 24719 27897 24731 27900
rect 24673 27891 24731 27897
rect 25130 27888 25136 27900
rect 25188 27928 25194 27940
rect 26602 27928 26608 27940
rect 25188 27900 26608 27928
rect 25188 27888 25194 27900
rect 26602 27888 26608 27900
rect 26660 27888 26666 27940
rect 19150 27860 19156 27872
rect 17267 27832 19012 27860
rect 19111 27832 19156 27860
rect 17267 27829 17279 27832
rect 17221 27823 17279 27829
rect 19150 27820 19156 27832
rect 19208 27820 19214 27872
rect 26694 27820 26700 27872
rect 26752 27860 26758 27872
rect 27062 27860 27068 27872
rect 26752 27832 27068 27860
rect 26752 27820 26758 27832
rect 27062 27820 27068 27832
rect 27120 27820 27126 27872
rect 28718 27820 28724 27872
rect 28776 27860 28782 27872
rect 29012 27869 29040 27968
rect 30285 27965 30297 27968
rect 30331 27996 30343 27999
rect 30466 27996 30472 28008
rect 30331 27968 30472 27996
rect 30331 27965 30343 27968
rect 30285 27959 30343 27965
rect 30466 27956 30472 27968
rect 30524 27956 30530 28008
rect 31297 27999 31355 28005
rect 31297 27965 31309 27999
rect 31343 27965 31355 27999
rect 33134 27996 33140 28008
rect 31297 27959 31355 27965
rect 31726 27968 33140 27996
rect 31312 27928 31340 27959
rect 31726 27928 31754 27968
rect 33134 27956 33140 27968
rect 33192 27996 33198 28008
rect 33594 27996 33600 28008
rect 33192 27968 33600 27996
rect 33192 27956 33198 27968
rect 33594 27956 33600 27968
rect 33652 27996 33658 28008
rect 34348 27996 34376 28027
rect 34514 28024 34520 28036
rect 34572 28024 34578 28076
rect 39689 28067 39747 28073
rect 39689 28033 39701 28067
rect 39735 28064 39747 28067
rect 39850 28064 39856 28076
rect 39735 28036 39856 28064
rect 39735 28033 39747 28036
rect 39689 28027 39747 28033
rect 39850 28024 39856 28036
rect 39908 28024 39914 28076
rect 39942 27996 39948 28008
rect 33652 27968 34376 27996
rect 39903 27968 39948 27996
rect 33652 27956 33658 27968
rect 39942 27956 39948 27968
rect 40000 27956 40006 28008
rect 58158 27928 58164 27940
rect 31312 27900 31754 27928
rect 58119 27900 58164 27928
rect 58158 27888 58164 27900
rect 58216 27888 58222 27940
rect 28997 27863 29055 27869
rect 28997 27860 29009 27863
rect 28776 27832 29009 27860
rect 28776 27820 28782 27832
rect 28997 27829 29009 27832
rect 29043 27829 29055 27863
rect 33962 27860 33968 27872
rect 33923 27832 33968 27860
rect 28997 27823 29055 27829
rect 33962 27820 33968 27832
rect 34020 27820 34026 27872
rect 38565 27863 38623 27869
rect 38565 27829 38577 27863
rect 38611 27860 38623 27863
rect 39022 27860 39028 27872
rect 38611 27832 39028 27860
rect 38611 27829 38623 27832
rect 38565 27823 38623 27829
rect 39022 27820 39028 27832
rect 39080 27820 39086 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 7650 27616 7656 27668
rect 7708 27656 7714 27668
rect 9033 27659 9091 27665
rect 9033 27656 9045 27659
rect 7708 27628 9045 27656
rect 7708 27616 7714 27628
rect 9033 27625 9045 27628
rect 9079 27656 9091 27659
rect 10410 27656 10416 27668
rect 9079 27628 10416 27656
rect 9079 27625 9091 27628
rect 9033 27619 9091 27625
rect 10410 27616 10416 27628
rect 10468 27616 10474 27668
rect 13446 27616 13452 27668
rect 13504 27656 13510 27668
rect 13541 27659 13599 27665
rect 13541 27656 13553 27659
rect 13504 27628 13553 27656
rect 13504 27616 13510 27628
rect 13541 27625 13553 27628
rect 13587 27625 13599 27659
rect 13541 27619 13599 27625
rect 16945 27659 17003 27665
rect 16945 27625 16957 27659
rect 16991 27656 17003 27659
rect 17218 27656 17224 27668
rect 16991 27628 17224 27656
rect 16991 27625 17003 27628
rect 16945 27619 17003 27625
rect 17218 27616 17224 27628
rect 17276 27616 17282 27668
rect 5442 27588 5448 27600
rect 5276 27560 5448 27588
rect 4890 27452 4896 27464
rect 4851 27424 4896 27452
rect 4890 27412 4896 27424
rect 4948 27412 4954 27464
rect 5276 27461 5304 27560
rect 5442 27548 5448 27560
rect 5500 27548 5506 27600
rect 6822 27548 6828 27600
rect 6880 27588 6886 27600
rect 9306 27588 9312 27600
rect 6880 27560 9312 27588
rect 6880 27548 6886 27560
rect 9306 27548 9312 27560
rect 9364 27548 9370 27600
rect 9674 27588 9680 27600
rect 9416 27560 9680 27588
rect 6840 27520 6868 27548
rect 6380 27492 6868 27520
rect 4986 27455 5044 27461
rect 4986 27421 4998 27455
rect 5032 27421 5044 27455
rect 4986 27415 5044 27421
rect 5261 27455 5319 27461
rect 5261 27421 5273 27455
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 5399 27455 5457 27461
rect 5399 27421 5411 27455
rect 5445 27452 5457 27455
rect 5534 27452 5540 27464
rect 5445 27424 5540 27452
rect 5445 27421 5457 27424
rect 5399 27415 5457 27421
rect 4062 27344 4068 27396
rect 4120 27384 4126 27396
rect 5000 27384 5028 27415
rect 5534 27412 5540 27424
rect 5592 27452 5598 27464
rect 6380 27452 6408 27492
rect 7098 27480 7104 27532
rect 7156 27520 7162 27532
rect 9416 27520 9444 27560
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 28994 27588 29000 27600
rect 28955 27560 29000 27588
rect 28994 27548 29000 27560
rect 29052 27548 29058 27600
rect 30466 27588 30472 27600
rect 30427 27560 30472 27588
rect 30466 27548 30472 27560
rect 30524 27588 30530 27600
rect 30524 27560 31064 27588
rect 30524 27548 30530 27560
rect 7156 27492 9444 27520
rect 9585 27523 9643 27529
rect 7156 27480 7162 27492
rect 9585 27489 9597 27523
rect 9631 27520 9643 27523
rect 9631 27492 10456 27520
rect 9631 27489 9643 27492
rect 9585 27483 9643 27489
rect 5592 27424 6408 27452
rect 5592 27412 5598 27424
rect 6454 27412 6460 27464
rect 6512 27452 6518 27464
rect 7285 27455 7343 27461
rect 7285 27452 7297 27455
rect 6512 27424 7297 27452
rect 6512 27412 6518 27424
rect 7285 27421 7297 27424
rect 7331 27421 7343 27455
rect 7285 27415 7343 27421
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27452 8447 27455
rect 8938 27452 8944 27464
rect 8435 27424 8944 27452
rect 8435 27421 8447 27424
rect 8389 27415 8447 27421
rect 8938 27412 8944 27424
rect 8996 27412 9002 27464
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27452 9183 27455
rect 9398 27452 9404 27464
rect 9171 27424 9404 27452
rect 9171 27421 9183 27424
rect 9125 27415 9183 27421
rect 4120 27356 5028 27384
rect 4120 27344 4126 27356
rect 5074 27344 5080 27396
rect 5132 27384 5138 27396
rect 5169 27387 5227 27393
rect 5169 27384 5181 27387
rect 5132 27356 5181 27384
rect 5132 27344 5138 27356
rect 5169 27353 5181 27356
rect 5215 27384 5227 27387
rect 6638 27384 6644 27396
rect 5215 27356 6644 27384
rect 5215 27353 5227 27356
rect 5169 27347 5227 27353
rect 6638 27344 6644 27356
rect 6696 27384 6702 27396
rect 7098 27384 7104 27396
rect 6696 27356 6960 27384
rect 7059 27356 7104 27384
rect 6696 27344 6702 27356
rect 5537 27319 5595 27325
rect 5537 27285 5549 27319
rect 5583 27316 5595 27319
rect 6822 27316 6828 27328
rect 5583 27288 6828 27316
rect 5583 27285 5595 27288
rect 5537 27279 5595 27285
rect 6822 27276 6828 27288
rect 6880 27276 6886 27328
rect 6932 27316 6960 27356
rect 7098 27344 7104 27356
rect 7156 27344 7162 27396
rect 9140 27384 9168 27415
rect 9398 27412 9404 27424
rect 9456 27412 9462 27464
rect 9490 27412 9496 27464
rect 9548 27452 9554 27464
rect 9861 27455 9919 27461
rect 9861 27452 9873 27455
rect 9548 27424 9873 27452
rect 9548 27412 9554 27424
rect 9861 27421 9873 27424
rect 9907 27421 9919 27455
rect 10428 27452 10456 27492
rect 10594 27480 10600 27532
rect 10652 27520 10658 27532
rect 12161 27523 12219 27529
rect 12161 27520 12173 27523
rect 10652 27492 12173 27520
rect 10652 27480 10658 27492
rect 12161 27489 12173 27492
rect 12207 27489 12219 27523
rect 12161 27483 12219 27489
rect 16022 27480 16028 27532
rect 16080 27520 16086 27532
rect 24394 27520 24400 27532
rect 16080 27492 24400 27520
rect 16080 27480 16086 27492
rect 24394 27480 24400 27492
rect 24452 27480 24458 27532
rect 31036 27529 31064 27560
rect 31021 27523 31079 27529
rect 31021 27489 31033 27523
rect 31067 27489 31079 27523
rect 34698 27520 34704 27532
rect 31021 27483 31079 27489
rect 32508 27492 33364 27520
rect 10686 27452 10692 27464
rect 10428 27424 10692 27452
rect 9861 27415 9919 27421
rect 10686 27412 10692 27424
rect 10744 27452 10750 27464
rect 10873 27455 10931 27461
rect 10873 27452 10885 27455
rect 10744 27424 10885 27452
rect 10744 27412 10750 27424
rect 10873 27421 10885 27424
rect 10919 27421 10931 27455
rect 10873 27415 10931 27421
rect 11149 27455 11207 27461
rect 11149 27421 11161 27455
rect 11195 27421 11207 27455
rect 11149 27415 11207 27421
rect 12428 27455 12486 27461
rect 12428 27421 12440 27455
rect 12474 27452 12486 27455
rect 12894 27452 12900 27464
rect 12474 27424 12900 27452
rect 12474 27421 12486 27424
rect 12428 27415 12486 27421
rect 7208 27356 9168 27384
rect 7208 27316 7236 27356
rect 6932 27288 7236 27316
rect 7469 27319 7527 27325
rect 7469 27285 7481 27319
rect 7515 27316 7527 27319
rect 7650 27316 7656 27328
rect 7515 27288 7656 27316
rect 7515 27285 7527 27288
rect 7469 27279 7527 27285
rect 7650 27276 7656 27288
rect 7708 27276 7714 27328
rect 11164 27316 11192 27415
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 17954 27452 17960 27464
rect 17819 27424 17960 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 17954 27412 17960 27424
rect 18012 27452 18018 27464
rect 18233 27455 18291 27461
rect 18233 27452 18245 27455
rect 18012 27424 18245 27452
rect 18012 27412 18018 27424
rect 18233 27421 18245 27424
rect 18279 27452 18291 27455
rect 19150 27452 19156 27464
rect 18279 27424 19156 27452
rect 18279 27421 18291 27424
rect 18233 27415 18291 27421
rect 19150 27412 19156 27424
rect 19208 27452 19214 27464
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 19208 27424 19257 27452
rect 19208 27412 19214 27424
rect 19245 27421 19257 27424
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 23385 27455 23443 27461
rect 23385 27452 23397 27455
rect 22879 27424 23397 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 23385 27421 23397 27424
rect 23431 27452 23443 27455
rect 26605 27455 26663 27461
rect 23431 27424 26556 27452
rect 23431 27421 23443 27424
rect 23385 27415 23443 27421
rect 20622 27344 20628 27396
rect 20680 27384 20686 27396
rect 21085 27387 21143 27393
rect 21085 27384 21097 27387
rect 20680 27356 21097 27384
rect 20680 27344 20686 27356
rect 21085 27353 21097 27356
rect 21131 27384 21143 27387
rect 21542 27384 21548 27396
rect 21131 27356 21548 27384
rect 21131 27353 21143 27356
rect 21085 27347 21143 27353
rect 21542 27344 21548 27356
rect 21600 27344 21606 27396
rect 25961 27387 26019 27393
rect 25961 27353 25973 27387
rect 26007 27353 26019 27387
rect 26142 27384 26148 27396
rect 26103 27356 26148 27384
rect 25961 27347 26019 27353
rect 12434 27316 12440 27328
rect 11164 27288 12440 27316
rect 12434 27276 12440 27288
rect 12492 27276 12498 27328
rect 16206 27276 16212 27328
rect 16264 27316 16270 27328
rect 16301 27319 16359 27325
rect 16301 27316 16313 27319
rect 16264 27288 16313 27316
rect 16264 27276 16270 27288
rect 16301 27285 16313 27288
rect 16347 27316 16359 27319
rect 16574 27316 16580 27328
rect 16347 27288 16580 27316
rect 16347 27285 16359 27288
rect 16301 27279 16359 27285
rect 16574 27276 16580 27288
rect 16632 27276 16638 27328
rect 18414 27316 18420 27328
rect 18375 27288 18420 27316
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 19429 27319 19487 27325
rect 19429 27285 19441 27319
rect 19475 27316 19487 27319
rect 19978 27316 19984 27328
rect 19475 27288 19984 27316
rect 19475 27285 19487 27288
rect 19429 27279 19487 27285
rect 19978 27276 19984 27288
rect 20036 27276 20042 27328
rect 24670 27316 24676 27328
rect 24631 27288 24676 27316
rect 24670 27276 24676 27288
rect 24728 27276 24734 27328
rect 24854 27276 24860 27328
rect 24912 27316 24918 27328
rect 25777 27319 25835 27325
rect 25777 27316 25789 27319
rect 24912 27288 25789 27316
rect 24912 27276 24918 27288
rect 25777 27285 25789 27288
rect 25823 27285 25835 27319
rect 25976 27316 26004 27347
rect 26142 27344 26148 27356
rect 26200 27344 26206 27396
rect 26528 27384 26556 27424
rect 26605 27421 26617 27455
rect 26651 27452 26663 27455
rect 26694 27452 26700 27464
rect 26651 27424 26700 27452
rect 26651 27421 26663 27424
rect 26605 27415 26663 27421
rect 26694 27412 26700 27424
rect 26752 27412 26758 27464
rect 28994 27452 29000 27464
rect 26804 27424 29000 27452
rect 26804 27384 26832 27424
rect 28994 27412 29000 27424
rect 29052 27412 29058 27464
rect 32508 27461 32536 27492
rect 31297 27455 31355 27461
rect 31297 27421 31309 27455
rect 31343 27452 31355 27455
rect 32493 27455 32551 27461
rect 32493 27452 32505 27455
rect 31343 27424 32505 27452
rect 31343 27421 31355 27424
rect 31297 27415 31355 27421
rect 32493 27421 32505 27424
rect 32539 27421 32551 27455
rect 32493 27415 32551 27421
rect 32585 27455 32643 27461
rect 32585 27421 32597 27455
rect 32631 27452 32643 27455
rect 32766 27452 32772 27464
rect 32631 27424 32772 27452
rect 32631 27421 32643 27424
rect 32585 27415 32643 27421
rect 32766 27412 32772 27424
rect 32824 27412 32830 27464
rect 32861 27455 32919 27461
rect 32861 27421 32873 27455
rect 32907 27452 32919 27455
rect 33226 27452 33232 27464
rect 32907 27424 33232 27452
rect 32907 27421 32919 27424
rect 32861 27415 32919 27421
rect 33226 27412 33232 27424
rect 33284 27412 33290 27464
rect 33336 27452 33364 27492
rect 33612 27492 34704 27520
rect 33410 27452 33416 27464
rect 33336 27424 33416 27452
rect 33410 27412 33416 27424
rect 33468 27461 33474 27464
rect 33612 27461 33640 27492
rect 34698 27480 34704 27492
rect 34756 27520 34762 27532
rect 34756 27492 34928 27520
rect 34756 27480 34762 27492
rect 33468 27455 33517 27461
rect 33468 27421 33471 27455
rect 33505 27452 33517 27455
rect 33597 27455 33655 27461
rect 33505 27424 33561 27452
rect 33505 27421 33517 27424
rect 33468 27415 33517 27421
rect 33597 27421 33609 27455
rect 33643 27421 33655 27455
rect 33597 27415 33655 27421
rect 33468 27412 33474 27415
rect 33778 27412 33784 27464
rect 33836 27452 33842 27464
rect 34900 27461 34928 27492
rect 33873 27455 33931 27461
rect 33873 27452 33885 27455
rect 33836 27424 33885 27452
rect 33836 27412 33842 27424
rect 33873 27421 33885 27424
rect 33919 27421 33931 27455
rect 33873 27415 33931 27421
rect 34885 27455 34943 27461
rect 34885 27421 34897 27455
rect 34931 27421 34943 27455
rect 34885 27415 34943 27421
rect 26878 27393 26884 27396
rect 26528 27356 26832 27384
rect 26872 27347 26884 27393
rect 26936 27384 26942 27396
rect 26936 27356 26972 27384
rect 26878 27344 26884 27347
rect 26936 27344 26942 27356
rect 27154 27344 27160 27396
rect 27212 27384 27218 27396
rect 28718 27384 28724 27396
rect 27212 27356 28724 27384
rect 27212 27344 27218 27356
rect 28718 27344 28724 27356
rect 28776 27344 28782 27396
rect 28813 27387 28871 27393
rect 28813 27353 28825 27387
rect 28859 27353 28871 27387
rect 28813 27347 28871 27353
rect 32677 27387 32735 27393
rect 32677 27353 32689 27387
rect 32723 27384 32735 27387
rect 33134 27384 33140 27396
rect 32723 27356 33140 27384
rect 32723 27353 32735 27356
rect 32677 27347 32735 27353
rect 27614 27316 27620 27328
rect 25976 27288 27620 27316
rect 25777 27279 25835 27285
rect 27614 27276 27620 27288
rect 27672 27276 27678 27328
rect 27982 27316 27988 27328
rect 27943 27288 27988 27316
rect 27982 27276 27988 27288
rect 28040 27276 28046 27328
rect 28626 27276 28632 27328
rect 28684 27316 28690 27328
rect 28828 27316 28856 27347
rect 33134 27344 33140 27356
rect 33192 27384 33198 27396
rect 33689 27387 33747 27393
rect 33689 27384 33701 27387
rect 33192 27356 33701 27384
rect 33192 27344 33198 27356
rect 33689 27353 33701 27356
rect 33735 27353 33747 27387
rect 33689 27347 33747 27353
rect 34606 27344 34612 27396
rect 34664 27384 34670 27396
rect 34701 27387 34759 27393
rect 34701 27384 34713 27387
rect 34664 27356 34713 27384
rect 34664 27344 34670 27356
rect 34701 27353 34713 27356
rect 34747 27353 34759 27387
rect 34701 27347 34759 27353
rect 29549 27319 29607 27325
rect 29549 27316 29561 27319
rect 28684 27288 29561 27316
rect 28684 27276 28690 27288
rect 29549 27285 29561 27288
rect 29595 27316 29607 27319
rect 29638 27316 29644 27328
rect 29595 27288 29644 27316
rect 29595 27285 29607 27288
rect 29549 27279 29607 27285
rect 29638 27276 29644 27288
rect 29696 27276 29702 27328
rect 32306 27316 32312 27328
rect 32267 27288 32312 27316
rect 32306 27276 32312 27288
rect 32364 27276 32370 27328
rect 33321 27319 33379 27325
rect 33321 27285 33333 27319
rect 33367 27316 33379 27319
rect 33502 27316 33508 27328
rect 33367 27288 33508 27316
rect 33367 27285 33379 27288
rect 33321 27279 33379 27285
rect 33502 27276 33508 27288
rect 33560 27276 33566 27328
rect 34422 27276 34428 27328
rect 34480 27316 34486 27328
rect 35069 27319 35127 27325
rect 35069 27316 35081 27319
rect 34480 27288 35081 27316
rect 34480 27276 34486 27288
rect 35069 27285 35081 27288
rect 35115 27285 35127 27319
rect 35069 27279 35127 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 2685 27115 2743 27121
rect 2685 27081 2697 27115
rect 2731 27112 2743 27115
rect 2774 27112 2780 27124
rect 2731 27084 2780 27112
rect 2731 27081 2743 27084
rect 2685 27075 2743 27081
rect 2774 27072 2780 27084
rect 2832 27072 2838 27124
rect 4614 27072 4620 27124
rect 4672 27112 4678 27124
rect 6365 27115 6423 27121
rect 4672 27084 5212 27112
rect 4672 27072 4678 27084
rect 3329 27047 3387 27053
rect 3329 27013 3341 27047
rect 3375 27044 3387 27047
rect 3970 27044 3976 27056
rect 3375 27016 3976 27044
rect 3375 27013 3387 27016
rect 3329 27007 3387 27013
rect 3970 27004 3976 27016
rect 4028 27044 4034 27056
rect 5074 27044 5080 27056
rect 4028 27016 4936 27044
rect 5035 27016 5080 27044
rect 4028 27004 4034 27016
rect 3513 26979 3571 26985
rect 3513 26945 3525 26979
rect 3559 26945 3571 26979
rect 4798 26976 4804 26988
rect 4759 26948 4804 26976
rect 3513 26939 3571 26945
rect 3528 26908 3556 26939
rect 4798 26936 4804 26948
rect 4856 26936 4862 26988
rect 4908 26985 4936 27016
rect 5074 27004 5080 27016
rect 5132 27004 5138 27056
rect 5184 27053 5212 27084
rect 6365 27081 6377 27115
rect 6411 27112 6423 27115
rect 6454 27112 6460 27124
rect 6411 27084 6460 27112
rect 6411 27081 6423 27084
rect 6365 27075 6423 27081
rect 6454 27072 6460 27084
rect 6512 27072 6518 27124
rect 10137 27115 10195 27121
rect 10137 27081 10149 27115
rect 10183 27112 10195 27115
rect 11514 27112 11520 27124
rect 10183 27084 11100 27112
rect 11475 27084 11520 27112
rect 10183 27081 10195 27084
rect 10137 27075 10195 27081
rect 5169 27047 5227 27053
rect 5169 27013 5181 27047
rect 5215 27013 5227 27047
rect 5169 27007 5227 27013
rect 5442 27004 5448 27056
rect 5500 27044 5506 27056
rect 7098 27044 7104 27056
rect 5500 27016 7104 27044
rect 5500 27004 5506 27016
rect 7098 27004 7104 27016
rect 7156 27004 7162 27056
rect 7742 27004 7748 27056
rect 7800 27044 7806 27056
rect 10152 27044 10180 27075
rect 10962 27044 10968 27056
rect 7800 27016 10180 27044
rect 10923 27016 10968 27044
rect 7800 27004 7806 27016
rect 4894 26979 4952 26985
rect 4894 26945 4906 26979
rect 4940 26945 4952 26979
rect 4894 26939 4952 26945
rect 5307 26979 5365 26985
rect 5307 26945 5319 26979
rect 5353 26976 5365 26979
rect 5534 26976 5540 26988
rect 5353 26948 5540 26976
rect 5353 26945 5365 26948
rect 5307 26939 5365 26945
rect 5534 26936 5540 26948
rect 5592 26936 5598 26988
rect 7466 26976 7472 26988
rect 7524 26985 7530 26988
rect 7436 26948 7472 26976
rect 7466 26936 7472 26948
rect 7524 26939 7536 26985
rect 9306 26976 9312 26988
rect 9267 26948 9312 26976
rect 7524 26936 7530 26939
rect 9306 26936 9312 26948
rect 9364 26936 9370 26988
rect 9508 26985 9536 27016
rect 10962 27004 10968 27016
rect 11020 27004 11026 27056
rect 11072 27044 11100 27084
rect 11514 27072 11520 27084
rect 11572 27072 11578 27124
rect 16022 27112 16028 27124
rect 12406 27084 15516 27112
rect 15983 27084 16028 27112
rect 12406 27044 12434 27084
rect 15488 27053 15516 27084
rect 16022 27072 16028 27084
rect 16080 27072 16086 27124
rect 16850 27072 16856 27124
rect 16908 27112 16914 27124
rect 17037 27115 17095 27121
rect 17037 27112 17049 27115
rect 16908 27084 17049 27112
rect 16908 27072 16914 27084
rect 17037 27081 17049 27084
rect 17083 27112 17095 27115
rect 17402 27112 17408 27124
rect 17083 27084 17408 27112
rect 17083 27081 17095 27084
rect 17037 27075 17095 27081
rect 17402 27072 17408 27084
rect 17460 27072 17466 27124
rect 18414 27072 18420 27124
rect 18472 27112 18478 27124
rect 25590 27112 25596 27124
rect 18472 27084 25596 27112
rect 18472 27072 18478 27084
rect 25590 27072 25596 27084
rect 25648 27072 25654 27124
rect 25685 27115 25743 27121
rect 25685 27081 25697 27115
rect 25731 27112 25743 27115
rect 26878 27112 26884 27124
rect 25731 27084 26884 27112
rect 25731 27081 25743 27084
rect 25685 27075 25743 27081
rect 26878 27072 26884 27084
rect 26936 27072 26942 27124
rect 31386 27112 31392 27124
rect 29012 27084 31392 27112
rect 11072 27016 12434 27044
rect 15473 27047 15531 27053
rect 15473 27013 15485 27047
rect 15519 27044 15531 27047
rect 18432 27044 18460 27072
rect 15519 27016 18460 27044
rect 15519 27013 15531 27016
rect 15473 27007 15531 27013
rect 9493 26979 9551 26985
rect 9493 26945 9505 26979
rect 9539 26945 9551 26979
rect 9493 26939 9551 26945
rect 9858 26936 9864 26988
rect 9916 26976 9922 26988
rect 10781 26979 10839 26985
rect 10781 26976 10793 26979
rect 9916 26948 10793 26976
rect 9916 26936 9922 26948
rect 10781 26945 10793 26948
rect 10827 26945 10839 26979
rect 10781 26939 10839 26945
rect 12345 26979 12403 26985
rect 12345 26945 12357 26979
rect 12391 26976 12403 26979
rect 12618 26976 12624 26988
rect 12391 26948 12624 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 12618 26936 12624 26948
rect 12676 26936 12682 26988
rect 15948 26985 15976 27016
rect 19610 27004 19616 27056
rect 19668 27044 19674 27056
rect 20530 27044 20536 27056
rect 19668 27016 20536 27044
rect 19668 27004 19674 27016
rect 20530 27004 20536 27016
rect 20588 27004 20594 27056
rect 21174 27044 21180 27056
rect 21135 27016 21180 27044
rect 21174 27004 21180 27016
rect 21232 27044 21238 27056
rect 21910 27044 21916 27056
rect 21232 27016 21916 27044
rect 21232 27004 21238 27016
rect 21910 27004 21916 27016
rect 21968 27044 21974 27056
rect 24489 27047 24547 27053
rect 24489 27044 24501 27047
rect 21968 27016 24501 27044
rect 21968 27004 21974 27016
rect 24489 27013 24501 27016
rect 24535 27013 24547 27047
rect 24489 27007 24547 27013
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26945 15991 26979
rect 15933 26939 15991 26945
rect 16117 26979 16175 26985
rect 16117 26945 16129 26979
rect 16163 26976 16175 26979
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 16163 26948 16865 26976
rect 16163 26945 16175 26948
rect 16117 26939 16175 26945
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 5442 26908 5448 26920
rect 3528 26880 5448 26908
rect 5442 26868 5448 26880
rect 5500 26868 5506 26920
rect 7742 26868 7748 26920
rect 7800 26908 7806 26920
rect 9766 26908 9772 26920
rect 7800 26880 9772 26908
rect 7800 26868 7806 26880
rect 9766 26868 9772 26880
rect 9824 26908 9830 26920
rect 10594 26908 10600 26920
rect 9824 26880 10600 26908
rect 9824 26868 9830 26880
rect 10594 26868 10600 26880
rect 10652 26868 10658 26920
rect 11974 26868 11980 26920
rect 12032 26908 12038 26920
rect 12069 26911 12127 26917
rect 12069 26908 12081 26911
rect 12032 26880 12081 26908
rect 12032 26868 12038 26880
rect 12069 26877 12081 26880
rect 12115 26877 12127 26911
rect 12069 26871 12127 26877
rect 13354 26868 13360 26920
rect 13412 26908 13418 26920
rect 16132 26908 16160 26939
rect 13412 26880 16160 26908
rect 13412 26868 13418 26880
rect 16206 26868 16212 26920
rect 16264 26908 16270 26920
rect 16669 26911 16727 26917
rect 16669 26908 16681 26911
rect 16264 26880 16681 26908
rect 16264 26868 16270 26880
rect 16669 26877 16681 26880
rect 16715 26877 16727 26911
rect 16868 26908 16896 26939
rect 17586 26936 17592 26988
rect 17644 26976 17650 26988
rect 17773 26979 17831 26985
rect 17773 26976 17785 26979
rect 17644 26948 17785 26976
rect 17644 26936 17650 26948
rect 17773 26945 17785 26948
rect 17819 26976 17831 26979
rect 18138 26976 18144 26988
rect 17819 26948 18144 26976
rect 17819 26945 17831 26948
rect 17773 26939 17831 26945
rect 18138 26936 18144 26948
rect 18196 26976 18202 26988
rect 18417 26979 18475 26985
rect 18417 26976 18429 26979
rect 18196 26948 18429 26976
rect 18196 26936 18202 26948
rect 18417 26945 18429 26948
rect 18463 26945 18475 26979
rect 18417 26939 18475 26945
rect 19886 26936 19892 26988
rect 19944 26976 19950 26988
rect 22462 26985 22468 26988
rect 20174 26979 20232 26985
rect 20174 26976 20186 26979
rect 19944 26948 20186 26976
rect 19944 26936 19950 26948
rect 20174 26945 20186 26948
rect 20220 26945 20232 26979
rect 20174 26939 20232 26945
rect 22456 26939 22468 26985
rect 22520 26976 22526 26988
rect 22520 26948 22556 26976
rect 22462 26936 22468 26939
rect 22520 26936 22526 26948
rect 18230 26908 18236 26920
rect 16868 26880 18236 26908
rect 16669 26871 16727 26877
rect 18230 26868 18236 26880
rect 18288 26868 18294 26920
rect 20441 26911 20499 26917
rect 20441 26877 20453 26911
rect 20487 26908 20499 26911
rect 20530 26908 20536 26920
rect 20487 26880 20536 26908
rect 20487 26877 20499 26880
rect 20441 26871 20499 26877
rect 20530 26868 20536 26880
rect 20588 26908 20594 26920
rect 22189 26911 22247 26917
rect 22189 26908 22201 26911
rect 20588 26880 22201 26908
rect 20588 26868 20594 26880
rect 22189 26877 22201 26880
rect 22235 26877 22247 26911
rect 22189 26871 22247 26877
rect 3234 26800 3240 26852
rect 3292 26840 3298 26852
rect 4065 26843 4123 26849
rect 4065 26840 4077 26843
rect 3292 26812 4077 26840
rect 3292 26800 3298 26812
rect 4065 26809 4077 26812
rect 4111 26840 4123 26843
rect 4111 26812 6132 26840
rect 4111 26809 4123 26812
rect 4065 26803 4123 26809
rect 6104 26784 6132 26812
rect 8478 26800 8484 26852
rect 8536 26840 8542 26852
rect 9309 26843 9367 26849
rect 9309 26840 9321 26843
rect 8536 26812 9321 26840
rect 8536 26800 8542 26812
rect 9309 26809 9321 26812
rect 9355 26809 9367 26843
rect 9309 26803 9367 26809
rect 17957 26843 18015 26849
rect 17957 26809 17969 26843
rect 18003 26840 18015 26843
rect 18322 26840 18328 26852
rect 18003 26812 18328 26840
rect 18003 26809 18015 26812
rect 17957 26803 18015 26809
rect 18322 26800 18328 26812
rect 18380 26800 18386 26852
rect 3050 26732 3056 26784
rect 3108 26772 3114 26784
rect 3145 26775 3203 26781
rect 3145 26772 3157 26775
rect 3108 26744 3157 26772
rect 3108 26732 3114 26744
rect 3145 26741 3157 26744
rect 3191 26741 3203 26775
rect 5442 26772 5448 26784
rect 5403 26744 5448 26772
rect 3145 26735 3203 26741
rect 5442 26732 5448 26744
rect 5500 26732 5506 26784
rect 6086 26732 6092 26784
rect 6144 26772 6150 26784
rect 9950 26772 9956 26784
rect 6144 26744 9956 26772
rect 6144 26732 6150 26744
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 18690 26732 18696 26784
rect 18748 26772 18754 26784
rect 19061 26775 19119 26781
rect 19061 26772 19073 26775
rect 18748 26744 19073 26772
rect 18748 26732 18754 26744
rect 19061 26741 19073 26744
rect 19107 26741 19119 26775
rect 19061 26735 19119 26741
rect 22554 26732 22560 26784
rect 22612 26772 22618 26784
rect 23569 26775 23627 26781
rect 23569 26772 23581 26775
rect 22612 26744 23581 26772
rect 22612 26732 22618 26744
rect 23569 26741 23581 26744
rect 23615 26741 23627 26775
rect 24504 26772 24532 27007
rect 25774 27004 25780 27056
rect 25832 27044 25838 27056
rect 29012 27044 29040 27084
rect 31386 27072 31392 27084
rect 31444 27072 31450 27124
rect 32398 27072 32404 27124
rect 32456 27112 32462 27124
rect 34238 27112 34244 27124
rect 32456 27084 34244 27112
rect 32456 27072 32462 27084
rect 34238 27072 34244 27084
rect 34296 27072 34302 27124
rect 25832 27016 29040 27044
rect 25832 27004 25838 27016
rect 29086 27004 29092 27056
rect 29144 27044 29150 27056
rect 29144 27016 29868 27044
rect 29144 27004 29150 27016
rect 24670 26936 24676 26988
rect 24728 26976 24734 26988
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 24728 26948 25053 26976
rect 24728 26936 24734 26948
rect 25041 26945 25053 26948
rect 25087 26945 25099 26979
rect 25041 26939 25099 26945
rect 25204 26982 25262 26988
rect 25204 26948 25216 26982
rect 25250 26948 25262 26982
rect 25204 26942 25262 26948
rect 25317 26979 25375 26985
rect 25317 26945 25329 26979
rect 25363 26945 25375 26979
rect 25455 26979 25513 26985
rect 25455 26976 25467 26979
rect 24762 26868 24768 26920
rect 24820 26908 24826 26920
rect 25219 26908 25247 26942
rect 25317 26939 25375 26945
rect 25444 26945 25467 26976
rect 25501 26945 25513 26979
rect 25444 26939 25513 26945
rect 24820 26880 25247 26908
rect 24820 26868 24826 26880
rect 25130 26800 25136 26852
rect 25188 26840 25194 26852
rect 25335 26840 25363 26939
rect 25444 26908 25472 26939
rect 27706 26936 27712 26988
rect 27764 26976 27770 26988
rect 29282 26979 29340 26985
rect 29282 26976 29294 26979
rect 27764 26948 29294 26976
rect 27764 26936 27770 26948
rect 29282 26945 29294 26948
rect 29328 26945 29340 26979
rect 29840 26976 29868 27016
rect 31202 27004 31208 27056
rect 31260 27044 31266 27056
rect 31481 27047 31539 27053
rect 31481 27044 31493 27047
rect 31260 27016 31493 27044
rect 31260 27004 31266 27016
rect 31481 27013 31493 27016
rect 31527 27044 31539 27047
rect 35618 27044 35624 27056
rect 31527 27016 32812 27044
rect 31527 27013 31539 27016
rect 31481 27007 31539 27013
rect 32398 26976 32404 26988
rect 29840 26948 32404 26976
rect 29282 26939 29340 26945
rect 32398 26936 32404 26948
rect 32456 26936 32462 26988
rect 32582 26976 32588 26988
rect 32543 26948 32588 26976
rect 32582 26936 32588 26948
rect 32640 26936 32646 26988
rect 32784 26985 32812 27016
rect 34532 27016 35624 27044
rect 32677 26979 32735 26985
rect 32677 26945 32689 26979
rect 32723 26945 32735 26979
rect 32677 26939 32735 26945
rect 32769 26979 32827 26985
rect 32769 26945 32781 26979
rect 32815 26945 32827 26979
rect 34238 26976 34244 26988
rect 34199 26948 34244 26976
rect 32769 26939 32827 26945
rect 25188 26812 25363 26840
rect 25424 26880 25472 26908
rect 29549 26911 29607 26917
rect 25188 26800 25194 26812
rect 25424 26772 25452 26880
rect 29549 26877 29561 26911
rect 29595 26908 29607 26911
rect 31938 26908 31944 26920
rect 29595 26880 31944 26908
rect 29595 26877 29607 26880
rect 29549 26871 29607 26877
rect 31938 26868 31944 26880
rect 31996 26868 32002 26920
rect 32692 26908 32720 26939
rect 34238 26936 34244 26948
rect 34296 26936 34302 26988
rect 34422 26976 34428 26988
rect 34383 26948 34428 26976
rect 34422 26936 34428 26948
rect 34480 26936 34486 26988
rect 34532 26985 34560 27016
rect 35618 27004 35624 27016
rect 35676 27004 35682 27056
rect 34517 26979 34575 26985
rect 34517 26945 34529 26979
rect 34563 26945 34575 26979
rect 34517 26939 34575 26945
rect 34609 26979 34667 26985
rect 34609 26945 34621 26979
rect 34655 26945 34667 26979
rect 34609 26939 34667 26945
rect 39689 26979 39747 26985
rect 39689 26945 39701 26979
rect 39735 26976 39747 26979
rect 40494 26976 40500 26988
rect 39735 26948 40500 26976
rect 39735 26945 39747 26948
rect 39689 26939 39747 26945
rect 34532 26908 34560 26939
rect 32692 26880 34560 26908
rect 31846 26800 31852 26852
rect 31904 26840 31910 26852
rect 32692 26840 32720 26880
rect 31904 26812 32720 26840
rect 31904 26800 31910 26812
rect 32858 26800 32864 26852
rect 32916 26840 32922 26852
rect 33781 26843 33839 26849
rect 33781 26840 33793 26843
rect 32916 26812 33793 26840
rect 32916 26800 32922 26812
rect 33781 26809 33793 26812
rect 33827 26840 33839 26843
rect 34624 26840 34652 26939
rect 40494 26936 40500 26948
rect 40552 26936 40558 26988
rect 39942 26908 39948 26920
rect 39903 26880 39948 26908
rect 39942 26868 39948 26880
rect 40000 26868 40006 26920
rect 33827 26812 34652 26840
rect 33827 26809 33839 26812
rect 33781 26803 33839 26809
rect 24504 26744 25452 26772
rect 23569 26735 23627 26741
rect 25590 26732 25596 26784
rect 25648 26772 25654 26784
rect 25866 26772 25872 26784
rect 25648 26744 25872 26772
rect 25648 26732 25654 26744
rect 25866 26732 25872 26744
rect 25924 26772 25930 26784
rect 26145 26775 26203 26781
rect 26145 26772 26157 26775
rect 25924 26744 26157 26772
rect 25924 26732 25930 26744
rect 26145 26741 26157 26744
rect 26191 26741 26203 26775
rect 28166 26772 28172 26784
rect 28127 26744 28172 26772
rect 26145 26735 26203 26741
rect 28166 26732 28172 26744
rect 28224 26732 28230 26784
rect 33045 26775 33103 26781
rect 33045 26741 33057 26775
rect 33091 26772 33103 26775
rect 33594 26772 33600 26784
rect 33091 26744 33600 26772
rect 33091 26741 33103 26744
rect 33045 26735 33103 26741
rect 33594 26732 33600 26744
rect 33652 26732 33658 26784
rect 34885 26775 34943 26781
rect 34885 26741 34897 26775
rect 34931 26772 34943 26775
rect 35802 26772 35808 26784
rect 34931 26744 35808 26772
rect 34931 26741 34943 26744
rect 34885 26735 34943 26741
rect 35802 26732 35808 26744
rect 35860 26732 35866 26784
rect 37090 26732 37096 26784
rect 37148 26772 37154 26784
rect 38565 26775 38623 26781
rect 38565 26772 38577 26775
rect 37148 26744 38577 26772
rect 37148 26732 37154 26744
rect 38565 26741 38577 26744
rect 38611 26772 38623 26775
rect 40034 26772 40040 26784
rect 38611 26744 40040 26772
rect 38611 26741 38623 26744
rect 38565 26735 38623 26741
rect 40034 26732 40040 26744
rect 40092 26732 40098 26784
rect 58158 26772 58164 26784
rect 58119 26744 58164 26772
rect 58158 26732 58164 26744
rect 58216 26732 58222 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 5077 26571 5135 26577
rect 5077 26537 5089 26571
rect 5123 26568 5135 26571
rect 5718 26568 5724 26580
rect 5123 26540 5724 26568
rect 5123 26537 5135 26540
rect 5077 26531 5135 26537
rect 5718 26528 5724 26540
rect 5776 26528 5782 26580
rect 7285 26571 7343 26577
rect 7285 26537 7297 26571
rect 7331 26568 7343 26571
rect 7466 26568 7472 26580
rect 7331 26540 7472 26568
rect 7331 26537 7343 26540
rect 7285 26531 7343 26537
rect 7466 26528 7472 26540
rect 7524 26528 7530 26580
rect 11698 26568 11704 26580
rect 11659 26540 11704 26568
rect 11698 26528 11704 26540
rect 11756 26528 11762 26580
rect 18322 26528 18328 26580
rect 18380 26568 18386 26580
rect 19886 26568 19892 26580
rect 18380 26540 19784 26568
rect 19847 26540 19892 26568
rect 18380 26528 18386 26540
rect 5629 26503 5687 26509
rect 5629 26469 5641 26503
rect 5675 26500 5687 26503
rect 6086 26500 6092 26512
rect 5675 26472 6092 26500
rect 5675 26469 5687 26472
rect 5629 26463 5687 26469
rect 6086 26460 6092 26472
rect 6144 26460 6150 26512
rect 7558 26460 7564 26512
rect 7616 26460 7622 26512
rect 7650 26460 7656 26512
rect 7708 26500 7714 26512
rect 12621 26503 12679 26509
rect 7708 26472 7788 26500
rect 7708 26460 7714 26472
rect 3142 26432 3148 26444
rect 2976 26404 3148 26432
rect 2774 26324 2780 26376
rect 2832 26364 2838 26376
rect 2976 26373 3004 26404
rect 3142 26392 3148 26404
rect 3200 26432 3206 26444
rect 7576 26432 7604 26460
rect 3200 26404 7696 26432
rect 3200 26392 3206 26404
rect 2869 26367 2927 26373
rect 2869 26364 2881 26367
rect 2832 26336 2881 26364
rect 2832 26324 2838 26336
rect 2869 26333 2881 26336
rect 2915 26333 2927 26367
rect 2869 26327 2927 26333
rect 2961 26367 3019 26373
rect 2961 26333 2973 26367
rect 3007 26333 3019 26367
rect 2961 26327 3019 26333
rect 3050 26324 3056 26376
rect 3108 26364 3114 26376
rect 3108 26336 3153 26364
rect 3108 26324 3114 26336
rect 3234 26324 3240 26376
rect 3292 26364 3298 26376
rect 3973 26367 4031 26373
rect 3292 26336 3337 26364
rect 3292 26324 3298 26336
rect 3973 26333 3985 26367
rect 4019 26364 4031 26367
rect 4062 26364 4068 26376
rect 4019 26336 4068 26364
rect 4019 26333 4031 26336
rect 3973 26327 4031 26333
rect 4062 26324 4068 26336
rect 4120 26324 4126 26376
rect 6086 26364 6092 26376
rect 6047 26336 6092 26364
rect 6086 26324 6092 26336
rect 6144 26324 6150 26376
rect 6270 26364 6276 26376
rect 6231 26336 6276 26364
rect 6270 26324 6276 26336
rect 6328 26324 6334 26376
rect 6380 26373 6408 26404
rect 6365 26367 6423 26373
rect 6365 26333 6377 26367
rect 6411 26333 6423 26367
rect 6365 26327 6423 26333
rect 6457 26367 6515 26373
rect 6457 26333 6469 26367
rect 6503 26333 6515 26367
rect 6457 26327 6515 26333
rect 2593 26299 2651 26305
rect 2593 26265 2605 26299
rect 2639 26296 2651 26299
rect 4157 26299 4215 26305
rect 2639 26268 2774 26296
rect 2639 26265 2651 26268
rect 2593 26259 2651 26265
rect 2746 26228 2774 26268
rect 4157 26265 4169 26299
rect 4203 26296 4215 26299
rect 5350 26296 5356 26308
rect 4203 26268 5356 26296
rect 4203 26265 4215 26268
rect 4157 26259 4215 26265
rect 5350 26256 5356 26268
rect 5408 26256 5414 26308
rect 5718 26256 5724 26308
rect 5776 26296 5782 26308
rect 6472 26296 6500 26327
rect 7466 26324 7472 26376
rect 7524 26364 7530 26376
rect 7668 26373 7696 26404
rect 7760 26373 7788 26472
rect 12621 26469 12633 26503
rect 12667 26500 12679 26503
rect 14550 26500 14556 26512
rect 12667 26472 14556 26500
rect 12667 26469 12679 26472
rect 12621 26463 12679 26469
rect 14550 26460 14556 26472
rect 14608 26460 14614 26512
rect 18049 26503 18107 26509
rect 18049 26469 18061 26503
rect 18095 26500 18107 26503
rect 19334 26500 19340 26512
rect 18095 26472 19340 26500
rect 18095 26469 18107 26472
rect 18049 26463 18107 26469
rect 19334 26460 19340 26472
rect 19392 26460 19398 26512
rect 19756 26500 19784 26540
rect 19886 26528 19892 26540
rect 19944 26528 19950 26580
rect 22189 26571 22247 26577
rect 20640 26540 22140 26568
rect 20640 26500 20668 26540
rect 22112 26500 22140 26540
rect 22189 26537 22201 26571
rect 22235 26568 22247 26571
rect 22462 26568 22468 26580
rect 22235 26540 22468 26568
rect 22235 26537 22247 26540
rect 22189 26531 22247 26537
rect 22462 26528 22468 26540
rect 22520 26528 22526 26580
rect 24302 26528 24308 26580
rect 24360 26568 24366 26580
rect 28626 26568 28632 26580
rect 24360 26540 28632 26568
rect 24360 26528 24366 26540
rect 28626 26528 28632 26540
rect 28684 26528 28690 26580
rect 28721 26571 28779 26577
rect 28721 26537 28733 26571
rect 28767 26568 28779 26571
rect 28994 26568 29000 26580
rect 28767 26540 29000 26568
rect 28767 26537 28779 26540
rect 28721 26531 28779 26537
rect 28994 26528 29000 26540
rect 29052 26568 29058 26580
rect 30282 26568 30288 26580
rect 29052 26540 30288 26568
rect 29052 26528 29058 26540
rect 30282 26528 30288 26540
rect 30340 26568 30346 26580
rect 31481 26571 31539 26577
rect 31481 26568 31493 26571
rect 30340 26540 31493 26568
rect 30340 26528 30346 26540
rect 31481 26537 31493 26540
rect 31527 26568 31539 26571
rect 34698 26568 34704 26580
rect 31527 26540 31754 26568
rect 34659 26540 34704 26568
rect 31527 26537 31539 26540
rect 31481 26531 31539 26537
rect 24854 26500 24860 26512
rect 19756 26472 20668 26500
rect 20732 26472 21864 26500
rect 22112 26472 24624 26500
rect 17770 26392 17776 26444
rect 17828 26432 17834 26444
rect 20732 26432 20760 26472
rect 17828 26404 20760 26432
rect 17828 26392 17834 26404
rect 7561 26367 7619 26373
rect 7561 26364 7573 26367
rect 7524 26336 7573 26364
rect 7524 26324 7530 26336
rect 7561 26333 7573 26336
rect 7607 26333 7619 26367
rect 7561 26327 7619 26333
rect 7653 26367 7711 26373
rect 7653 26333 7665 26367
rect 7699 26333 7711 26367
rect 7653 26327 7711 26333
rect 7745 26367 7803 26373
rect 7745 26333 7757 26367
rect 7791 26333 7803 26367
rect 7745 26327 7803 26333
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26364 7987 26367
rect 8202 26364 8208 26376
rect 7975 26336 8208 26364
rect 7975 26333 7987 26336
rect 7929 26327 7987 26333
rect 8202 26324 8208 26336
rect 8260 26324 8266 26376
rect 9309 26367 9367 26373
rect 9309 26333 9321 26367
rect 9355 26364 9367 26367
rect 11514 26364 11520 26376
rect 9355 26336 11520 26364
rect 9355 26333 9367 26336
rect 9309 26327 9367 26333
rect 5776 26268 6500 26296
rect 5776 26256 5782 26268
rect 6546 26256 6552 26308
rect 6604 26296 6610 26308
rect 9324 26296 9352 26327
rect 11514 26324 11520 26336
rect 11572 26324 11578 26376
rect 16669 26367 16727 26373
rect 16669 26333 16681 26367
rect 16715 26364 16727 26367
rect 17402 26364 17408 26376
rect 16715 26336 17408 26364
rect 16715 26333 16727 26336
rect 16669 26327 16727 26333
rect 17402 26324 17408 26336
rect 17460 26324 17466 26376
rect 17954 26324 17960 26376
rect 18012 26364 18018 26376
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 18012 26336 19257 26364
rect 18012 26324 18018 26336
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 19426 26364 19432 26376
rect 19387 26336 19432 26364
rect 19245 26327 19303 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 19536 26373 19564 26404
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26333 19579 26367
rect 19521 26327 19579 26333
rect 19610 26324 19616 26376
rect 19668 26364 19674 26376
rect 20070 26364 20076 26376
rect 19668 26336 20076 26364
rect 19668 26324 19674 26336
rect 20070 26324 20076 26336
rect 20128 26324 20134 26376
rect 20438 26364 20444 26376
rect 20399 26336 20444 26364
rect 20438 26324 20444 26336
rect 20496 26324 20502 26376
rect 20622 26364 20628 26376
rect 20583 26336 20628 26364
rect 20622 26324 20628 26336
rect 20680 26324 20686 26376
rect 20732 26373 20760 26404
rect 20717 26367 20775 26373
rect 20717 26333 20729 26367
rect 20763 26333 20775 26367
rect 20717 26327 20775 26333
rect 20806 26324 20812 26376
rect 20864 26364 20870 26376
rect 21545 26367 21603 26373
rect 21545 26364 21557 26367
rect 20864 26336 20909 26364
rect 21008 26336 21557 26364
rect 20864 26324 20870 26336
rect 6604 26268 9352 26296
rect 11793 26299 11851 26305
rect 6604 26256 6610 26268
rect 11793 26265 11805 26299
rect 11839 26296 11851 26299
rect 11974 26296 11980 26308
rect 11839 26268 11980 26296
rect 11839 26265 11851 26268
rect 11793 26259 11851 26265
rect 11974 26256 11980 26268
rect 12032 26256 12038 26308
rect 12434 26256 12440 26308
rect 12492 26296 12498 26308
rect 16936 26299 16994 26305
rect 12492 26268 12537 26296
rect 12492 26256 12498 26268
rect 16936 26265 16948 26299
rect 16982 26296 16994 26299
rect 17310 26296 17316 26308
rect 16982 26268 17316 26296
rect 16982 26265 16994 26268
rect 16936 26259 16994 26265
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 20456 26296 20484 26324
rect 21008 26296 21036 26336
rect 21545 26333 21557 26336
rect 21591 26333 21603 26367
rect 21726 26364 21732 26376
rect 21687 26336 21732 26364
rect 21545 26327 21603 26333
rect 21726 26324 21732 26336
rect 21784 26324 21790 26376
rect 21836 26373 21864 26472
rect 22462 26392 22468 26444
rect 22520 26432 22526 26444
rect 23017 26435 23075 26441
rect 23017 26432 23029 26435
rect 22520 26404 23029 26432
rect 22520 26392 22526 26404
rect 23017 26401 23029 26404
rect 23063 26401 23075 26435
rect 23017 26395 23075 26401
rect 24596 26376 24624 26472
rect 24688 26472 24860 26500
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26333 21879 26367
rect 21821 26327 21879 26333
rect 21910 26324 21916 26376
rect 21968 26364 21974 26376
rect 21968 26336 22013 26364
rect 21968 26324 21974 26336
rect 22554 26324 22560 26376
rect 22612 26364 22618 26376
rect 22833 26367 22891 26373
rect 22833 26364 22845 26367
rect 22612 26336 22845 26364
rect 22612 26324 22618 26336
rect 22833 26333 22845 26336
rect 22879 26333 22891 26367
rect 24578 26364 24584 26376
rect 24491 26336 24584 26364
rect 22833 26327 22891 26333
rect 24578 26324 24584 26336
rect 24636 26324 24642 26376
rect 24688 26358 24716 26472
rect 24854 26460 24860 26472
rect 24912 26460 24918 26512
rect 27065 26503 27123 26509
rect 27065 26469 27077 26503
rect 27111 26469 27123 26503
rect 27065 26463 27123 26469
rect 25130 26432 25136 26444
rect 24872 26404 25136 26432
rect 24872 26373 24900 26404
rect 25130 26392 25136 26404
rect 25188 26392 25194 26444
rect 27080 26432 27108 26463
rect 27614 26432 27620 26444
rect 27080 26404 27620 26432
rect 27614 26392 27620 26404
rect 27672 26432 27678 26444
rect 28718 26432 28724 26444
rect 27672 26404 28724 26432
rect 27672 26392 27678 26404
rect 28718 26392 28724 26404
rect 28776 26392 28782 26444
rect 24857 26367 24915 26373
rect 24744 26361 24802 26367
rect 24744 26358 24756 26361
rect 24688 26330 24756 26358
rect 24744 26327 24756 26330
rect 24790 26327 24802 26361
rect 24857 26333 24869 26367
rect 24903 26333 24915 26367
rect 24857 26327 24915 26333
rect 24995 26367 25053 26373
rect 24995 26333 25007 26367
rect 25041 26364 25053 26367
rect 25590 26364 25596 26376
rect 25041 26336 25596 26364
rect 25041 26333 25053 26336
rect 24995 26327 25053 26333
rect 24744 26321 24802 26327
rect 25590 26324 25596 26336
rect 25648 26324 25654 26376
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26364 25743 26367
rect 26786 26364 26792 26376
rect 25731 26336 26792 26364
rect 25731 26333 25743 26336
rect 25685 26327 25743 26333
rect 26786 26324 26792 26336
rect 26844 26324 26850 26376
rect 31726 26364 31754 26540
rect 34698 26528 34704 26540
rect 34756 26528 34762 26580
rect 31938 26392 31944 26444
rect 31996 26432 32002 26444
rect 32033 26435 32091 26441
rect 32033 26432 32045 26435
rect 31996 26404 32045 26432
rect 31996 26392 32002 26404
rect 32033 26401 32045 26404
rect 32079 26401 32091 26435
rect 32033 26395 32091 26401
rect 33781 26367 33839 26373
rect 33781 26364 33793 26367
rect 31726 26336 33793 26364
rect 33781 26333 33793 26336
rect 33827 26333 33839 26367
rect 33781 26327 33839 26333
rect 35802 26324 35808 26376
rect 35860 26373 35866 26376
rect 35860 26364 35872 26373
rect 36081 26367 36139 26373
rect 35860 26336 35905 26364
rect 35860 26327 35872 26336
rect 36081 26333 36093 26367
rect 36127 26364 36139 26367
rect 37182 26364 37188 26376
rect 36127 26336 37188 26364
rect 36127 26333 36139 26336
rect 36081 26327 36139 26333
rect 35860 26324 35866 26327
rect 37182 26324 37188 26336
rect 37240 26324 37246 26376
rect 37366 26324 37372 26376
rect 37424 26364 37430 26376
rect 38933 26367 38991 26373
rect 38933 26364 38945 26367
rect 37424 26336 38945 26364
rect 37424 26324 37430 26336
rect 38933 26333 38945 26336
rect 38979 26364 38991 26367
rect 39301 26367 39359 26373
rect 38979 26336 39252 26364
rect 38979 26333 38991 26336
rect 38933 26327 38991 26333
rect 20456 26268 21036 26296
rect 21085 26299 21143 26305
rect 21085 26265 21097 26299
rect 21131 26296 21143 26299
rect 21634 26296 21640 26308
rect 21131 26268 21640 26296
rect 21131 26265 21143 26268
rect 21085 26259 21143 26265
rect 21634 26256 21640 26268
rect 21692 26256 21698 26308
rect 22649 26299 22707 26305
rect 22649 26265 22661 26299
rect 22695 26265 22707 26299
rect 22649 26259 22707 26265
rect 25225 26299 25283 26305
rect 25225 26265 25237 26299
rect 25271 26296 25283 26299
rect 25930 26299 25988 26305
rect 25930 26296 25942 26299
rect 25271 26268 25942 26296
rect 25271 26265 25283 26268
rect 25225 26259 25283 26265
rect 25930 26265 25942 26268
rect 25976 26265 25988 26299
rect 25930 26259 25988 26265
rect 2866 26228 2872 26240
rect 2746 26200 2872 26228
rect 2866 26188 2872 26200
rect 2924 26188 2930 26240
rect 3050 26188 3056 26240
rect 3108 26228 3114 26240
rect 3789 26231 3847 26237
rect 3789 26228 3801 26231
rect 3108 26200 3801 26228
rect 3108 26188 3114 26200
rect 3789 26197 3801 26200
rect 3835 26197 3847 26231
rect 6730 26228 6736 26240
rect 6691 26200 6736 26228
rect 3789 26191 3847 26197
rect 6730 26188 6736 26200
rect 6788 26188 6794 26240
rect 10594 26228 10600 26240
rect 10555 26200 10600 26228
rect 10594 26188 10600 26200
rect 10652 26188 10658 26240
rect 12342 26188 12348 26240
rect 12400 26228 12406 26240
rect 13081 26231 13139 26237
rect 13081 26228 13093 26231
rect 12400 26200 13093 26228
rect 12400 26188 12406 26200
rect 13081 26197 13093 26200
rect 13127 26197 13139 26231
rect 13081 26191 13139 26197
rect 20254 26188 20260 26240
rect 20312 26228 20318 26240
rect 21450 26228 21456 26240
rect 20312 26200 21456 26228
rect 20312 26188 20318 26200
rect 21450 26188 21456 26200
rect 21508 26228 21514 26240
rect 22664 26228 22692 26259
rect 26142 26256 26148 26308
rect 26200 26296 26206 26308
rect 27525 26299 27583 26305
rect 27525 26296 27537 26299
rect 26200 26268 27537 26296
rect 26200 26256 26206 26268
rect 27525 26265 27537 26268
rect 27571 26265 27583 26299
rect 27525 26259 27583 26265
rect 27709 26299 27767 26305
rect 27709 26265 27721 26299
rect 27755 26296 27767 26299
rect 28166 26296 28172 26308
rect 27755 26268 28172 26296
rect 27755 26265 27767 26268
rect 27709 26259 27767 26265
rect 28166 26256 28172 26268
rect 28224 26296 28230 26308
rect 29730 26296 29736 26308
rect 28224 26268 29736 26296
rect 28224 26256 28230 26268
rect 29730 26256 29736 26268
rect 29788 26256 29794 26308
rect 39114 26296 39120 26308
rect 39075 26268 39120 26296
rect 39114 26256 39120 26268
rect 39172 26256 39178 26308
rect 39224 26296 39252 26336
rect 39301 26333 39313 26367
rect 39347 26364 39359 26367
rect 40310 26364 40316 26376
rect 39347 26336 40316 26364
rect 39347 26333 39359 26336
rect 39301 26327 39359 26333
rect 40310 26324 40316 26336
rect 40368 26324 40374 26376
rect 39853 26299 39911 26305
rect 39853 26296 39865 26299
rect 39224 26268 39865 26296
rect 39853 26265 39865 26268
rect 39899 26265 39911 26299
rect 40034 26296 40040 26308
rect 39995 26268 40040 26296
rect 39853 26259 39911 26265
rect 40034 26256 40040 26268
rect 40092 26256 40098 26308
rect 21508 26200 22692 26228
rect 21508 26188 21514 26200
rect 25774 26188 25780 26240
rect 25832 26228 25838 26240
rect 27893 26231 27951 26237
rect 27893 26228 27905 26231
rect 25832 26200 27905 26228
rect 25832 26188 25838 26200
rect 27893 26197 27905 26200
rect 27939 26197 27951 26231
rect 27893 26191 27951 26197
rect 40221 26231 40279 26237
rect 40221 26197 40233 26231
rect 40267 26228 40279 26231
rect 41138 26228 41144 26240
rect 40267 26200 41144 26228
rect 40267 26197 40279 26200
rect 40221 26191 40279 26197
rect 41138 26188 41144 26200
rect 41196 26188 41202 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 3970 26024 3976 26036
rect 3931 25996 3976 26024
rect 3970 25984 3976 25996
rect 4028 25984 4034 26036
rect 5813 26027 5871 26033
rect 5813 25993 5825 26027
rect 5859 26024 5871 26027
rect 6270 26024 6276 26036
rect 5859 25996 6276 26024
rect 5859 25993 5871 25996
rect 5813 25987 5871 25993
rect 6270 25984 6276 25996
rect 6328 25984 6334 26036
rect 9490 25984 9496 26036
rect 9548 26024 9554 26036
rect 12434 26024 12440 26036
rect 9548 25996 12440 26024
rect 9548 25984 9554 25996
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 13541 26027 13599 26033
rect 13541 25993 13553 26027
rect 13587 26024 13599 26027
rect 13630 26024 13636 26036
rect 13587 25996 13636 26024
rect 13587 25993 13599 25996
rect 13541 25987 13599 25993
rect 13630 25984 13636 25996
rect 13688 25984 13694 26036
rect 17310 26024 17316 26036
rect 17271 25996 17316 26024
rect 17310 25984 17316 25996
rect 17368 25984 17374 26036
rect 17770 25984 17776 26036
rect 17828 25984 17834 26036
rect 18877 26027 18935 26033
rect 18877 25993 18889 26027
rect 18923 26024 18935 26027
rect 19426 26024 19432 26036
rect 18923 25996 19432 26024
rect 18923 25993 18935 25996
rect 18877 25987 18935 25993
rect 19426 25984 19432 25996
rect 19484 25984 19490 26036
rect 20622 25984 20628 26036
rect 20680 26024 20686 26036
rect 20901 26027 20959 26033
rect 20901 26024 20913 26027
rect 20680 25996 20913 26024
rect 20680 25984 20686 25996
rect 20901 25993 20913 25996
rect 20947 25993 20959 26027
rect 26237 26027 26295 26033
rect 20901 25987 20959 25993
rect 21008 25996 26197 26024
rect 2866 25965 2872 25968
rect 2860 25919 2872 25965
rect 2924 25956 2930 25968
rect 2924 25928 2960 25956
rect 2866 25916 2872 25919
rect 2924 25916 2930 25928
rect 5350 25916 5356 25968
rect 5408 25956 5414 25968
rect 5445 25959 5503 25965
rect 5445 25956 5457 25959
rect 5408 25928 5457 25956
rect 5408 25916 5414 25928
rect 5445 25925 5457 25928
rect 5491 25925 5503 25959
rect 5445 25919 5503 25925
rect 5629 25959 5687 25965
rect 5629 25925 5641 25959
rect 5675 25956 5687 25959
rect 7282 25956 7288 25968
rect 5675 25928 7052 25956
rect 7243 25928 7288 25956
rect 5675 25925 5687 25928
rect 5629 25919 5687 25925
rect 2590 25888 2596 25900
rect 2551 25860 2596 25888
rect 2590 25848 2596 25860
rect 2648 25848 2654 25900
rect 6914 25888 6920 25900
rect 6875 25860 6920 25888
rect 6914 25848 6920 25860
rect 6972 25848 6978 25900
rect 7024 25897 7052 25928
rect 7282 25916 7288 25928
rect 7340 25916 7346 25968
rect 9306 25956 9312 25968
rect 9267 25928 9312 25956
rect 9306 25916 9312 25928
rect 9364 25916 9370 25968
rect 9398 25916 9404 25968
rect 9456 25956 9462 25968
rect 17788 25956 17816 25984
rect 9456 25928 10364 25956
rect 9456 25916 9462 25928
rect 7010 25891 7068 25897
rect 7010 25857 7022 25891
rect 7056 25888 7068 25891
rect 7098 25888 7104 25900
rect 7056 25860 7104 25888
rect 7056 25857 7068 25860
rect 7010 25851 7068 25857
rect 7098 25848 7104 25860
rect 7156 25848 7162 25900
rect 7193 25891 7251 25897
rect 7193 25857 7205 25891
rect 7239 25857 7251 25891
rect 7193 25851 7251 25857
rect 7423 25891 7481 25897
rect 7423 25857 7435 25891
rect 7469 25888 7481 25891
rect 9324 25888 9352 25916
rect 7469 25860 9352 25888
rect 7469 25857 7481 25860
rect 7423 25851 7481 25857
rect 7208 25820 7236 25851
rect 9416 25820 9444 25916
rect 9490 25848 9496 25900
rect 9548 25888 9554 25900
rect 10336 25897 10364 25928
rect 17696 25928 17816 25956
rect 18509 25959 18567 25965
rect 10321 25891 10379 25897
rect 9548 25860 9593 25888
rect 9548 25848 9554 25860
rect 10321 25857 10333 25891
rect 10367 25857 10379 25891
rect 10321 25851 10379 25857
rect 11885 25891 11943 25897
rect 11885 25857 11897 25891
rect 11931 25888 11943 25891
rect 12342 25888 12348 25900
rect 11931 25860 12348 25888
rect 11931 25857 11943 25860
rect 11885 25851 11943 25857
rect 12342 25848 12348 25860
rect 12400 25848 12406 25900
rect 13262 25848 13268 25900
rect 13320 25888 13326 25900
rect 13633 25891 13691 25897
rect 13633 25888 13645 25891
rect 13320 25860 13645 25888
rect 13320 25848 13326 25860
rect 13633 25857 13645 25860
rect 13679 25857 13691 25891
rect 13633 25851 13691 25857
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25888 15715 25891
rect 16022 25888 16028 25900
rect 15703 25860 16028 25888
rect 15703 25857 15715 25860
rect 15657 25851 15715 25857
rect 16022 25848 16028 25860
rect 16080 25848 16086 25900
rect 16850 25888 16856 25900
rect 16811 25860 16856 25888
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 17126 25848 17132 25900
rect 17184 25888 17190 25900
rect 17494 25888 17500 25900
rect 17184 25860 17500 25888
rect 17184 25848 17190 25860
rect 17494 25848 17500 25860
rect 17552 25888 17558 25900
rect 17696 25897 17724 25928
rect 18509 25925 18521 25959
rect 18555 25956 18567 25959
rect 18782 25956 18788 25968
rect 18555 25928 18788 25956
rect 18555 25925 18567 25928
rect 18509 25919 18567 25925
rect 18782 25916 18788 25928
rect 18840 25956 18846 25968
rect 19705 25959 19763 25965
rect 19705 25956 19717 25959
rect 18840 25928 19717 25956
rect 18840 25916 18846 25928
rect 19705 25925 19717 25928
rect 19751 25956 19763 25959
rect 20254 25956 20260 25968
rect 19751 25928 20260 25956
rect 19751 25925 19763 25928
rect 19705 25919 19763 25925
rect 20254 25916 20260 25928
rect 20312 25916 20318 25968
rect 20441 25959 20499 25965
rect 20441 25925 20453 25959
rect 20487 25956 20499 25959
rect 20806 25956 20812 25968
rect 20487 25928 20812 25956
rect 20487 25925 20499 25928
rect 20441 25919 20499 25925
rect 20806 25916 20812 25928
rect 20864 25956 20870 25968
rect 21008 25956 21036 25996
rect 20864 25928 21036 25956
rect 21269 25959 21327 25965
rect 20864 25916 20870 25928
rect 21269 25925 21281 25959
rect 21315 25956 21327 25959
rect 21450 25956 21456 25968
rect 21315 25928 21456 25956
rect 21315 25925 21327 25928
rect 21269 25919 21327 25925
rect 21450 25916 21456 25928
rect 21508 25916 21514 25968
rect 21634 25916 21640 25968
rect 21692 25956 21698 25968
rect 22066 25959 22124 25965
rect 22066 25956 22078 25959
rect 21692 25928 22078 25956
rect 21692 25916 21698 25928
rect 22066 25925 22078 25928
rect 22112 25925 22124 25959
rect 22066 25919 22124 25925
rect 25130 25916 25136 25968
rect 25188 25956 25194 25968
rect 26169 25956 26197 25996
rect 26237 25993 26249 26027
rect 26283 26024 26295 26027
rect 27706 26024 27712 26036
rect 26283 25996 27712 26024
rect 26283 25993 26295 25996
rect 26237 25987 26295 25993
rect 27706 25984 27712 25996
rect 27764 25984 27770 26036
rect 32766 26024 32772 26036
rect 32727 25996 32772 26024
rect 32766 25984 32772 25996
rect 32824 25984 32830 26036
rect 37274 25984 37280 26036
rect 37332 26024 37338 26036
rect 38197 26027 38255 26033
rect 38197 26024 38209 26027
rect 37332 25996 38209 26024
rect 37332 25984 37338 25996
rect 38197 25993 38209 25996
rect 38243 26024 38255 26027
rect 38243 25996 38792 26024
rect 38243 25993 38255 25996
rect 38197 25987 38255 25993
rect 26973 25959 27031 25965
rect 26973 25956 26985 25959
rect 25188 25928 25912 25956
rect 25188 25916 25194 25928
rect 25884 25900 25912 25928
rect 26169 25928 26985 25956
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17552 25860 17601 25888
rect 17552 25848 17558 25860
rect 17589 25857 17601 25860
rect 17635 25857 17647 25891
rect 17589 25851 17647 25857
rect 17681 25891 17739 25897
rect 17681 25857 17693 25891
rect 17727 25857 17739 25891
rect 17681 25851 17739 25857
rect 17773 25891 17831 25897
rect 17773 25857 17785 25891
rect 17819 25857 17831 25891
rect 17773 25851 17831 25857
rect 17957 25891 18015 25897
rect 17957 25857 17969 25891
rect 18003 25888 18015 25891
rect 18138 25888 18144 25900
rect 18003 25860 18144 25888
rect 18003 25857 18015 25860
rect 17957 25851 18015 25857
rect 7208 25792 9444 25820
rect 9858 25780 9864 25832
rect 9916 25820 9922 25832
rect 10045 25823 10103 25829
rect 10045 25820 10057 25823
rect 9916 25792 10057 25820
rect 9916 25780 9922 25792
rect 10045 25789 10057 25792
rect 10091 25789 10103 25823
rect 10045 25783 10103 25789
rect 10870 25780 10876 25832
rect 10928 25820 10934 25832
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 10928 25792 12173 25820
rect 10928 25780 10934 25792
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 13722 25780 13728 25832
rect 13780 25820 13786 25832
rect 15381 25823 15439 25829
rect 15381 25820 15393 25823
rect 13780 25792 15393 25820
rect 13780 25780 13786 25792
rect 15381 25789 15393 25792
rect 15427 25789 15439 25823
rect 17788 25820 17816 25851
rect 18138 25848 18144 25860
rect 18196 25848 18202 25900
rect 18690 25888 18696 25900
rect 18651 25860 18696 25888
rect 18690 25848 18696 25860
rect 18748 25848 18754 25900
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19521 25891 19579 25897
rect 19521 25888 19533 25891
rect 19484 25860 19533 25888
rect 19484 25848 19490 25860
rect 19521 25857 19533 25860
rect 19567 25857 19579 25891
rect 19521 25851 19579 25857
rect 21085 25891 21143 25897
rect 21085 25857 21097 25891
rect 21131 25888 21143 25891
rect 21131 25860 22875 25888
rect 21131 25857 21143 25860
rect 21085 25851 21143 25857
rect 19337 25823 19395 25829
rect 19337 25820 19349 25823
rect 17788 25792 19349 25820
rect 15381 25783 15439 25789
rect 19337 25789 19349 25792
rect 19383 25789 19395 25823
rect 19337 25783 19395 25789
rect 20530 25780 20536 25832
rect 20588 25820 20594 25832
rect 21821 25823 21879 25829
rect 21821 25820 21833 25823
rect 20588 25792 21833 25820
rect 20588 25780 20594 25792
rect 21821 25789 21833 25792
rect 21867 25789 21879 25823
rect 21821 25783 21879 25789
rect 7561 25755 7619 25761
rect 7561 25721 7573 25755
rect 7607 25752 7619 25755
rect 8294 25752 8300 25764
rect 7607 25724 8300 25752
rect 7607 25721 7619 25724
rect 7561 25715 7619 25721
rect 8294 25712 8300 25724
rect 8352 25712 8358 25764
rect 17310 25712 17316 25764
rect 17368 25752 17374 25764
rect 19058 25752 19064 25764
rect 17368 25724 19064 25752
rect 17368 25712 17374 25724
rect 19058 25712 19064 25724
rect 19116 25712 19122 25764
rect 22847 25696 22875 25860
rect 24578 25848 24584 25900
rect 24636 25888 24642 25900
rect 24946 25888 24952 25900
rect 24636 25860 24952 25888
rect 24636 25848 24642 25860
rect 24946 25848 24952 25860
rect 25004 25888 25010 25900
rect 25774 25897 25780 25900
rect 25593 25891 25651 25897
rect 25593 25888 25605 25891
rect 25004 25860 25605 25888
rect 25004 25848 25010 25860
rect 25593 25857 25605 25860
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 25756 25891 25780 25897
rect 25756 25857 25768 25891
rect 25756 25851 25780 25857
rect 25774 25848 25780 25851
rect 25832 25848 25838 25900
rect 25866 25848 25872 25900
rect 25924 25888 25930 25900
rect 26007 25891 26065 25897
rect 25924 25860 25969 25888
rect 25924 25848 25930 25860
rect 26007 25857 26019 25891
rect 26053 25888 26065 25891
rect 26169 25888 26197 25928
rect 26973 25925 26985 25928
rect 27019 25956 27031 25959
rect 27062 25956 27068 25968
rect 27019 25928 27068 25956
rect 27019 25925 27031 25928
rect 26973 25919 27031 25925
rect 27062 25916 27068 25928
rect 27120 25916 27126 25968
rect 28626 25956 28632 25968
rect 28539 25928 28632 25956
rect 28626 25916 28632 25928
rect 28684 25956 28690 25968
rect 29825 25959 29883 25965
rect 29825 25956 29837 25959
rect 28684 25928 29837 25956
rect 28684 25916 28690 25928
rect 29825 25925 29837 25928
rect 29871 25925 29883 25959
rect 29825 25919 29883 25925
rect 33594 25916 33600 25968
rect 33652 25956 33658 25968
rect 38764 25965 38792 25996
rect 33882 25959 33940 25965
rect 33882 25956 33894 25959
rect 33652 25928 33894 25956
rect 33652 25916 33658 25928
rect 33882 25925 33894 25928
rect 33928 25925 33940 25959
rect 33882 25919 33940 25925
rect 38749 25959 38807 25965
rect 38749 25925 38761 25959
rect 38795 25925 38807 25959
rect 38749 25919 38807 25925
rect 26053 25860 26197 25888
rect 28813 25891 28871 25897
rect 26053 25857 26065 25860
rect 26007 25851 26065 25857
rect 28813 25857 28825 25891
rect 28859 25888 28871 25891
rect 28902 25888 28908 25900
rect 28859 25860 28908 25888
rect 28859 25857 28871 25860
rect 28813 25851 28871 25857
rect 28902 25848 28908 25860
rect 28960 25848 28966 25900
rect 30006 25888 30012 25900
rect 29967 25860 30012 25888
rect 30006 25848 30012 25860
rect 30064 25848 30070 25900
rect 34146 25820 34152 25832
rect 34107 25792 34152 25820
rect 34146 25780 34152 25792
rect 34204 25780 34210 25832
rect 37182 25712 37188 25764
rect 37240 25752 37246 25764
rect 39942 25752 39948 25764
rect 37240 25724 39948 25752
rect 37240 25712 37246 25724
rect 39942 25712 39948 25724
rect 40000 25752 40006 25764
rect 40037 25755 40095 25761
rect 40037 25752 40049 25755
rect 40000 25724 40049 25752
rect 40000 25712 40006 25724
rect 40037 25721 40049 25724
rect 40083 25721 40095 25755
rect 40037 25715 40095 25721
rect 6178 25644 6184 25696
rect 6236 25684 6242 25696
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 6236 25656 6377 25684
rect 6236 25644 6242 25656
rect 6365 25653 6377 25656
rect 6411 25684 6423 25687
rect 7466 25684 7472 25696
rect 6411 25656 7472 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 7466 25644 7472 25656
rect 7524 25644 7530 25696
rect 8113 25687 8171 25693
rect 8113 25653 8125 25687
rect 8159 25684 8171 25687
rect 8202 25684 8208 25696
rect 8159 25656 8208 25684
rect 8159 25653 8171 25656
rect 8113 25647 8171 25653
rect 8202 25644 8208 25656
rect 8260 25644 8266 25696
rect 15010 25644 15016 25696
rect 15068 25684 15074 25696
rect 16669 25687 16727 25693
rect 16669 25684 16681 25687
rect 15068 25656 16681 25684
rect 15068 25644 15074 25656
rect 16669 25653 16681 25656
rect 16715 25653 16727 25687
rect 16669 25647 16727 25653
rect 17218 25644 17224 25696
rect 17276 25684 17282 25696
rect 18138 25684 18144 25696
rect 17276 25656 18144 25684
rect 17276 25644 17282 25656
rect 18138 25644 18144 25656
rect 18196 25684 18202 25696
rect 20438 25684 20444 25696
rect 18196 25656 20444 25684
rect 18196 25644 18202 25656
rect 20438 25644 20444 25656
rect 20496 25644 20502 25696
rect 22830 25684 22836 25696
rect 22743 25656 22836 25684
rect 22830 25644 22836 25656
rect 22888 25684 22894 25696
rect 23201 25687 23259 25693
rect 23201 25684 23213 25687
rect 22888 25656 23213 25684
rect 22888 25644 22894 25656
rect 23201 25653 23213 25656
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 28997 25687 29055 25693
rect 28997 25653 29009 25687
rect 29043 25684 29055 25687
rect 29546 25684 29552 25696
rect 29043 25656 29552 25684
rect 29043 25653 29055 25656
rect 28997 25647 29055 25653
rect 29546 25644 29552 25656
rect 29604 25644 29610 25696
rect 30193 25687 30251 25693
rect 30193 25653 30205 25687
rect 30239 25684 30251 25687
rect 30466 25684 30472 25696
rect 30239 25656 30472 25684
rect 30239 25653 30251 25656
rect 30193 25647 30251 25653
rect 30466 25644 30472 25656
rect 30524 25644 30530 25696
rect 31113 25687 31171 25693
rect 31113 25653 31125 25687
rect 31159 25684 31171 25687
rect 31294 25684 31300 25696
rect 31159 25656 31300 25684
rect 31159 25653 31171 25656
rect 31113 25647 31171 25653
rect 31294 25644 31300 25656
rect 31352 25644 31358 25696
rect 37461 25687 37519 25693
rect 37461 25653 37473 25687
rect 37507 25684 37519 25687
rect 37826 25684 37832 25696
rect 37507 25656 37832 25684
rect 37507 25653 37519 25656
rect 37461 25647 37519 25653
rect 37826 25644 37832 25656
rect 37884 25644 37890 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 7098 25440 7104 25492
rect 7156 25480 7162 25492
rect 7745 25483 7803 25489
rect 7745 25480 7757 25483
rect 7156 25452 7757 25480
rect 7156 25440 7162 25452
rect 7745 25449 7757 25452
rect 7791 25449 7803 25483
rect 7745 25443 7803 25449
rect 16298 25440 16304 25492
rect 16356 25480 16362 25492
rect 22186 25480 22192 25492
rect 16356 25452 22192 25480
rect 16356 25440 16362 25452
rect 22186 25440 22192 25452
rect 22244 25480 22250 25492
rect 24670 25480 24676 25492
rect 22244 25452 24676 25480
rect 22244 25440 22250 25452
rect 24670 25440 24676 25452
rect 24728 25440 24734 25492
rect 24762 25440 24768 25492
rect 24820 25480 24826 25492
rect 25777 25483 25835 25489
rect 25777 25480 25789 25483
rect 24820 25452 25789 25480
rect 24820 25440 24826 25452
rect 25777 25449 25789 25452
rect 25823 25449 25835 25483
rect 25777 25443 25835 25449
rect 31294 25440 31300 25492
rect 31352 25480 31358 25492
rect 39209 25483 39267 25489
rect 39209 25480 39221 25483
rect 31352 25452 39221 25480
rect 31352 25440 31358 25452
rect 39209 25449 39221 25452
rect 39255 25449 39267 25483
rect 39850 25480 39856 25492
rect 39811 25452 39856 25480
rect 39209 25443 39267 25449
rect 9950 25372 9956 25424
rect 10008 25412 10014 25424
rect 10597 25415 10655 25421
rect 10597 25412 10609 25415
rect 10008 25384 10609 25412
rect 10008 25372 10014 25384
rect 10597 25381 10609 25384
rect 10643 25381 10655 25415
rect 20070 25412 20076 25424
rect 20031 25384 20076 25412
rect 10597 25375 10655 25381
rect 20070 25372 20076 25384
rect 20128 25372 20134 25424
rect 21542 25372 21548 25424
rect 21600 25412 21606 25424
rect 27798 25412 27804 25424
rect 21600 25384 27804 25412
rect 21600 25372 21606 25384
rect 27798 25372 27804 25384
rect 27856 25372 27862 25424
rect 30006 25412 30012 25424
rect 28966 25384 30012 25412
rect 2133 25347 2191 25353
rect 2133 25313 2145 25347
rect 2179 25344 2191 25347
rect 3142 25344 3148 25356
rect 2179 25316 2912 25344
rect 2179 25313 2191 25316
rect 2133 25307 2191 25313
rect 2884 25288 2912 25316
rect 2976 25316 3148 25344
rect 2590 25236 2596 25288
rect 2648 25236 2654 25288
rect 2866 25276 2872 25288
rect 2827 25248 2872 25276
rect 2866 25236 2872 25248
rect 2924 25236 2930 25288
rect 2976 25285 3004 25316
rect 3142 25304 3148 25316
rect 3200 25304 3206 25356
rect 11790 25304 11796 25356
rect 11848 25344 11854 25356
rect 15841 25347 15899 25353
rect 15841 25344 15853 25347
rect 11848 25316 15853 25344
rect 11848 25304 11854 25316
rect 15841 25313 15853 25316
rect 15887 25344 15899 25347
rect 17586 25344 17592 25356
rect 15887 25316 17592 25344
rect 15887 25313 15899 25316
rect 15841 25307 15899 25313
rect 17586 25304 17592 25316
rect 17644 25304 17650 25356
rect 18049 25347 18107 25353
rect 18049 25313 18061 25347
rect 18095 25344 18107 25347
rect 18230 25344 18236 25356
rect 18095 25316 18236 25344
rect 18095 25313 18107 25316
rect 18049 25307 18107 25313
rect 18230 25304 18236 25316
rect 18288 25304 18294 25356
rect 18325 25347 18383 25353
rect 18325 25313 18337 25347
rect 18371 25344 18383 25347
rect 18414 25344 18420 25356
rect 18371 25316 18420 25344
rect 18371 25313 18383 25316
rect 18325 25307 18383 25313
rect 18414 25304 18420 25316
rect 18472 25344 18478 25356
rect 19242 25344 19248 25356
rect 18472 25316 19248 25344
rect 18472 25304 18478 25316
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 28966 25344 28994 25384
rect 30006 25372 30012 25384
rect 30064 25412 30070 25424
rect 31389 25415 31447 25421
rect 31389 25412 31401 25415
rect 30064 25384 31401 25412
rect 30064 25372 30070 25384
rect 31389 25381 31401 25384
rect 31435 25381 31447 25415
rect 39224 25412 39252 25443
rect 39850 25440 39856 25452
rect 39908 25440 39914 25492
rect 40494 25440 40500 25492
rect 40552 25480 40558 25492
rect 41601 25483 41659 25489
rect 41601 25480 41613 25483
rect 40552 25452 41613 25480
rect 40552 25440 40558 25452
rect 41601 25449 41613 25452
rect 41647 25449 41659 25483
rect 41601 25443 41659 25449
rect 40126 25412 40132 25424
rect 39224 25384 40132 25412
rect 31389 25375 31447 25381
rect 40126 25372 40132 25384
rect 40184 25372 40190 25424
rect 40862 25344 40868 25356
rect 21836 25316 28994 25344
rect 37936 25316 40868 25344
rect 2961 25279 3019 25285
rect 2961 25245 2973 25279
rect 3007 25245 3019 25279
rect 2961 25239 3019 25245
rect 3050 25236 3056 25288
rect 3108 25276 3114 25288
rect 3108 25248 3153 25276
rect 3108 25236 3114 25248
rect 3234 25236 3240 25288
rect 3292 25276 3298 25288
rect 6365 25279 6423 25285
rect 3292 25248 3337 25276
rect 3292 25236 3298 25248
rect 6365 25245 6377 25279
rect 6411 25276 6423 25279
rect 7742 25276 7748 25288
rect 6411 25248 7748 25276
rect 6411 25245 6423 25248
rect 6365 25239 6423 25245
rect 7742 25236 7748 25248
rect 7800 25236 7806 25288
rect 10781 25279 10839 25285
rect 10781 25245 10793 25279
rect 10827 25276 10839 25279
rect 10870 25276 10876 25288
rect 10827 25248 10876 25276
rect 10827 25245 10839 25248
rect 10781 25239 10839 25245
rect 10870 25236 10876 25248
rect 10928 25276 10934 25288
rect 11517 25279 11575 25285
rect 11517 25276 11529 25279
rect 10928 25248 11529 25276
rect 10928 25236 10934 25248
rect 11517 25245 11529 25248
rect 11563 25245 11575 25279
rect 11517 25239 11575 25245
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 15657 25279 15715 25285
rect 15657 25276 15669 25279
rect 12400 25248 15669 25276
rect 12400 25236 12406 25248
rect 15657 25245 15669 25248
rect 15703 25276 15715 25279
rect 16301 25279 16359 25285
rect 16301 25276 16313 25279
rect 15703 25248 16313 25276
rect 15703 25245 15715 25248
rect 15657 25239 15715 25245
rect 16301 25245 16313 25248
rect 16347 25245 16359 25279
rect 16301 25239 16359 25245
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 18748 25248 20208 25276
rect 18748 25236 18754 25248
rect 2608 25208 2636 25236
rect 4157 25211 4215 25217
rect 4157 25208 4169 25211
rect 2608 25180 4169 25208
rect 4157 25177 4169 25180
rect 4203 25177 4215 25211
rect 4157 25171 4215 25177
rect 5905 25211 5963 25217
rect 5905 25177 5917 25211
rect 5951 25208 5963 25211
rect 6454 25208 6460 25220
rect 5951 25180 6460 25208
rect 5951 25177 5963 25180
rect 5905 25171 5963 25177
rect 6454 25168 6460 25180
rect 6512 25168 6518 25220
rect 6632 25211 6690 25217
rect 6632 25177 6644 25211
rect 6678 25208 6690 25211
rect 6730 25208 6736 25220
rect 6678 25180 6736 25208
rect 6678 25177 6690 25180
rect 6632 25171 6690 25177
rect 6730 25168 6736 25180
rect 6788 25168 6794 25220
rect 14921 25211 14979 25217
rect 14921 25177 14933 25211
rect 14967 25177 14979 25211
rect 14921 25171 14979 25177
rect 2593 25143 2651 25149
rect 2593 25109 2605 25143
rect 2639 25140 2651 25143
rect 2866 25140 2872 25152
rect 2639 25112 2872 25140
rect 2639 25109 2651 25112
rect 2593 25103 2651 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 11422 25140 11428 25152
rect 11383 25112 11428 25140
rect 11422 25100 11428 25112
rect 11480 25100 11486 25152
rect 13262 25140 13268 25152
rect 13223 25112 13268 25140
rect 13262 25100 13268 25112
rect 13320 25100 13326 25152
rect 14642 25100 14648 25152
rect 14700 25140 14706 25152
rect 14737 25143 14795 25149
rect 14737 25140 14749 25143
rect 14700 25112 14749 25140
rect 14700 25100 14706 25112
rect 14737 25109 14749 25112
rect 14783 25109 14795 25143
rect 14936 25140 14964 25171
rect 15010 25168 15016 25220
rect 15068 25208 15074 25220
rect 15105 25211 15163 25217
rect 15105 25208 15117 25211
rect 15068 25180 15117 25208
rect 15068 25168 15074 25180
rect 15105 25177 15117 25180
rect 15151 25177 15163 25211
rect 20180 25208 20208 25248
rect 21358 25236 21364 25288
rect 21416 25276 21422 25288
rect 21836 25285 21864 25316
rect 21683 25279 21741 25285
rect 21683 25276 21695 25279
rect 21416 25248 21695 25276
rect 21416 25236 21422 25248
rect 21683 25245 21695 25248
rect 21729 25245 21741 25279
rect 21683 25239 21741 25245
rect 21821 25279 21879 25285
rect 21821 25245 21833 25279
rect 21867 25245 21879 25279
rect 21821 25239 21879 25245
rect 22051 25279 22109 25285
rect 22051 25245 22063 25279
rect 22097 25245 22109 25279
rect 22051 25239 22109 25245
rect 22189 25279 22247 25285
rect 22189 25245 22201 25279
rect 22235 25276 22247 25279
rect 22646 25276 22652 25288
rect 22235 25248 22652 25276
rect 22235 25245 22247 25248
rect 22189 25239 22247 25245
rect 21910 25208 21916 25220
rect 20180 25180 21680 25208
rect 21871 25180 21916 25208
rect 15105 25171 15163 25177
rect 15562 25140 15568 25152
rect 14936 25112 15568 25140
rect 14737 25103 14795 25109
rect 15562 25100 15568 25112
rect 15620 25100 15626 25152
rect 17037 25143 17095 25149
rect 17037 25109 17049 25143
rect 17083 25140 17095 25143
rect 17126 25140 17132 25152
rect 17083 25112 17132 25140
rect 17083 25109 17095 25112
rect 17037 25103 17095 25109
rect 17126 25100 17132 25112
rect 17184 25100 17190 25152
rect 19334 25100 19340 25152
rect 19392 25140 19398 25152
rect 19392 25112 19437 25140
rect 19392 25100 19398 25112
rect 20806 25100 20812 25152
rect 20864 25140 20870 25152
rect 21545 25143 21603 25149
rect 21545 25140 21557 25143
rect 20864 25112 21557 25140
rect 20864 25100 20870 25112
rect 21545 25109 21557 25112
rect 21591 25109 21603 25143
rect 21652 25140 21680 25180
rect 21910 25168 21916 25180
rect 21968 25168 21974 25220
rect 22066 25140 22094 25239
rect 22646 25236 22652 25248
rect 22704 25236 22710 25288
rect 25222 25236 25228 25288
rect 25280 25276 25286 25288
rect 26142 25276 26148 25288
rect 25280 25248 26148 25276
rect 25280 25236 25286 25248
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 28537 25279 28595 25285
rect 28537 25245 28549 25279
rect 28583 25276 28595 25279
rect 28994 25276 29000 25288
rect 28583 25248 29000 25276
rect 28583 25245 28595 25248
rect 28537 25239 28595 25245
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 30285 25279 30343 25285
rect 30285 25276 30297 25279
rect 29840 25248 30297 25276
rect 25961 25211 26019 25217
rect 25961 25177 25973 25211
rect 26007 25177 26019 25211
rect 26786 25208 26792 25220
rect 26747 25180 26792 25208
rect 25961 25171 26019 25177
rect 21652 25112 22094 25140
rect 25976 25140 26004 25171
rect 26786 25168 26792 25180
rect 26844 25168 26850 25220
rect 29840 25152 29868 25248
rect 30285 25245 30297 25248
rect 30331 25245 30343 25279
rect 30466 25276 30472 25288
rect 30427 25248 30472 25276
rect 30285 25239 30343 25245
rect 30466 25236 30472 25248
rect 30524 25236 30530 25288
rect 30558 25236 30564 25288
rect 30616 25276 30622 25288
rect 30699 25279 30757 25285
rect 30616 25248 30661 25276
rect 30616 25236 30622 25248
rect 30699 25245 30711 25279
rect 30745 25276 30757 25279
rect 31294 25276 31300 25288
rect 30745 25248 31300 25276
rect 30745 25245 30757 25248
rect 30699 25239 30757 25245
rect 31294 25236 31300 25248
rect 31352 25236 31358 25288
rect 31938 25236 31944 25288
rect 31996 25276 32002 25288
rect 32769 25279 32827 25285
rect 32769 25276 32781 25279
rect 31996 25248 32781 25276
rect 31996 25236 32002 25248
rect 32769 25245 32781 25248
rect 32815 25276 32827 25279
rect 34146 25276 34152 25288
rect 32815 25248 34152 25276
rect 32815 25245 32827 25248
rect 32769 25239 32827 25245
rect 34146 25236 34152 25248
rect 34204 25236 34210 25288
rect 37093 25279 37151 25285
rect 37093 25245 37105 25279
rect 37139 25276 37151 25279
rect 37182 25276 37188 25288
rect 37139 25248 37188 25276
rect 37139 25245 37151 25248
rect 37093 25239 37151 25245
rect 37182 25236 37188 25248
rect 37240 25236 37246 25288
rect 37826 25276 37832 25288
rect 37787 25248 37832 25276
rect 37826 25236 37832 25248
rect 37884 25236 37890 25288
rect 37936 25285 37964 25316
rect 37921 25279 37979 25285
rect 37921 25245 37933 25279
rect 37967 25245 37979 25279
rect 37921 25239 37979 25245
rect 38010 25236 38016 25288
rect 38068 25276 38074 25288
rect 38197 25279 38255 25285
rect 38068 25248 38113 25276
rect 38068 25236 38074 25248
rect 38197 25245 38209 25279
rect 38243 25245 38255 25279
rect 40126 25276 40132 25288
rect 40087 25248 40132 25276
rect 38197 25239 38255 25245
rect 30929 25211 30987 25217
rect 30929 25177 30941 25211
rect 30975 25208 30987 25211
rect 32502 25211 32560 25217
rect 32502 25208 32514 25211
rect 30975 25180 32514 25208
rect 30975 25177 30987 25180
rect 30929 25171 30987 25177
rect 32502 25177 32514 25180
rect 32548 25177 32560 25211
rect 32502 25171 32560 25177
rect 36848 25211 36906 25217
rect 36848 25177 36860 25211
rect 36894 25208 36906 25211
rect 37553 25211 37611 25217
rect 37553 25208 37565 25211
rect 36894 25180 37565 25208
rect 36894 25177 36906 25180
rect 36848 25171 36906 25177
rect 37553 25177 37565 25180
rect 37599 25177 37611 25211
rect 38212 25208 38240 25239
rect 40126 25236 40132 25248
rect 40184 25236 40190 25288
rect 40236 25285 40264 25316
rect 40862 25304 40868 25316
rect 40920 25344 40926 25356
rect 40920 25316 41276 25344
rect 40920 25304 40926 25316
rect 40221 25279 40279 25285
rect 40221 25245 40233 25279
rect 40267 25245 40279 25279
rect 40221 25239 40279 25245
rect 40310 25236 40316 25288
rect 40368 25276 40374 25288
rect 40497 25279 40555 25285
rect 40368 25248 40413 25276
rect 40368 25236 40374 25248
rect 40497 25245 40509 25279
rect 40543 25276 40555 25279
rect 40957 25279 41015 25285
rect 40957 25276 40969 25279
rect 40543 25248 40969 25276
rect 40543 25245 40555 25248
rect 40497 25239 40555 25245
rect 40957 25245 40969 25248
rect 41003 25245 41015 25279
rect 41138 25276 41144 25288
rect 41099 25248 41144 25276
rect 40957 25239 41015 25245
rect 39758 25208 39764 25220
rect 38212 25180 39764 25208
rect 37553 25171 37611 25177
rect 39758 25168 39764 25180
rect 39816 25208 39822 25220
rect 40512 25208 40540 25239
rect 41138 25236 41144 25248
rect 41196 25236 41202 25288
rect 41248 25282 41276 25316
rect 41233 25276 41291 25282
rect 41233 25242 41245 25276
rect 41279 25242 41291 25276
rect 41233 25236 41291 25242
rect 41371 25279 41429 25285
rect 41371 25245 41383 25279
rect 41417 25245 41429 25279
rect 58158 25276 58164 25288
rect 58119 25248 58164 25276
rect 41371 25239 41429 25245
rect 39816 25180 40540 25208
rect 39816 25168 39822 25180
rect 27982 25140 27988 25152
rect 25976 25112 27988 25140
rect 21545 25103 21603 25109
rect 27982 25100 27988 25112
rect 28040 25140 28046 25152
rect 28994 25140 29000 25152
rect 28040 25112 29000 25140
rect 28040 25100 28046 25112
rect 28994 25100 29000 25112
rect 29052 25100 29058 25152
rect 29822 25140 29828 25152
rect 29783 25112 29828 25140
rect 29822 25100 29828 25112
rect 29880 25100 29886 25152
rect 35713 25143 35771 25149
rect 35713 25109 35725 25143
rect 35759 25140 35771 25143
rect 36170 25140 36176 25152
rect 35759 25112 36176 25140
rect 35759 25109 35771 25112
rect 35713 25103 35771 25109
rect 36170 25100 36176 25112
rect 36228 25100 36234 25152
rect 41230 25100 41236 25152
rect 41288 25140 41294 25152
rect 41386 25140 41414 25239
rect 58158 25236 58164 25248
rect 58216 25236 58222 25288
rect 41288 25112 41414 25140
rect 41288 25100 41294 25112
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 6457 24939 6515 24945
rect 6457 24905 6469 24939
rect 6503 24936 6515 24939
rect 6546 24936 6552 24948
rect 6503 24908 6552 24936
rect 6503 24905 6515 24908
rect 6457 24899 6515 24905
rect 6546 24896 6552 24908
rect 6604 24896 6610 24948
rect 8202 24896 8208 24948
rect 8260 24936 8266 24948
rect 11422 24936 11428 24948
rect 8260 24908 11428 24936
rect 8260 24896 8266 24908
rect 11422 24896 11428 24908
rect 11480 24936 11486 24948
rect 16298 24936 16304 24948
rect 11480 24908 16304 24936
rect 11480 24896 11486 24908
rect 16298 24896 16304 24908
rect 16356 24896 16362 24948
rect 19334 24936 19340 24948
rect 18984 24908 19340 24936
rect 2866 24877 2872 24880
rect 2860 24831 2872 24877
rect 2924 24868 2930 24880
rect 9674 24868 9680 24880
rect 2924 24840 2960 24868
rect 2866 24828 2872 24831
rect 2924 24828 2930 24840
rect 9646 24828 9680 24868
rect 9732 24828 9738 24880
rect 15378 24868 15384 24880
rect 12817 24840 15384 24868
rect 2590 24800 2596 24812
rect 2551 24772 2596 24800
rect 2590 24760 2596 24772
rect 2648 24760 2654 24812
rect 3326 24760 3332 24812
rect 3384 24800 3390 24812
rect 6270 24800 6276 24812
rect 3384 24772 6276 24800
rect 3384 24760 3390 24772
rect 6270 24760 6276 24772
rect 6328 24760 6334 24812
rect 7006 24760 7012 24812
rect 7064 24800 7070 24812
rect 9646 24800 9674 24828
rect 9841 24803 9899 24809
rect 9841 24800 9853 24803
rect 7064 24772 9674 24800
rect 9784 24772 9853 24800
rect 7064 24760 7070 24772
rect 7926 24692 7932 24744
rect 7984 24732 7990 24744
rect 8202 24732 8208 24744
rect 7984 24704 8208 24732
rect 7984 24692 7990 24704
rect 8202 24692 8208 24704
rect 8260 24692 8266 24744
rect 9030 24692 9036 24744
rect 9088 24732 9094 24744
rect 9784 24732 9812 24772
rect 9841 24769 9853 24772
rect 9887 24769 9899 24803
rect 9841 24763 9899 24769
rect 9931 24760 9937 24812
rect 9989 24809 9995 24812
rect 9989 24803 10008 24809
rect 9996 24769 10008 24803
rect 9989 24763 10008 24769
rect 10050 24803 10108 24809
rect 10050 24769 10062 24803
rect 10096 24800 10108 24803
rect 10229 24803 10287 24809
rect 10096 24772 10180 24800
rect 10096 24769 10108 24772
rect 10050 24763 10108 24769
rect 9989 24760 9995 24763
rect 9088 24704 9812 24732
rect 10152 24732 10180 24772
rect 10229 24769 10241 24803
rect 10275 24800 10287 24803
rect 10318 24800 10324 24812
rect 10275 24772 10324 24800
rect 10275 24769 10287 24772
rect 10229 24763 10287 24769
rect 10318 24760 10324 24772
rect 10376 24800 10382 24812
rect 12817 24800 12845 24840
rect 15378 24828 15384 24840
rect 15436 24828 15442 24880
rect 10376 24772 12845 24800
rect 10376 24760 10382 24772
rect 14090 24760 14096 24812
rect 14148 24800 14154 24812
rect 14441 24803 14499 24809
rect 14441 24800 14453 24803
rect 14148 24772 14453 24800
rect 14148 24760 14154 24772
rect 14441 24769 14453 24772
rect 14487 24769 14499 24803
rect 17954 24800 17960 24812
rect 17915 24772 17960 24800
rect 14441 24763 14499 24769
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 18138 24800 18144 24812
rect 18099 24772 18144 24800
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 18233 24803 18291 24809
rect 18233 24769 18245 24803
rect 18279 24769 18291 24803
rect 18233 24763 18291 24769
rect 18325 24803 18383 24809
rect 18325 24769 18337 24803
rect 18371 24800 18383 24803
rect 18984 24800 19012 24908
rect 19334 24896 19340 24908
rect 19392 24936 19398 24948
rect 23658 24936 23664 24948
rect 19392 24908 23664 24936
rect 19392 24896 19398 24908
rect 23658 24896 23664 24908
rect 23716 24936 23722 24948
rect 24397 24939 24455 24945
rect 24397 24936 24409 24939
rect 23716 24908 24409 24936
rect 23716 24896 23722 24908
rect 24397 24905 24409 24908
rect 24443 24905 24455 24939
rect 24397 24899 24455 24905
rect 37645 24939 37703 24945
rect 37645 24905 37657 24939
rect 37691 24936 37703 24939
rect 38010 24936 38016 24948
rect 37691 24908 38016 24936
rect 37691 24905 37703 24908
rect 37645 24899 37703 24905
rect 20530 24868 20536 24880
rect 19168 24840 20536 24868
rect 18371 24772 19012 24800
rect 19061 24803 19119 24809
rect 18371 24769 18383 24772
rect 18325 24763 18383 24769
rect 19061 24769 19073 24803
rect 19107 24800 19119 24803
rect 19168 24800 19196 24840
rect 20530 24828 20536 24840
rect 20588 24828 20594 24880
rect 21910 24828 21916 24880
rect 21968 24868 21974 24880
rect 21968 24840 22692 24868
rect 21968 24828 21974 24840
rect 22664 24812 22692 24840
rect 19334 24809 19340 24812
rect 19328 24800 19340 24809
rect 19107 24772 19196 24800
rect 19295 24772 19340 24800
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 19328 24763 19340 24772
rect 10778 24732 10784 24744
rect 10152 24704 10784 24732
rect 9088 24692 9094 24704
rect 10778 24692 10784 24704
rect 10836 24692 10842 24744
rect 14185 24735 14243 24741
rect 14185 24701 14197 24735
rect 14231 24701 14243 24735
rect 14185 24695 14243 24701
rect 3973 24667 4031 24673
rect 3973 24633 3985 24667
rect 4019 24664 4031 24667
rect 4062 24664 4068 24676
rect 4019 24636 4068 24664
rect 4019 24633 4031 24636
rect 3973 24627 4031 24633
rect 4062 24624 4068 24636
rect 4120 24624 4126 24676
rect 8220 24664 8248 24692
rect 13630 24664 13636 24676
rect 8220 24636 13636 24664
rect 13630 24624 13636 24636
rect 13688 24624 13694 24676
rect 14200 24608 14228 24695
rect 17770 24692 17776 24744
rect 17828 24732 17834 24744
rect 18248 24732 18276 24763
rect 19334 24760 19340 24763
rect 19392 24760 19398 24812
rect 21358 24760 21364 24812
rect 21416 24800 21422 24812
rect 22421 24803 22479 24809
rect 22421 24800 22433 24803
rect 21416 24772 22433 24800
rect 21416 24760 21422 24772
rect 22421 24769 22433 24772
rect 22467 24769 22479 24803
rect 22421 24763 22479 24769
rect 22557 24803 22615 24809
rect 22557 24769 22569 24803
rect 22603 24769 22615 24803
rect 22557 24763 22615 24769
rect 17828 24704 18276 24732
rect 17828 24692 17834 24704
rect 17402 24664 17408 24676
rect 15120 24636 17408 24664
rect 6270 24556 6276 24608
rect 6328 24596 6334 24608
rect 9030 24596 9036 24608
rect 6328 24568 9036 24596
rect 6328 24556 6334 24568
rect 9030 24556 9036 24568
rect 9088 24556 9094 24608
rect 9582 24596 9588 24608
rect 9543 24568 9588 24596
rect 9582 24556 9588 24568
rect 9640 24556 9646 24608
rect 11606 24596 11612 24608
rect 11567 24568 11612 24596
rect 11606 24556 11612 24568
rect 11664 24556 11670 24608
rect 12621 24599 12679 24605
rect 12621 24565 12633 24599
rect 12667 24596 12679 24599
rect 12894 24596 12900 24608
rect 12667 24568 12900 24596
rect 12667 24565 12679 24568
rect 12621 24559 12679 24565
rect 12894 24556 12900 24568
rect 12952 24596 12958 24608
rect 13081 24599 13139 24605
rect 13081 24596 13093 24599
rect 12952 24568 13093 24596
rect 12952 24556 12958 24568
rect 13081 24565 13093 24568
rect 13127 24565 13139 24599
rect 14182 24596 14188 24608
rect 14095 24568 14188 24596
rect 13081 24559 13139 24565
rect 14182 24556 14188 24568
rect 14240 24596 14246 24608
rect 15120 24596 15148 24636
rect 17402 24624 17408 24636
rect 17460 24624 17466 24676
rect 22572 24664 22600 24763
rect 22646 24760 22652 24812
rect 22704 24800 22710 24812
rect 22830 24800 22836 24812
rect 22704 24772 22749 24800
rect 22791 24772 22836 24800
rect 22704 24760 22710 24772
rect 22830 24760 22836 24772
rect 22888 24760 22894 24812
rect 22922 24760 22928 24812
rect 22980 24800 22986 24812
rect 22980 24772 23025 24800
rect 22980 24760 22986 24772
rect 24412 24732 24440 24899
rect 38010 24896 38016 24908
rect 38068 24896 38074 24948
rect 24670 24828 24676 24880
rect 24728 24868 24734 24880
rect 25866 24868 25872 24880
rect 24728 24840 25872 24868
rect 24728 24828 24734 24840
rect 24946 24800 24952 24812
rect 24907 24772 24952 24800
rect 24946 24760 24952 24772
rect 25004 24760 25010 24812
rect 25130 24800 25136 24812
rect 25091 24772 25136 24800
rect 25130 24760 25136 24772
rect 25188 24760 25194 24812
rect 25240 24809 25268 24840
rect 25866 24828 25872 24840
rect 25924 24828 25930 24880
rect 30466 24828 30472 24880
rect 30524 24868 30530 24880
rect 32493 24871 32551 24877
rect 30524 24840 30785 24868
rect 30524 24828 30530 24840
rect 30757 24812 30785 24840
rect 32493 24837 32505 24871
rect 32539 24868 32551 24871
rect 32766 24868 32772 24880
rect 32539 24840 32772 24868
rect 32539 24837 32551 24840
rect 32493 24831 32551 24837
rect 32766 24828 32772 24840
rect 32824 24828 32830 24880
rect 39960 24840 40264 24868
rect 25225 24803 25283 24809
rect 25225 24769 25237 24803
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 25317 24803 25375 24809
rect 25317 24769 25329 24803
rect 25363 24769 25375 24803
rect 25317 24763 25375 24769
rect 25332 24732 25360 24763
rect 26786 24760 26792 24812
rect 26844 24800 26850 24812
rect 28537 24803 28595 24809
rect 28537 24800 28549 24803
rect 26844 24772 28549 24800
rect 26844 24760 26850 24772
rect 28537 24769 28549 24772
rect 28583 24769 28595 24803
rect 28537 24763 28595 24769
rect 28804 24803 28862 24809
rect 28804 24769 28816 24803
rect 28850 24800 28862 24803
rect 29086 24800 29092 24812
rect 28850 24772 29092 24800
rect 28850 24769 28862 24772
rect 28804 24763 28862 24769
rect 29086 24760 29092 24772
rect 29144 24760 29150 24812
rect 30558 24760 30564 24812
rect 30616 24800 30622 24812
rect 30653 24803 30711 24809
rect 30653 24800 30665 24803
rect 30616 24772 30665 24800
rect 30616 24760 30622 24772
rect 30653 24769 30665 24772
rect 30699 24769 30711 24803
rect 30653 24763 30711 24769
rect 30742 24806 30800 24812
rect 30742 24772 30754 24806
rect 30788 24772 30800 24806
rect 30742 24766 30800 24772
rect 30842 24803 30900 24809
rect 30842 24769 30854 24803
rect 30888 24769 30900 24803
rect 30842 24763 30900 24769
rect 31021 24806 31079 24809
rect 31021 24803 31248 24806
rect 31021 24769 31033 24803
rect 31067 24778 31248 24803
rect 31067 24769 31079 24778
rect 31021 24763 31079 24769
rect 25590 24732 25596 24744
rect 24412 24704 25360 24732
rect 25551 24704 25596 24732
rect 25590 24692 25596 24704
rect 25648 24692 25654 24744
rect 29638 24692 29644 24744
rect 29696 24732 29702 24744
rect 30852 24732 30880 24763
rect 29696 24704 30880 24732
rect 29696 24692 29702 24704
rect 28534 24664 28540 24676
rect 22572 24636 28540 24664
rect 28534 24624 28540 24636
rect 28592 24624 28598 24676
rect 29822 24624 29828 24676
rect 29880 24664 29886 24676
rect 31220 24664 31248 24778
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32324 24732 32352 24763
rect 32582 24760 32588 24812
rect 32640 24800 32646 24812
rect 32677 24803 32735 24809
rect 32677 24800 32689 24803
rect 32640 24772 32689 24800
rect 32640 24760 32646 24772
rect 32677 24769 32689 24772
rect 32723 24769 32735 24803
rect 32677 24763 32735 24769
rect 37277 24803 37335 24809
rect 37277 24769 37289 24803
rect 37323 24800 37335 24803
rect 37366 24800 37372 24812
rect 37323 24772 37372 24800
rect 37323 24769 37335 24772
rect 37277 24763 37335 24769
rect 37366 24760 37372 24772
rect 37424 24760 37430 24812
rect 37461 24803 37519 24809
rect 37461 24769 37473 24803
rect 37507 24769 37519 24803
rect 37461 24763 37519 24769
rect 39873 24803 39931 24809
rect 39873 24769 39885 24803
rect 39919 24800 39931 24803
rect 39960 24800 39988 24840
rect 40236 24812 40264 24840
rect 39919 24772 39988 24800
rect 39919 24769 39931 24772
rect 39873 24763 39931 24769
rect 34606 24732 34612 24744
rect 32324 24704 34612 24732
rect 34606 24692 34612 24704
rect 34664 24692 34670 24744
rect 36170 24692 36176 24744
rect 36228 24732 36234 24744
rect 37476 24732 37504 24763
rect 40034 24760 40040 24812
rect 40092 24800 40098 24812
rect 40129 24803 40187 24809
rect 40129 24800 40141 24803
rect 40092 24772 40141 24800
rect 40092 24760 40098 24772
rect 40129 24769 40141 24772
rect 40175 24769 40187 24803
rect 40129 24763 40187 24769
rect 40218 24760 40224 24812
rect 40276 24760 40282 24812
rect 36228 24704 37504 24732
rect 36228 24692 36234 24704
rect 29880 24636 31248 24664
rect 29880 24624 29886 24636
rect 15562 24596 15568 24608
rect 14240 24568 15148 24596
rect 15523 24568 15568 24596
rect 14240 24556 14246 24568
rect 15562 24556 15568 24568
rect 15620 24556 15626 24608
rect 18601 24599 18659 24605
rect 18601 24565 18613 24599
rect 18647 24596 18659 24599
rect 19334 24596 19340 24608
rect 18647 24568 19340 24596
rect 18647 24565 18659 24568
rect 18601 24559 18659 24565
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 20441 24599 20499 24605
rect 20441 24565 20453 24599
rect 20487 24596 20499 24599
rect 21726 24596 21732 24608
rect 20487 24568 21732 24596
rect 20487 24565 20499 24568
rect 20441 24559 20499 24565
rect 21726 24556 21732 24568
rect 21784 24556 21790 24608
rect 22094 24556 22100 24608
rect 22152 24596 22158 24608
rect 22281 24599 22339 24605
rect 22281 24596 22293 24599
rect 22152 24568 22293 24596
rect 22152 24556 22158 24568
rect 22281 24565 22293 24568
rect 22327 24565 22339 24599
rect 22281 24559 22339 24565
rect 28902 24556 28908 24608
rect 28960 24596 28966 24608
rect 29917 24599 29975 24605
rect 29917 24596 29929 24599
rect 28960 24568 29929 24596
rect 28960 24556 28966 24568
rect 29917 24565 29929 24568
rect 29963 24565 29975 24599
rect 30374 24596 30380 24608
rect 30335 24568 30380 24596
rect 29917 24559 29975 24565
rect 30374 24556 30380 24568
rect 30432 24556 30438 24608
rect 30558 24556 30564 24608
rect 30616 24596 30622 24608
rect 31478 24596 31484 24608
rect 30616 24568 31484 24596
rect 30616 24556 30622 24568
rect 31478 24556 31484 24568
rect 31536 24556 31542 24608
rect 38746 24596 38752 24608
rect 38707 24568 38752 24596
rect 38746 24556 38752 24568
rect 38804 24556 38810 24608
rect 40865 24599 40923 24605
rect 40865 24565 40877 24599
rect 40911 24596 40923 24599
rect 41230 24596 41236 24608
rect 40911 24568 41236 24596
rect 40911 24565 40923 24568
rect 40865 24559 40923 24565
rect 41230 24556 41236 24568
rect 41288 24556 41294 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 3234 24352 3240 24404
rect 3292 24392 3298 24404
rect 3789 24395 3847 24401
rect 3789 24392 3801 24395
rect 3292 24364 3801 24392
rect 3292 24352 3298 24364
rect 3789 24361 3801 24364
rect 3835 24361 3847 24395
rect 3789 24355 3847 24361
rect 5442 24352 5448 24404
rect 5500 24392 5506 24404
rect 7926 24392 7932 24404
rect 5500 24364 7932 24392
rect 5500 24352 5506 24364
rect 7926 24352 7932 24364
rect 7984 24352 7990 24404
rect 10778 24392 10784 24404
rect 10739 24364 10784 24392
rect 10778 24352 10784 24364
rect 10836 24352 10842 24404
rect 12986 24352 12992 24404
rect 13044 24392 13050 24404
rect 14090 24392 14096 24404
rect 13044 24364 13952 24392
rect 14051 24364 14096 24392
rect 13044 24352 13050 24364
rect 13924 24324 13952 24364
rect 14090 24352 14096 24364
rect 14148 24352 14154 24404
rect 14918 24352 14924 24404
rect 14976 24392 14982 24404
rect 16117 24395 16175 24401
rect 16117 24392 16129 24395
rect 14976 24364 16129 24392
rect 14976 24352 14982 24364
rect 16117 24361 16129 24364
rect 16163 24361 16175 24395
rect 16117 24355 16175 24361
rect 18138 24352 18144 24404
rect 18196 24392 18202 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 18196 24364 19257 24392
rect 18196 24352 18202 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 19245 24355 19303 24361
rect 24673 24395 24731 24401
rect 24673 24361 24685 24395
rect 24719 24392 24731 24395
rect 25130 24392 25136 24404
rect 24719 24364 25136 24392
rect 24719 24361 24731 24364
rect 24673 24355 24731 24361
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 28902 24392 28908 24404
rect 25516 24364 28908 24392
rect 15010 24324 15016 24336
rect 13004 24296 13216 24324
rect 13924 24296 15016 24324
rect 8941 24191 8999 24197
rect 8941 24157 8953 24191
rect 8987 24188 8999 24191
rect 9674 24188 9680 24200
rect 8987 24160 9680 24188
rect 8987 24157 8999 24160
rect 8941 24151 8999 24157
rect 9674 24148 9680 24160
rect 9732 24188 9738 24200
rect 10594 24188 10600 24200
rect 9732 24160 10600 24188
rect 9732 24148 9738 24160
rect 10594 24148 10600 24160
rect 10652 24148 10658 24200
rect 11606 24148 11612 24200
rect 11664 24188 11670 24200
rect 12069 24191 12127 24197
rect 12069 24188 12081 24191
rect 11664 24160 12081 24188
rect 11664 24148 11670 24160
rect 12069 24157 12081 24160
rect 12115 24157 12127 24191
rect 12069 24151 12127 24157
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 9208 24123 9266 24129
rect 9208 24089 9220 24123
rect 9254 24120 9266 24123
rect 9582 24120 9588 24132
rect 9254 24092 9588 24120
rect 9254 24089 9266 24092
rect 9208 24083 9266 24089
rect 9582 24080 9588 24092
rect 9640 24080 9646 24132
rect 10965 24123 11023 24129
rect 10965 24089 10977 24123
rect 11011 24089 11023 24123
rect 11146 24120 11152 24132
rect 11107 24092 11152 24120
rect 10965 24083 11023 24089
rect 10226 24012 10232 24064
rect 10284 24052 10290 24064
rect 10321 24055 10379 24061
rect 10321 24052 10333 24055
rect 10284 24024 10333 24052
rect 10284 24012 10290 24024
rect 10321 24021 10333 24024
rect 10367 24052 10379 24055
rect 10980 24052 11008 24083
rect 11146 24080 11152 24092
rect 11204 24080 11210 24132
rect 11330 24080 11336 24132
rect 11388 24120 11394 24132
rect 12176 24120 12204 24151
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 12437 24191 12495 24197
rect 12308 24160 12353 24188
rect 12308 24148 12314 24160
rect 12437 24157 12449 24191
rect 12483 24188 12495 24191
rect 12894 24188 12900 24200
rect 12483 24160 12900 24188
rect 12483 24157 12495 24160
rect 12437 24151 12495 24157
rect 12894 24148 12900 24160
rect 12952 24148 12958 24200
rect 13004 24188 13032 24296
rect 13188 24256 13216 24296
rect 15010 24284 15016 24296
rect 15068 24324 15074 24336
rect 15068 24296 15332 24324
rect 15068 24284 15074 24296
rect 15197 24259 15255 24265
rect 15197 24256 15209 24259
rect 13188 24228 15209 24256
rect 15197 24225 15209 24228
rect 15243 24225 15255 24259
rect 15197 24219 15255 24225
rect 13081 24191 13139 24197
rect 13081 24188 13093 24191
rect 13004 24160 13093 24188
rect 13081 24157 13093 24160
rect 13127 24157 13139 24191
rect 13081 24151 13139 24157
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24157 13231 24191
rect 13173 24151 13231 24157
rect 13311 24191 13369 24197
rect 13311 24157 13323 24191
rect 13357 24188 13369 24191
rect 13538 24188 13544 24200
rect 13357 24160 13544 24188
rect 13357 24157 13369 24160
rect 13311 24151 13369 24157
rect 13188 24120 13216 24151
rect 13538 24148 13544 24160
rect 13596 24148 13602 24200
rect 13630 24148 13636 24200
rect 13688 24188 13694 24200
rect 14323 24191 14381 24197
rect 14323 24188 14335 24191
rect 13688 24160 14335 24188
rect 13688 24148 13694 24160
rect 14323 24157 14335 24160
rect 14369 24157 14381 24191
rect 14323 24151 14381 24157
rect 14458 24185 14516 24191
rect 14458 24151 14470 24185
rect 14504 24151 14516 24185
rect 14458 24145 14516 24151
rect 14553 24188 14611 24194
rect 14642 24188 14648 24200
rect 14553 24154 14565 24188
rect 14599 24160 14648 24188
rect 14599 24154 14611 24160
rect 14553 24148 14611 24154
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24184 14795 24191
rect 14826 24184 14832 24200
rect 14783 24157 14832 24184
rect 14737 24156 14832 24157
rect 14737 24151 14795 24156
rect 14826 24148 14832 24156
rect 14884 24148 14890 24200
rect 15304 24188 15332 24296
rect 17126 24284 17132 24336
rect 17184 24324 17190 24336
rect 18693 24327 18751 24333
rect 17184 24296 18644 24324
rect 17184 24284 17190 24296
rect 16850 24216 16856 24268
rect 16908 24256 16914 24268
rect 18616 24256 18644 24296
rect 18693 24293 18705 24327
rect 18739 24324 18751 24327
rect 18782 24324 18788 24336
rect 18739 24296 18788 24324
rect 18739 24293 18751 24296
rect 18693 24287 18751 24293
rect 18782 24284 18788 24296
rect 18840 24284 18846 24336
rect 24946 24324 24952 24336
rect 19352 24296 24952 24324
rect 19352 24256 19380 24296
rect 24946 24284 24952 24296
rect 25004 24284 25010 24336
rect 25516 24256 25544 24364
rect 28902 24352 28908 24364
rect 28960 24352 28966 24404
rect 28997 24395 29055 24401
rect 28997 24361 29009 24395
rect 29043 24392 29055 24395
rect 29638 24392 29644 24404
rect 29043 24364 29644 24392
rect 29043 24361 29055 24364
rect 28997 24355 29055 24361
rect 29638 24352 29644 24364
rect 29696 24352 29702 24404
rect 29914 24352 29920 24404
rect 29972 24392 29978 24404
rect 31110 24392 31116 24404
rect 29972 24364 31116 24392
rect 29972 24352 29978 24364
rect 31110 24352 31116 24364
rect 31168 24352 31174 24404
rect 29549 24327 29607 24333
rect 29549 24324 29561 24327
rect 16908 24228 17954 24256
rect 18616 24228 19380 24256
rect 19444 24228 21772 24256
rect 16908 24216 16914 24228
rect 15565 24191 15623 24197
rect 15565 24188 15577 24191
rect 15304 24160 15577 24188
rect 15565 24157 15577 24160
rect 15611 24157 15623 24191
rect 16298 24188 16304 24200
rect 16259 24160 16304 24188
rect 15565 24151 15623 24157
rect 16298 24148 16304 24160
rect 16356 24148 16362 24200
rect 17770 24188 17776 24200
rect 17731 24160 17776 24188
rect 17770 24148 17776 24160
rect 17828 24148 17834 24200
rect 17926 24188 17954 24228
rect 18049 24191 18107 24197
rect 18049 24188 18061 24191
rect 17926 24160 18061 24188
rect 18049 24157 18061 24160
rect 18095 24188 18107 24191
rect 18138 24188 18144 24200
rect 18095 24160 18144 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 19444 24197 19472 24228
rect 21744 24200 21772 24228
rect 22066 24228 25544 24256
rect 28966 24296 29561 24324
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24157 18567 24191
rect 18509 24151 18567 24157
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 13722 24120 13728 24132
rect 11388 24092 13728 24120
rect 11388 24080 11394 24092
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 10367 24024 11008 24052
rect 10367 24021 10379 24024
rect 10321 24015 10379 24021
rect 11238 24012 11244 24064
rect 11296 24052 11302 24064
rect 11793 24055 11851 24061
rect 11793 24052 11805 24055
rect 11296 24024 11805 24052
rect 11296 24012 11302 24024
rect 11793 24021 11805 24024
rect 11839 24021 11851 24055
rect 11793 24015 11851 24021
rect 13446 24012 13452 24064
rect 13504 24052 13510 24064
rect 13541 24055 13599 24061
rect 13541 24052 13553 24055
rect 13504 24024 13553 24052
rect 13504 24012 13510 24024
rect 13541 24021 13553 24024
rect 13587 24021 13599 24055
rect 13740 24052 13768 24080
rect 14473 24052 14501 24145
rect 14918 24080 14924 24132
rect 14976 24120 14982 24132
rect 15381 24123 15439 24129
rect 15381 24120 15393 24123
rect 14976 24092 15393 24120
rect 14976 24080 14982 24092
rect 15381 24089 15393 24092
rect 15427 24089 15439 24123
rect 15381 24083 15439 24089
rect 17126 24080 17132 24132
rect 17184 24120 17190 24132
rect 17494 24120 17500 24132
rect 17184 24092 17500 24120
rect 17184 24080 17190 24092
rect 17494 24080 17500 24092
rect 17552 24120 17558 24132
rect 18524 24120 18552 24151
rect 21358 24148 21364 24200
rect 21416 24197 21422 24200
rect 21416 24191 21465 24197
rect 21416 24157 21419 24191
rect 21453 24157 21465 24191
rect 21416 24151 21465 24157
rect 21416 24148 21422 24151
rect 21726 24148 21732 24200
rect 21784 24197 21790 24200
rect 21784 24191 21823 24197
rect 21811 24157 21823 24191
rect 21910 24188 21916 24200
rect 21871 24160 21916 24188
rect 21784 24151 21823 24157
rect 21784 24148 21790 24151
rect 21910 24148 21916 24160
rect 21968 24148 21974 24200
rect 17552 24092 18552 24120
rect 17552 24080 17558 24092
rect 18782 24080 18788 24132
rect 18840 24120 18846 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 18840 24092 19625 24120
rect 18840 24080 18846 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 19613 24083 19671 24089
rect 21545 24123 21603 24129
rect 21545 24089 21557 24123
rect 21591 24089 21603 24123
rect 21545 24083 21603 24089
rect 13740 24024 14501 24052
rect 13541 24015 13599 24021
rect 17218 24012 17224 24064
rect 17276 24052 17282 24064
rect 17770 24052 17776 24064
rect 17276 24024 17776 24052
rect 17276 24012 17282 24024
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 18230 24012 18236 24064
rect 18288 24052 18294 24064
rect 18506 24052 18512 24064
rect 18288 24024 18512 24052
rect 18288 24012 18294 24024
rect 18506 24012 18512 24024
rect 18564 24012 18570 24064
rect 21174 24012 21180 24064
rect 21232 24052 21238 24064
rect 21269 24055 21327 24061
rect 21269 24052 21281 24055
rect 21232 24024 21281 24052
rect 21232 24012 21238 24024
rect 21269 24021 21281 24024
rect 21315 24021 21327 24055
rect 21560 24052 21588 24083
rect 21634 24080 21640 24132
rect 21692 24120 21698 24132
rect 21692 24092 21737 24120
rect 21692 24080 21698 24092
rect 22066 24052 22094 24228
rect 25498 24188 25504 24200
rect 25459 24160 25504 24188
rect 25498 24148 25504 24160
rect 25556 24188 25562 24200
rect 26786 24188 26792 24200
rect 25556 24160 26792 24188
rect 25556 24148 25562 24160
rect 26786 24148 26792 24160
rect 26844 24148 26850 24200
rect 28534 24148 28540 24200
rect 28592 24188 28598 24200
rect 28813 24191 28871 24197
rect 28813 24188 28825 24191
rect 28592 24160 28825 24188
rect 28592 24148 28598 24160
rect 28813 24157 28825 24160
rect 28859 24188 28871 24191
rect 28966 24188 28994 24296
rect 29549 24293 29561 24296
rect 29595 24293 29607 24327
rect 29549 24287 29607 24293
rect 30929 24259 30987 24265
rect 30929 24225 30941 24259
rect 30975 24256 30987 24259
rect 31938 24256 31944 24268
rect 30975 24228 31944 24256
rect 30975 24225 30987 24228
rect 30929 24219 30987 24225
rect 31938 24216 31944 24228
rect 31996 24216 32002 24268
rect 28859 24160 28994 24188
rect 28859 24157 28871 24160
rect 28813 24151 28871 24157
rect 30374 24148 30380 24200
rect 30432 24188 30438 24200
rect 30662 24191 30720 24197
rect 30662 24188 30674 24191
rect 30432 24160 30674 24188
rect 30432 24148 30438 24160
rect 30662 24157 30674 24160
rect 30708 24157 30720 24191
rect 30662 24151 30720 24157
rect 38746 24148 38752 24200
rect 38804 24188 38810 24200
rect 41233 24191 41291 24197
rect 41233 24188 41245 24191
rect 38804 24160 41245 24188
rect 38804 24148 38810 24160
rect 41233 24157 41245 24160
rect 41279 24157 41291 24191
rect 58158 24188 58164 24200
rect 58119 24160 58164 24188
rect 41233 24151 41291 24157
rect 58158 24148 58164 24160
rect 58216 24148 58222 24200
rect 24857 24123 24915 24129
rect 24857 24089 24869 24123
rect 24903 24089 24915 24123
rect 24857 24083 24915 24089
rect 25041 24123 25099 24129
rect 25041 24089 25053 24123
rect 25087 24120 25099 24123
rect 25222 24120 25228 24132
rect 25087 24092 25228 24120
rect 25087 24089 25099 24092
rect 25041 24083 25099 24089
rect 21560 24024 22094 24052
rect 24872 24052 24900 24083
rect 25222 24080 25228 24092
rect 25280 24080 25286 24132
rect 25590 24080 25596 24132
rect 25648 24120 25654 24132
rect 25746 24123 25804 24129
rect 25746 24120 25758 24123
rect 25648 24092 25758 24120
rect 25648 24080 25654 24092
rect 25746 24089 25758 24092
rect 25792 24089 25804 24123
rect 28626 24120 28632 24132
rect 28587 24092 28632 24120
rect 25746 24083 25804 24089
rect 28626 24080 28632 24092
rect 28684 24080 28690 24132
rect 40126 24080 40132 24132
rect 40184 24120 40190 24132
rect 40221 24123 40279 24129
rect 40221 24120 40233 24123
rect 40184 24092 40233 24120
rect 40184 24080 40190 24092
rect 40221 24089 40233 24092
rect 40267 24089 40279 24123
rect 40402 24120 40408 24132
rect 40363 24092 40408 24120
rect 40221 24083 40279 24089
rect 26878 24052 26884 24064
rect 24872 24024 26884 24052
rect 21269 24015 21327 24021
rect 26878 24012 26884 24024
rect 26936 24012 26942 24064
rect 27246 24012 27252 24064
rect 27304 24052 27310 24064
rect 32306 24052 32312 24064
rect 27304 24024 32312 24052
rect 27304 24012 27310 24024
rect 32306 24012 32312 24024
rect 32364 24012 32370 24064
rect 40236 24052 40264 24083
rect 40402 24080 40408 24092
rect 40460 24080 40466 24132
rect 41049 24123 41107 24129
rect 41049 24120 41061 24123
rect 40512 24092 41061 24120
rect 40512 24052 40540 24092
rect 41049 24089 41061 24092
rect 41095 24089 41107 24123
rect 41049 24083 41107 24089
rect 40236 24024 40540 24052
rect 40589 24055 40647 24061
rect 40589 24021 40601 24055
rect 40635 24052 40647 24055
rect 40954 24052 40960 24064
rect 40635 24024 40960 24052
rect 40635 24021 40647 24024
rect 40589 24015 40647 24021
rect 40954 24012 40960 24024
rect 41012 24012 41018 24064
rect 41414 24052 41420 24064
rect 41375 24024 41420 24052
rect 41414 24012 41420 24024
rect 41472 24012 41478 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 5258 23808 5264 23860
rect 5316 23848 5322 23860
rect 8570 23848 8576 23860
rect 5316 23820 8576 23848
rect 5316 23808 5322 23820
rect 8570 23808 8576 23820
rect 8628 23848 8634 23860
rect 8941 23851 8999 23857
rect 8941 23848 8953 23851
rect 8628 23820 8953 23848
rect 8628 23808 8634 23820
rect 8941 23817 8953 23820
rect 8987 23817 8999 23851
rect 9950 23848 9956 23860
rect 9863 23820 9956 23848
rect 8941 23811 8999 23817
rect 2222 23712 2228 23724
rect 2183 23684 2228 23712
rect 2222 23672 2228 23684
rect 2280 23672 2286 23724
rect 2409 23715 2467 23721
rect 2409 23681 2421 23715
rect 2455 23712 2467 23715
rect 3234 23712 3240 23724
rect 2455 23684 3240 23712
rect 2455 23681 2467 23684
rect 2409 23675 2467 23681
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 8956 23712 8984 23811
rect 9582 23712 9588 23724
rect 8956 23684 9588 23712
rect 9582 23672 9588 23684
rect 9640 23712 9646 23724
rect 9876 23721 9904 23820
rect 9950 23808 9956 23820
rect 10008 23848 10014 23860
rect 11330 23848 11336 23860
rect 10008 23820 11336 23848
rect 10008 23808 10014 23820
rect 11330 23808 11336 23820
rect 11388 23808 11394 23860
rect 12069 23851 12127 23857
rect 12069 23817 12081 23851
rect 12115 23848 12127 23851
rect 12250 23848 12256 23860
rect 12115 23820 12256 23848
rect 12115 23817 12127 23820
rect 12069 23811 12127 23817
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12434 23808 12440 23860
rect 12492 23848 12498 23860
rect 21542 23848 21548 23860
rect 12492 23820 14320 23848
rect 12492 23808 12498 23820
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 11146 23780 11152 23792
rect 11011 23752 11152 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 11146 23740 11152 23752
rect 11204 23780 11210 23792
rect 11701 23783 11759 23789
rect 11701 23780 11713 23783
rect 11204 23752 11713 23780
rect 11204 23740 11210 23752
rect 11701 23749 11713 23752
rect 11747 23780 11759 23783
rect 12986 23780 12992 23792
rect 11747 23752 12992 23780
rect 11747 23749 11759 23752
rect 11701 23743 11759 23749
rect 12986 23740 12992 23752
rect 13044 23740 13050 23792
rect 14182 23780 14188 23792
rect 13188 23752 14188 23780
rect 9769 23715 9827 23721
rect 9769 23712 9781 23715
rect 9640 23684 9781 23712
rect 9640 23672 9646 23684
rect 9769 23681 9781 23684
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 9861 23715 9919 23721
rect 9861 23681 9873 23715
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23681 10011 23715
rect 9953 23675 10011 23681
rect 10137 23715 10195 23721
rect 10137 23681 10149 23715
rect 10183 23712 10195 23715
rect 10318 23712 10324 23724
rect 10183 23684 10324 23712
rect 10183 23681 10195 23684
rect 10137 23675 10195 23681
rect 6086 23604 6092 23656
rect 6144 23644 6150 23656
rect 7377 23647 7435 23653
rect 7377 23644 7389 23647
rect 6144 23616 7389 23644
rect 6144 23604 6150 23616
rect 7377 23613 7389 23616
rect 7423 23613 7435 23647
rect 7377 23607 7435 23613
rect 7653 23647 7711 23653
rect 7653 23613 7665 23647
rect 7699 23613 7711 23647
rect 9968 23644 9996 23675
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 10778 23712 10784 23724
rect 10739 23684 10784 23712
rect 10778 23672 10784 23684
rect 10836 23672 10842 23724
rect 13188 23721 13216 23752
rect 14182 23740 14188 23752
rect 14240 23740 14246 23792
rect 14292 23780 14320 23820
rect 14752 23820 21548 23848
rect 14752 23780 14780 23820
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22186 23808 22192 23860
rect 22244 23848 22250 23860
rect 24397 23851 24455 23857
rect 24397 23848 24409 23851
rect 22244 23820 24409 23848
rect 22244 23808 22250 23820
rect 24397 23817 24409 23820
rect 24443 23848 24455 23851
rect 24762 23848 24768 23860
rect 24443 23820 24768 23848
rect 24443 23817 24455 23820
rect 24397 23811 24455 23817
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 24946 23848 24952 23860
rect 24907 23820 24952 23848
rect 24946 23808 24952 23820
rect 25004 23848 25010 23860
rect 29086 23848 29092 23860
rect 25004 23820 25973 23848
rect 29047 23820 29092 23848
rect 25004 23808 25010 23820
rect 14292 23752 14780 23780
rect 17037 23783 17095 23789
rect 17037 23749 17049 23783
rect 17083 23780 17095 23783
rect 17126 23780 17132 23792
rect 17083 23752 17132 23780
rect 17083 23749 17095 23752
rect 17037 23743 17095 23749
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 17405 23783 17463 23789
rect 17405 23749 17417 23783
rect 17451 23780 17463 23783
rect 22646 23780 22652 23792
rect 17451 23752 18000 23780
rect 22607 23752 22652 23780
rect 17451 23749 17463 23752
rect 17405 23743 17463 23749
rect 13446 23721 13452 23724
rect 11885 23715 11943 23721
rect 11885 23712 11897 23715
rect 11716 23684 11897 23712
rect 11716 23656 11744 23684
rect 11885 23681 11897 23684
rect 11931 23681 11943 23715
rect 11885 23675 11943 23681
rect 13173 23715 13231 23721
rect 13173 23681 13185 23715
rect 13219 23681 13231 23715
rect 13440 23712 13452 23721
rect 13407 23684 13452 23712
rect 13173 23675 13231 23681
rect 13440 23675 13452 23684
rect 13446 23672 13452 23675
rect 13504 23672 13510 23724
rect 17218 23712 17224 23724
rect 17179 23684 17224 23712
rect 17218 23672 17224 23684
rect 17276 23672 17282 23724
rect 17770 23672 17776 23724
rect 17828 23712 17834 23724
rect 17865 23715 17923 23721
rect 17865 23712 17877 23715
rect 17828 23684 17877 23712
rect 17828 23672 17834 23684
rect 17865 23681 17877 23684
rect 17911 23681 17923 23715
rect 17972 23712 18000 23752
rect 22646 23740 22652 23752
rect 22704 23740 22710 23792
rect 22741 23783 22799 23789
rect 22741 23749 22753 23783
rect 22787 23780 22799 23783
rect 25314 23780 25320 23792
rect 22787 23752 25320 23780
rect 22787 23749 22799 23752
rect 22741 23743 22799 23749
rect 25314 23740 25320 23752
rect 25372 23740 25378 23792
rect 18028 23715 18086 23721
rect 18028 23712 18040 23715
rect 17972 23684 18040 23712
rect 17865 23675 17923 23681
rect 18028 23681 18040 23684
rect 18074 23681 18086 23715
rect 18028 23675 18086 23681
rect 18128 23715 18186 23721
rect 18128 23681 18140 23715
rect 18174 23712 18186 23715
rect 18174 23681 18187 23712
rect 18128 23675 18187 23681
rect 10597 23647 10655 23653
rect 10597 23644 10609 23647
rect 9968 23616 10609 23644
rect 7653 23607 7711 23613
rect 10597 23613 10609 23616
rect 10643 23613 10655 23647
rect 10597 23607 10655 23613
rect 7668 23576 7696 23607
rect 11698 23604 11704 23656
rect 11756 23604 11762 23656
rect 14826 23604 14832 23656
rect 14884 23644 14890 23656
rect 14884 23616 15148 23644
rect 14884 23604 14890 23616
rect 8205 23579 8263 23585
rect 8205 23576 8217 23579
rect 7668 23548 8217 23576
rect 8205 23545 8217 23548
rect 8251 23576 8263 23579
rect 11790 23576 11796 23588
rect 8251 23548 11796 23576
rect 8251 23545 8263 23548
rect 8205 23539 8263 23545
rect 11790 23536 11796 23548
rect 11848 23536 11854 23588
rect 14458 23536 14464 23588
rect 14516 23576 14522 23588
rect 14553 23579 14611 23585
rect 14553 23576 14565 23579
rect 14516 23548 14565 23576
rect 14516 23536 14522 23548
rect 14553 23545 14565 23548
rect 14599 23576 14611 23579
rect 14918 23576 14924 23588
rect 14599 23548 14924 23576
rect 14599 23545 14611 23548
rect 14553 23539 14611 23545
rect 14918 23536 14924 23548
rect 14976 23536 14982 23588
rect 15120 23585 15148 23616
rect 18159 23588 18187 23675
rect 18230 23672 18236 23724
rect 18288 23721 18294 23724
rect 18288 23715 18311 23721
rect 18299 23681 18311 23715
rect 22370 23712 22376 23724
rect 22331 23684 22376 23712
rect 18288 23675 18311 23681
rect 18288 23672 18294 23675
rect 22370 23672 22376 23684
rect 22428 23672 22434 23724
rect 22554 23721 22560 23724
rect 22521 23715 22560 23721
rect 22521 23681 22533 23715
rect 22521 23675 22560 23681
rect 22554 23672 22560 23675
rect 22612 23672 22618 23724
rect 22838 23715 22896 23721
rect 22838 23681 22850 23715
rect 22884 23681 22896 23715
rect 22838 23675 22896 23681
rect 18506 23604 18512 23656
rect 18564 23644 18570 23656
rect 19334 23644 19340 23656
rect 18564 23616 19340 23644
rect 18564 23604 18570 23616
rect 19334 23604 19340 23616
rect 19392 23604 19398 23656
rect 21358 23604 21364 23656
rect 21416 23644 21422 23656
rect 22853 23644 22881 23675
rect 24946 23672 24952 23724
rect 25004 23712 25010 23724
rect 25501 23715 25559 23721
rect 25501 23712 25513 23715
rect 25004 23684 25513 23712
rect 25004 23672 25010 23684
rect 25501 23681 25513 23684
rect 25547 23681 25559 23715
rect 25682 23712 25688 23724
rect 25643 23684 25688 23712
rect 25501 23675 25559 23681
rect 25682 23672 25688 23684
rect 25740 23672 25746 23724
rect 25945 23721 25973 23820
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 30834 23808 30840 23860
rect 30892 23848 30898 23860
rect 33962 23848 33968 23860
rect 30892 23820 33968 23848
rect 30892 23808 30898 23820
rect 33962 23808 33968 23820
rect 34020 23808 34026 23860
rect 41230 23848 41236 23860
rect 40880 23820 41236 23848
rect 31570 23740 31576 23792
rect 31628 23780 31634 23792
rect 32950 23780 32956 23792
rect 31628 23752 32812 23780
rect 32911 23752 32956 23780
rect 31628 23740 31634 23752
rect 25780 23715 25838 23721
rect 25780 23681 25792 23715
rect 25826 23681 25838 23715
rect 25780 23675 25838 23681
rect 25889 23715 25973 23721
rect 25889 23681 25901 23715
rect 25935 23684 25973 23715
rect 25935 23681 25947 23684
rect 25889 23675 25947 23681
rect 21416 23616 22881 23644
rect 21416 23604 21422 23616
rect 24670 23604 24676 23656
rect 24728 23644 24734 23656
rect 25792 23644 25820 23675
rect 28810 23672 28816 23724
rect 28868 23712 28874 23724
rect 29319 23715 29377 23721
rect 29319 23712 29331 23715
rect 28868 23684 29331 23712
rect 28868 23672 28874 23684
rect 29319 23681 29331 23684
rect 29365 23681 29377 23715
rect 29319 23675 29377 23681
rect 29457 23715 29515 23721
rect 29457 23681 29469 23715
rect 29503 23681 29515 23715
rect 29457 23675 29515 23681
rect 24728 23616 25820 23644
rect 24728 23604 24734 23616
rect 28258 23604 28264 23656
rect 28316 23644 28322 23656
rect 29472 23644 29500 23675
rect 29546 23672 29552 23724
rect 29604 23721 29610 23724
rect 32784 23721 32812 23752
rect 32950 23740 32956 23752
rect 33008 23740 33014 23792
rect 33318 23740 33324 23792
rect 33376 23780 33382 23792
rect 33413 23783 33471 23789
rect 33413 23780 33425 23783
rect 33376 23752 33425 23780
rect 33376 23740 33382 23752
rect 33413 23749 33425 23752
rect 33459 23749 33471 23783
rect 33413 23743 33471 23749
rect 35897 23783 35955 23789
rect 35897 23749 35909 23783
rect 35943 23780 35955 23783
rect 36078 23780 36084 23792
rect 35943 23752 36084 23780
rect 35943 23749 35955 23752
rect 35897 23743 35955 23749
rect 36078 23740 36084 23752
rect 36136 23740 36142 23792
rect 39884 23783 39942 23789
rect 39884 23749 39896 23783
rect 39930 23780 39942 23783
rect 40589 23783 40647 23789
rect 40589 23780 40601 23783
rect 39930 23752 40601 23780
rect 39930 23749 39942 23752
rect 39884 23743 39942 23749
rect 40589 23749 40601 23752
rect 40635 23749 40647 23783
rect 40880 23780 40908 23820
rect 41230 23808 41236 23820
rect 41288 23848 41294 23860
rect 41693 23851 41751 23857
rect 41693 23848 41705 23851
rect 41288 23820 41705 23848
rect 41288 23808 41294 23820
rect 41693 23817 41705 23820
rect 41739 23817 41751 23851
rect 41693 23811 41751 23817
rect 40589 23743 40647 23749
rect 40860 23752 40908 23780
rect 29604 23712 29612 23721
rect 29733 23715 29791 23721
rect 29604 23684 29649 23712
rect 29604 23675 29612 23684
rect 29733 23681 29745 23715
rect 29779 23681 29791 23715
rect 29733 23675 29791 23681
rect 32677 23715 32735 23721
rect 32677 23681 32689 23715
rect 32723 23681 32735 23715
rect 32677 23675 32735 23681
rect 32769 23715 32827 23721
rect 32769 23681 32781 23715
rect 32815 23681 32827 23715
rect 32769 23675 32827 23681
rect 33689 23715 33747 23721
rect 33689 23681 33701 23715
rect 33735 23712 33747 23715
rect 35618 23712 35624 23724
rect 33735 23684 35624 23712
rect 33735 23681 33747 23684
rect 33689 23675 33747 23681
rect 29604 23672 29610 23675
rect 29748 23644 29776 23675
rect 29822 23644 29828 23656
rect 28316 23616 29500 23644
rect 29735 23616 29828 23644
rect 28316 23604 28322 23616
rect 15105 23579 15163 23585
rect 15105 23545 15117 23579
rect 15151 23576 15163 23579
rect 15151 23548 16436 23576
rect 15151 23545 15163 23548
rect 15105 23539 15163 23545
rect 2498 23468 2504 23520
rect 2556 23508 2562 23520
rect 2593 23511 2651 23517
rect 2593 23508 2605 23511
rect 2556 23480 2605 23508
rect 2556 23468 2562 23480
rect 2593 23477 2605 23480
rect 2639 23477 2651 23511
rect 9490 23508 9496 23520
rect 9451 23480 9496 23508
rect 2593 23471 2651 23477
rect 9490 23468 9496 23480
rect 9548 23468 9554 23520
rect 9582 23468 9588 23520
rect 9640 23508 9646 23520
rect 12434 23508 12440 23520
rect 9640 23480 12440 23508
rect 9640 23468 9646 23480
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 12526 23468 12532 23520
rect 12584 23508 12590 23520
rect 12621 23511 12679 23517
rect 12621 23508 12633 23511
rect 12584 23480 12633 23508
rect 12584 23468 12590 23480
rect 12621 23477 12633 23480
rect 12667 23508 12679 23511
rect 13538 23508 13544 23520
rect 12667 23480 13544 23508
rect 12667 23477 12679 23480
rect 12621 23471 12679 23477
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 15378 23468 15384 23520
rect 15436 23508 15442 23520
rect 15841 23511 15899 23517
rect 15841 23508 15853 23511
rect 15436 23480 15853 23508
rect 15436 23468 15442 23480
rect 15841 23477 15853 23480
rect 15887 23508 15899 23511
rect 16298 23508 16304 23520
rect 15887 23480 16304 23508
rect 15887 23477 15899 23480
rect 15841 23471 15899 23477
rect 16298 23468 16304 23480
rect 16356 23468 16362 23520
rect 16408 23508 16436 23548
rect 18138 23536 18144 23588
rect 18196 23536 18202 23588
rect 21450 23576 21456 23588
rect 18239 23548 21456 23576
rect 18239 23508 18267 23548
rect 21450 23536 21456 23548
rect 21508 23536 21514 23588
rect 18506 23508 18512 23520
rect 16408 23480 18267 23508
rect 18467 23480 18512 23508
rect 18506 23468 18512 23480
rect 18564 23468 18570 23520
rect 23017 23511 23075 23517
rect 23017 23477 23029 23511
rect 23063 23508 23075 23511
rect 23198 23508 23204 23520
rect 23063 23480 23204 23508
rect 23063 23477 23075 23480
rect 23017 23471 23075 23477
rect 23198 23468 23204 23480
rect 23256 23468 23262 23520
rect 26142 23508 26148 23520
rect 26103 23480 26148 23508
rect 26142 23468 26148 23480
rect 26200 23468 26206 23520
rect 28629 23511 28687 23517
rect 28629 23477 28641 23511
rect 28675 23508 28687 23511
rect 28810 23508 28816 23520
rect 28675 23480 28816 23508
rect 28675 23477 28687 23480
rect 28629 23471 28687 23477
rect 28810 23468 28816 23480
rect 28868 23468 28874 23520
rect 29380 23508 29408 23616
rect 29454 23536 29460 23588
rect 29512 23576 29518 23588
rect 29748 23576 29776 23616
rect 29822 23604 29828 23616
rect 29880 23644 29886 23656
rect 30193 23647 30251 23653
rect 30193 23644 30205 23647
rect 29880 23616 30205 23644
rect 29880 23604 29886 23616
rect 30193 23613 30205 23616
rect 30239 23613 30251 23647
rect 30193 23607 30251 23613
rect 29512 23548 29776 23576
rect 32692 23576 32720 23675
rect 35618 23672 35624 23684
rect 35676 23672 35682 23724
rect 35802 23712 35808 23724
rect 35763 23684 35808 23712
rect 35802 23672 35808 23684
rect 35860 23672 35866 23724
rect 35986 23712 35992 23724
rect 35947 23684 35992 23712
rect 35986 23672 35992 23684
rect 36044 23672 36050 23724
rect 36170 23712 36176 23724
rect 36131 23684 36176 23712
rect 36170 23672 36176 23684
rect 36228 23672 36234 23724
rect 40034 23672 40040 23724
rect 40092 23712 40098 23724
rect 40860 23721 40888 23752
rect 40129 23715 40187 23721
rect 40129 23712 40141 23715
rect 40092 23684 40141 23712
rect 40092 23672 40098 23684
rect 40129 23681 40141 23684
rect 40175 23681 40187 23715
rect 40129 23675 40187 23681
rect 40845 23715 40903 23721
rect 40845 23681 40857 23715
rect 40891 23681 40903 23715
rect 40845 23675 40903 23681
rect 40957 23715 41015 23721
rect 40957 23681 40969 23715
rect 41003 23681 41015 23715
rect 40957 23675 41015 23681
rect 33597 23647 33655 23653
rect 33597 23613 33609 23647
rect 33643 23644 33655 23647
rect 34238 23644 34244 23656
rect 33643 23616 34244 23644
rect 33643 23613 33655 23616
rect 33597 23607 33655 23613
rect 34238 23604 34244 23616
rect 34296 23604 34302 23656
rect 37918 23644 37924 23656
rect 37879 23616 37924 23644
rect 37918 23604 37924 23616
rect 37976 23604 37982 23656
rect 40972 23588 41000 23675
rect 41046 23672 41052 23724
rect 41104 23721 41110 23724
rect 41104 23712 41112 23721
rect 41233 23715 41291 23721
rect 41104 23684 41149 23712
rect 41104 23675 41112 23684
rect 41233 23681 41245 23715
rect 41279 23681 41291 23715
rect 41233 23675 41291 23681
rect 41104 23672 41110 23675
rect 41248 23644 41276 23675
rect 41064 23616 41276 23644
rect 41064 23588 41092 23616
rect 35621 23579 35679 23585
rect 35621 23576 35633 23579
rect 32692 23548 35633 23576
rect 29512 23536 29518 23548
rect 35621 23545 35633 23548
rect 35667 23545 35679 23579
rect 35621 23539 35679 23545
rect 37461 23579 37519 23585
rect 37461 23545 37473 23579
rect 37507 23576 37519 23579
rect 38378 23576 38384 23588
rect 37507 23548 38384 23576
rect 37507 23545 37519 23548
rect 37461 23539 37519 23545
rect 38378 23536 38384 23548
rect 38436 23536 38442 23588
rect 40954 23536 40960 23588
rect 41012 23536 41018 23588
rect 41046 23536 41052 23588
rect 41104 23536 41110 23588
rect 30466 23508 30472 23520
rect 29380 23480 30472 23508
rect 30466 23468 30472 23480
rect 30524 23468 30530 23520
rect 32490 23508 32496 23520
rect 32451 23480 32496 23508
rect 32490 23468 32496 23480
rect 32548 23468 32554 23520
rect 32674 23508 32680 23520
rect 32635 23480 32680 23508
rect 32674 23468 32680 23480
rect 32732 23468 32738 23520
rect 32766 23468 32772 23520
rect 32824 23508 32830 23520
rect 33413 23511 33471 23517
rect 33413 23508 33425 23511
rect 32824 23480 33425 23508
rect 32824 23468 32830 23480
rect 33413 23477 33425 23480
rect 33459 23477 33471 23511
rect 33413 23471 33471 23477
rect 33502 23468 33508 23520
rect 33560 23508 33566 23520
rect 33873 23511 33931 23517
rect 33873 23508 33885 23511
rect 33560 23480 33885 23508
rect 33560 23468 33566 23480
rect 33873 23477 33885 23480
rect 33919 23477 33931 23511
rect 33873 23471 33931 23477
rect 35894 23468 35900 23520
rect 35952 23508 35958 23520
rect 38749 23511 38807 23517
rect 38749 23508 38761 23511
rect 35952 23480 38761 23508
rect 35952 23468 35958 23480
rect 38749 23477 38761 23480
rect 38795 23508 38807 23511
rect 40402 23508 40408 23520
rect 38795 23480 40408 23508
rect 38795 23477 38807 23480
rect 38749 23471 38807 23477
rect 40402 23468 40408 23480
rect 40460 23468 40466 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 2958 23264 2964 23316
rect 3016 23304 3022 23316
rect 3789 23307 3847 23313
rect 3789 23304 3801 23307
rect 3016 23276 3801 23304
rect 3016 23264 3022 23276
rect 3789 23273 3801 23276
rect 3835 23304 3847 23307
rect 3970 23304 3976 23316
rect 3835 23276 3976 23304
rect 3835 23273 3847 23276
rect 3789 23267 3847 23273
rect 3970 23264 3976 23276
rect 4028 23264 4034 23316
rect 18230 23304 18236 23316
rect 18191 23276 18236 23304
rect 18230 23264 18236 23276
rect 18288 23264 18294 23316
rect 23106 23264 23112 23316
rect 23164 23304 23170 23316
rect 23201 23307 23259 23313
rect 23201 23304 23213 23307
rect 23164 23276 23213 23304
rect 23164 23264 23170 23276
rect 23201 23273 23213 23276
rect 23247 23273 23259 23307
rect 29546 23304 29552 23316
rect 23201 23267 23259 23273
rect 23308 23276 29552 23304
rect 2976 23168 3004 23264
rect 2424 23140 3004 23168
rect 12406 23140 16068 23168
rect 2424 23100 2452 23140
rect 2547 23103 2605 23109
rect 2547 23100 2559 23103
rect 2424 23072 2559 23100
rect 2547 23069 2559 23072
rect 2593 23069 2605 23103
rect 2682 23100 2688 23112
rect 2643 23072 2688 23100
rect 2547 23063 2605 23069
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 2774 23060 2780 23112
rect 2832 23100 2838 23112
rect 2832 23072 2877 23100
rect 2832 23060 2838 23072
rect 2958 23060 2964 23112
rect 3016 23100 3022 23112
rect 7374 23100 7380 23112
rect 3016 23072 3061 23100
rect 7335 23072 7380 23100
rect 3016 23060 3022 23072
rect 7374 23060 7380 23072
rect 7432 23060 7438 23112
rect 7653 23103 7711 23109
rect 7653 23069 7665 23103
rect 7699 23100 7711 23103
rect 8941 23103 8999 23109
rect 7699 23072 8248 23100
rect 7699 23069 7711 23072
rect 7653 23063 7711 23069
rect 2222 22992 2228 23044
rect 2280 23032 2286 23044
rect 4614 23032 4620 23044
rect 2280 23004 4620 23032
rect 2280 22992 2286 23004
rect 4614 22992 4620 23004
rect 4672 23032 4678 23044
rect 4672 23004 7696 23032
rect 4672 22992 4678 23004
rect 7668 22976 7696 23004
rect 2317 22967 2375 22973
rect 2317 22933 2329 22967
rect 2363 22964 2375 22967
rect 2682 22964 2688 22976
rect 2363 22936 2688 22964
rect 2363 22933 2375 22936
rect 2317 22927 2375 22933
rect 2682 22924 2688 22936
rect 2740 22924 2746 22976
rect 7650 22924 7656 22976
rect 7708 22924 7714 22976
rect 8220 22973 8248 23072
rect 8941 23069 8953 23103
rect 8987 23100 8999 23103
rect 9674 23100 9680 23112
rect 8987 23072 9680 23100
rect 8987 23069 8999 23072
rect 8941 23063 8999 23069
rect 9674 23060 9680 23072
rect 9732 23100 9738 23112
rect 11238 23109 11244 23112
rect 10965 23103 11023 23109
rect 10965 23100 10977 23103
rect 9732 23072 10977 23100
rect 9732 23060 9738 23072
rect 10965 23069 10977 23072
rect 11011 23069 11023 23103
rect 11232 23100 11244 23109
rect 11199 23072 11244 23100
rect 10965 23063 11023 23069
rect 11232 23063 11244 23072
rect 11238 23060 11244 23063
rect 11296 23060 11302 23112
rect 11514 23060 11520 23112
rect 11572 23100 11578 23112
rect 12406 23100 12434 23140
rect 14826 23100 14832 23112
rect 11572 23072 12434 23100
rect 14787 23072 14832 23100
rect 11572 23060 11578 23072
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 15197 23103 15255 23109
rect 15197 23100 15209 23103
rect 14936 23072 15209 23100
rect 9208 23035 9266 23041
rect 9208 23001 9220 23035
rect 9254 23032 9266 23035
rect 9490 23032 9496 23044
rect 9254 23004 9496 23032
rect 9254 23001 9266 23004
rect 9208 22995 9266 23001
rect 9490 22992 9496 23004
rect 9548 22992 9554 23044
rect 11882 23032 11888 23044
rect 10060 23004 11888 23032
rect 8205 22967 8263 22973
rect 8205 22933 8217 22967
rect 8251 22964 8263 22967
rect 10060 22964 10088 23004
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 14366 23032 14372 23044
rect 14279 23004 14372 23032
rect 14366 22992 14372 23004
rect 14424 23032 14430 23044
rect 14936 23032 14964 23072
rect 15197 23069 15209 23072
rect 15243 23100 15255 23103
rect 15243 23072 15884 23100
rect 15243 23069 15255 23072
rect 15197 23063 15255 23069
rect 14424 23004 14964 23032
rect 15013 23035 15071 23041
rect 14424 22992 14430 23004
rect 15013 23001 15025 23035
rect 15059 23001 15071 23035
rect 15013 22995 15071 23001
rect 15105 23035 15163 23041
rect 15105 23001 15117 23035
rect 15151 23032 15163 23035
rect 15562 23032 15568 23044
rect 15151 23004 15568 23032
rect 15151 23001 15163 23004
rect 15105 22995 15163 23001
rect 8251 22936 10088 22964
rect 8251 22933 8263 22936
rect 8205 22927 8263 22933
rect 10134 22924 10140 22976
rect 10192 22964 10198 22976
rect 10321 22967 10379 22973
rect 10321 22964 10333 22967
rect 10192 22936 10333 22964
rect 10192 22924 10198 22936
rect 10321 22933 10333 22936
rect 10367 22964 10379 22967
rect 10778 22964 10784 22976
rect 10367 22936 10784 22964
rect 10367 22933 10379 22936
rect 10321 22927 10379 22933
rect 10778 22924 10784 22936
rect 10836 22924 10842 22976
rect 11698 22924 11704 22976
rect 11756 22964 11762 22976
rect 12345 22967 12403 22973
rect 12345 22964 12357 22967
rect 11756 22936 12357 22964
rect 11756 22924 11762 22936
rect 12345 22933 12357 22936
rect 12391 22933 12403 22967
rect 12345 22927 12403 22933
rect 14918 22924 14924 22976
rect 14976 22964 14982 22976
rect 15028 22964 15056 22995
rect 15562 22992 15568 23004
rect 15620 22992 15626 23044
rect 15856 23032 15884 23072
rect 15930 23060 15936 23112
rect 15988 23100 15994 23112
rect 16040 23109 16068 23140
rect 17586 23128 17592 23180
rect 17644 23168 17650 23180
rect 23106 23168 23112 23180
rect 17644 23140 23112 23168
rect 17644 23128 17650 23140
rect 23106 23128 23112 23140
rect 23164 23128 23170 23180
rect 16025 23103 16083 23109
rect 16025 23100 16037 23103
rect 15988 23072 16037 23100
rect 15988 23060 15994 23072
rect 16025 23069 16037 23072
rect 16071 23069 16083 23103
rect 22738 23100 22744 23112
rect 16025 23063 16083 23069
rect 16132 23072 22744 23100
rect 16132 23032 16160 23072
rect 22738 23060 22744 23072
rect 22796 23060 22802 23112
rect 23198 23100 23204 23112
rect 23159 23072 23204 23100
rect 23198 23060 23204 23072
rect 23256 23060 23262 23112
rect 23308 23109 23336 23276
rect 29546 23264 29552 23276
rect 29604 23264 29610 23316
rect 39114 23304 39120 23316
rect 36280 23276 39120 23304
rect 35897 23239 35955 23245
rect 35897 23205 35909 23239
rect 35943 23236 35955 23239
rect 36078 23236 36084 23248
rect 35943 23208 36084 23236
rect 35943 23205 35955 23208
rect 35897 23199 35955 23205
rect 36078 23196 36084 23208
rect 36136 23196 36142 23248
rect 25498 23128 25504 23180
rect 25556 23168 25562 23180
rect 25869 23171 25927 23177
rect 25869 23168 25881 23171
rect 25556 23140 25881 23168
rect 25556 23128 25562 23140
rect 25869 23137 25881 23140
rect 25915 23137 25927 23171
rect 34146 23168 34152 23180
rect 34107 23140 34152 23168
rect 25869 23131 25927 23137
rect 34146 23128 34152 23140
rect 34204 23128 34210 23180
rect 35802 23168 35808 23180
rect 35084 23140 35808 23168
rect 23293 23103 23351 23109
rect 23293 23069 23305 23103
rect 23339 23069 23351 23103
rect 23293 23063 23351 23069
rect 23382 23060 23388 23112
rect 23440 23100 23446 23112
rect 24397 23103 24455 23109
rect 24397 23100 24409 23103
rect 23440 23072 24409 23100
rect 23440 23060 23446 23072
rect 24397 23069 24409 23072
rect 24443 23069 24455 23103
rect 24670 23100 24676 23112
rect 24631 23072 24676 23100
rect 24397 23063 24455 23069
rect 24670 23060 24676 23072
rect 24728 23060 24734 23112
rect 26142 23109 26148 23112
rect 26136 23100 26148 23109
rect 26103 23072 26148 23100
rect 26136 23063 26148 23072
rect 26142 23060 26148 23063
rect 26200 23060 26206 23112
rect 35084 23109 35112 23140
rect 35802 23128 35808 23140
rect 35860 23128 35866 23180
rect 35069 23103 35127 23109
rect 35069 23069 35081 23103
rect 35115 23069 35127 23103
rect 35069 23063 35127 23069
rect 35437 23103 35495 23109
rect 35437 23069 35449 23103
rect 35483 23100 35495 23103
rect 36280 23100 36308 23276
rect 39114 23264 39120 23276
rect 39172 23264 39178 23316
rect 40129 23307 40187 23313
rect 40129 23273 40141 23307
rect 40175 23304 40187 23307
rect 40218 23304 40224 23316
rect 40175 23276 40224 23304
rect 40175 23273 40187 23276
rect 40129 23267 40187 23273
rect 40218 23264 40224 23276
rect 40276 23264 40282 23316
rect 41414 23168 41420 23180
rect 38120 23140 40540 23168
rect 35483 23072 36308 23100
rect 35483 23069 35495 23072
rect 35437 23063 35495 23069
rect 37182 23060 37188 23112
rect 37240 23100 37246 23112
rect 37277 23103 37335 23109
rect 37277 23100 37289 23103
rect 37240 23072 37289 23100
rect 37240 23060 37246 23072
rect 37277 23069 37289 23072
rect 37323 23069 37335 23103
rect 37277 23063 37335 23069
rect 37918 23060 37924 23112
rect 37976 23100 37982 23112
rect 38120 23109 38148 23140
rect 38013 23103 38071 23109
rect 38013 23100 38025 23103
rect 37976 23072 38025 23100
rect 37976 23060 37982 23072
rect 38013 23069 38025 23072
rect 38059 23069 38071 23103
rect 38013 23063 38071 23069
rect 38105 23103 38163 23109
rect 38105 23069 38117 23103
rect 38151 23069 38163 23103
rect 38105 23063 38163 23069
rect 38194 23060 38200 23112
rect 38252 23100 38258 23112
rect 38252 23072 38297 23100
rect 38252 23060 38258 23072
rect 38378 23060 38384 23112
rect 38436 23100 38442 23112
rect 40402 23109 40408 23112
rect 40385 23103 40408 23109
rect 38436 23072 38481 23100
rect 38436 23060 38442 23072
rect 40385 23069 40397 23103
rect 40385 23063 40408 23069
rect 40402 23060 40408 23063
rect 40460 23060 40466 23112
rect 40512 23109 40540 23140
rect 40604 23140 41420 23168
rect 40604 23109 40632 23140
rect 41414 23128 41420 23140
rect 41472 23128 41478 23180
rect 40497 23103 40555 23109
rect 40497 23069 40509 23103
rect 40543 23069 40555 23103
rect 40497 23063 40555 23069
rect 40594 23103 40652 23109
rect 40594 23069 40606 23103
rect 40640 23069 40652 23103
rect 40594 23063 40652 23069
rect 40773 23103 40831 23109
rect 40773 23069 40785 23103
rect 40819 23100 40831 23103
rect 41046 23100 41052 23112
rect 40819 23072 41052 23100
rect 40819 23069 40831 23072
rect 40773 23063 40831 23069
rect 20438 23032 20444 23044
rect 15856 23004 16160 23032
rect 20399 23004 20444 23032
rect 20438 22992 20444 23004
rect 20496 23032 20502 23044
rect 20993 23035 21051 23041
rect 20993 23032 21005 23035
rect 20496 23004 21005 23032
rect 20496 22992 20502 23004
rect 20993 23001 21005 23004
rect 21039 23001 21051 23035
rect 20993 22995 21051 23001
rect 22066 23004 23612 23032
rect 14976 22936 15056 22964
rect 14976 22924 14982 22936
rect 15286 22924 15292 22976
rect 15344 22964 15350 22976
rect 15381 22967 15439 22973
rect 15381 22964 15393 22967
rect 15344 22936 15393 22964
rect 15344 22924 15350 22936
rect 15381 22933 15393 22936
rect 15427 22933 15439 22967
rect 15381 22927 15439 22933
rect 17313 22967 17371 22973
rect 17313 22933 17325 22967
rect 17359 22964 17371 22967
rect 17402 22964 17408 22976
rect 17359 22936 17408 22964
rect 17359 22933 17371 22936
rect 17313 22927 17371 22933
rect 17402 22924 17408 22936
rect 17460 22924 17466 22976
rect 20530 22924 20536 22976
rect 20588 22964 20594 22976
rect 22066 22964 22094 23004
rect 22278 22964 22284 22976
rect 20588 22936 22094 22964
rect 22239 22936 22284 22964
rect 20588 22924 20594 22936
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 23584 22973 23612 23004
rect 25314 22992 25320 23044
rect 25372 23032 25378 23044
rect 28442 23032 28448 23044
rect 25372 23004 28448 23032
rect 25372 22992 25378 23004
rect 28442 22992 28448 23004
rect 28500 22992 28506 23044
rect 33410 22992 33416 23044
rect 33468 23032 33474 23044
rect 33882 23035 33940 23041
rect 33882 23032 33894 23035
rect 33468 23004 33894 23032
rect 33468 22992 33474 23004
rect 33882 23001 33894 23004
rect 33928 23001 33940 23035
rect 33882 22995 33940 23001
rect 35161 23035 35219 23041
rect 35161 23001 35173 23035
rect 35207 23001 35219 23035
rect 35161 22995 35219 23001
rect 35253 23035 35311 23041
rect 35253 23001 35265 23035
rect 35299 23032 35311 23035
rect 35986 23032 35992 23044
rect 35299 23004 35992 23032
rect 35299 23001 35311 23004
rect 35253 22995 35311 23001
rect 23569 22967 23627 22973
rect 23569 22933 23581 22967
rect 23615 22933 23627 22967
rect 23569 22927 23627 22933
rect 27249 22967 27307 22973
rect 27249 22933 27261 22967
rect 27295 22964 27307 22967
rect 27614 22964 27620 22976
rect 27295 22936 27620 22964
rect 27295 22933 27307 22936
rect 27249 22927 27307 22933
rect 27614 22924 27620 22936
rect 27672 22924 27678 22976
rect 28813 22967 28871 22973
rect 28813 22933 28825 22967
rect 28859 22964 28871 22967
rect 29362 22964 29368 22976
rect 28859 22936 29368 22964
rect 28859 22933 28871 22936
rect 28813 22927 28871 22933
rect 29362 22924 29368 22936
rect 29420 22924 29426 22976
rect 32306 22924 32312 22976
rect 32364 22964 32370 22976
rect 32769 22967 32827 22973
rect 32769 22964 32781 22967
rect 32364 22936 32781 22964
rect 32364 22924 32370 22936
rect 32769 22933 32781 22936
rect 32815 22964 32827 22967
rect 32858 22964 32864 22976
rect 32815 22936 32864 22964
rect 32815 22933 32827 22936
rect 32769 22927 32827 22933
rect 32858 22924 32864 22936
rect 32916 22924 32922 22976
rect 34146 22924 34152 22976
rect 34204 22964 34210 22976
rect 34885 22967 34943 22973
rect 34885 22964 34897 22967
rect 34204 22936 34897 22964
rect 34204 22924 34210 22936
rect 34885 22933 34897 22936
rect 34931 22933 34943 22967
rect 35176 22964 35204 22995
rect 35986 22992 35992 23004
rect 36044 22992 36050 23044
rect 37032 23035 37090 23041
rect 36096 23004 36952 23032
rect 36096 22964 36124 23004
rect 35176 22936 36124 22964
rect 36924 22964 36952 23004
rect 37032 23001 37044 23035
rect 37078 23032 37090 23035
rect 37737 23035 37795 23041
rect 37737 23032 37749 23035
rect 37078 23004 37749 23032
rect 37078 23001 37090 23004
rect 37032 22995 37090 23001
rect 37737 23001 37749 23004
rect 37783 23001 37795 23035
rect 40512 23032 40540 23063
rect 41046 23060 41052 23072
rect 41104 23060 41110 23112
rect 40954 23032 40960 23044
rect 40512 23004 40960 23032
rect 37737 22995 37795 23001
rect 40954 22992 40960 23004
rect 41012 22992 41018 23044
rect 38746 22964 38752 22976
rect 36924 22936 38752 22964
rect 34885 22927 34943 22933
rect 38746 22924 38752 22936
rect 38804 22924 38810 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1581 22763 1639 22769
rect 1581 22729 1593 22763
rect 1627 22760 1639 22763
rect 2774 22760 2780 22772
rect 1627 22732 2780 22760
rect 1627 22729 1639 22732
rect 1581 22723 1639 22729
rect 2774 22720 2780 22732
rect 2832 22720 2838 22772
rect 3786 22760 3792 22772
rect 3699 22732 3792 22760
rect 3786 22720 3792 22732
rect 3844 22760 3850 22772
rect 9214 22760 9220 22772
rect 3844 22732 9220 22760
rect 3844 22720 3850 22732
rect 9214 22720 9220 22732
rect 9272 22720 9278 22772
rect 11054 22720 11060 22772
rect 11112 22760 11118 22772
rect 15930 22760 15936 22772
rect 11112 22732 14780 22760
rect 15891 22732 15936 22760
rect 11112 22720 11118 22732
rect 1949 22695 2007 22701
rect 1949 22661 1961 22695
rect 1995 22692 2007 22695
rect 2222 22692 2228 22704
rect 1995 22664 2228 22692
rect 1995 22661 2007 22664
rect 1949 22655 2007 22661
rect 2222 22652 2228 22664
rect 2280 22652 2286 22704
rect 2590 22692 2596 22704
rect 2424 22664 2596 22692
rect 2424 22633 2452 22664
rect 2590 22652 2596 22664
rect 2648 22692 2654 22704
rect 2648 22664 6592 22692
rect 2648 22652 2654 22664
rect 2682 22633 2688 22636
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22593 1823 22627
rect 1765 22587 1823 22593
rect 2409 22627 2467 22633
rect 2409 22593 2421 22627
rect 2455 22593 2467 22627
rect 2676 22624 2688 22633
rect 2643 22596 2688 22624
rect 2409 22587 2467 22593
rect 2676 22587 2688 22596
rect 1780 22420 1808 22587
rect 2682 22584 2688 22587
rect 2740 22584 2746 22636
rect 4433 22627 4491 22633
rect 4433 22593 4445 22627
rect 4479 22593 4491 22627
rect 4614 22624 4620 22636
rect 4575 22596 4620 22624
rect 4433 22587 4491 22593
rect 4448 22556 4476 22587
rect 4614 22584 4620 22596
rect 4672 22624 4678 22636
rect 6564 22633 6592 22664
rect 8662 22652 8668 22704
rect 8720 22692 8726 22704
rect 9493 22695 9551 22701
rect 9493 22692 9505 22695
rect 8720 22664 9505 22692
rect 8720 22652 8726 22664
rect 9493 22661 9505 22664
rect 9539 22692 9551 22695
rect 10229 22695 10287 22701
rect 10229 22692 10241 22695
rect 9539 22664 10241 22692
rect 9539 22661 9551 22664
rect 9493 22655 9551 22661
rect 10229 22661 10241 22664
rect 10275 22692 10287 22695
rect 13262 22692 13268 22704
rect 10275 22664 13268 22692
rect 10275 22661 10287 22664
rect 10229 22655 10287 22661
rect 13262 22652 13268 22664
rect 13320 22652 13326 22704
rect 14458 22692 14464 22704
rect 14419 22664 14464 22692
rect 14458 22652 14464 22664
rect 14516 22652 14522 22704
rect 6822 22633 6828 22636
rect 5445 22627 5503 22633
rect 5445 22624 5457 22627
rect 4672 22596 5457 22624
rect 4672 22584 4678 22596
rect 5445 22593 5457 22596
rect 5491 22593 5503 22627
rect 5445 22587 5503 22593
rect 5629 22627 5687 22633
rect 5629 22593 5641 22627
rect 5675 22624 5687 22627
rect 6549 22627 6607 22633
rect 5675 22596 6500 22624
rect 5675 22593 5687 22596
rect 5629 22587 5687 22593
rect 4706 22556 4712 22568
rect 4448 22528 4712 22556
rect 4706 22516 4712 22528
rect 4764 22516 4770 22568
rect 3786 22420 3792 22432
rect 1780 22392 3792 22420
rect 3786 22380 3792 22392
rect 3844 22380 3850 22432
rect 4249 22423 4307 22429
rect 4249 22389 4261 22423
rect 4295 22420 4307 22423
rect 4614 22420 4620 22432
rect 4295 22392 4620 22420
rect 4295 22389 4307 22392
rect 4249 22383 4307 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 5813 22423 5871 22429
rect 5813 22389 5825 22423
rect 5859 22420 5871 22423
rect 6362 22420 6368 22432
rect 5859 22392 6368 22420
rect 5859 22389 5871 22392
rect 5813 22383 5871 22389
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 6472 22420 6500 22596
rect 6549 22593 6561 22627
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 6816 22587 6828 22633
rect 6880 22624 6886 22636
rect 8573 22627 8631 22633
rect 6880 22596 6916 22624
rect 6822 22584 6828 22587
rect 6880 22584 6886 22596
rect 8573 22593 8585 22627
rect 8619 22624 8631 22627
rect 9030 22624 9036 22636
rect 8619 22596 9036 22624
rect 8619 22593 8631 22596
rect 8573 22587 8631 22593
rect 9030 22584 9036 22596
rect 9088 22584 9094 22636
rect 9677 22627 9735 22633
rect 9677 22593 9689 22627
rect 9723 22624 9735 22627
rect 10042 22624 10048 22636
rect 9723 22596 10048 22624
rect 9723 22593 9735 22596
rect 9677 22587 9735 22593
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22593 11851 22627
rect 11793 22587 11851 22593
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22624 12035 22627
rect 12158 22624 12164 22636
rect 12023 22596 12164 22624
rect 12023 22593 12035 22596
rect 11977 22587 12035 22593
rect 7650 22516 7656 22568
rect 7708 22556 7714 22568
rect 8018 22556 8024 22568
rect 7708 22528 8024 22556
rect 7708 22516 7714 22528
rect 8018 22516 8024 22528
rect 8076 22516 8082 22568
rect 8938 22516 8944 22568
rect 8996 22556 9002 22568
rect 11808 22556 11836 22587
rect 12158 22584 12164 22596
rect 12216 22584 12222 22636
rect 14366 22624 14372 22636
rect 14327 22596 14372 22624
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 14752 22633 14780 22732
rect 15930 22720 15936 22732
rect 15988 22720 15994 22772
rect 16316 22732 18644 22760
rect 15381 22695 15439 22701
rect 15381 22661 15393 22695
rect 15427 22692 15439 22695
rect 16316 22692 16344 22732
rect 15427 22664 16344 22692
rect 18224 22695 18282 22701
rect 15427 22661 15439 22664
rect 15381 22655 15439 22661
rect 18224 22661 18236 22695
rect 18270 22692 18282 22695
rect 18506 22692 18512 22704
rect 18270 22664 18512 22692
rect 18270 22661 18282 22664
rect 18224 22655 18282 22661
rect 14553 22627 14611 22633
rect 14553 22593 14565 22627
rect 14599 22593 14611 22627
rect 14553 22587 14611 22593
rect 14737 22627 14795 22633
rect 14737 22593 14749 22627
rect 14783 22593 14795 22627
rect 14737 22587 14795 22593
rect 12529 22559 12587 22565
rect 12529 22556 12541 22559
rect 8996 22528 12541 22556
rect 8996 22516 9002 22528
rect 12529 22525 12541 22528
rect 12575 22556 12587 22559
rect 14182 22556 14188 22568
rect 12575 22528 14188 22556
rect 12575 22525 12587 22528
rect 12529 22519 12587 22525
rect 14182 22516 14188 22528
rect 14240 22516 14246 22568
rect 14568 22556 14596 22587
rect 14918 22556 14924 22568
rect 14568 22528 14924 22556
rect 14918 22516 14924 22528
rect 14976 22556 14982 22568
rect 15396 22556 15424 22655
rect 18506 22652 18512 22664
rect 18564 22652 18570 22704
rect 18616 22692 18644 22732
rect 19334 22720 19340 22772
rect 19392 22760 19398 22772
rect 20622 22760 20628 22772
rect 19392 22732 20628 22760
rect 19392 22720 19398 22732
rect 20622 22720 20628 22732
rect 20680 22720 20686 22772
rect 23106 22720 23112 22772
rect 23164 22760 23170 22772
rect 23753 22763 23811 22769
rect 23753 22760 23765 22763
rect 23164 22732 23765 22760
rect 23164 22720 23170 22732
rect 23753 22729 23765 22732
rect 23799 22760 23811 22763
rect 25222 22760 25228 22772
rect 23799 22732 24440 22760
rect 25183 22732 25228 22760
rect 23799 22729 23811 22732
rect 23753 22723 23811 22729
rect 23290 22692 23296 22704
rect 18616 22664 23296 22692
rect 23290 22652 23296 22664
rect 23348 22652 23354 22704
rect 24412 22701 24440 22732
rect 25222 22720 25228 22732
rect 25280 22760 25286 22772
rect 31573 22763 31631 22769
rect 25280 22732 26832 22760
rect 25280 22720 25286 22732
rect 24397 22695 24455 22701
rect 24397 22661 24409 22695
rect 24443 22661 24455 22695
rect 24397 22655 24455 22661
rect 24581 22695 24639 22701
rect 24581 22661 24593 22695
rect 24627 22692 24639 22695
rect 26694 22692 26700 22704
rect 24627 22664 26700 22692
rect 24627 22661 24639 22664
rect 24581 22655 24639 22661
rect 26694 22652 26700 22664
rect 26752 22652 26758 22704
rect 17402 22584 17408 22636
rect 17460 22624 17466 22636
rect 17957 22627 18015 22633
rect 17957 22624 17969 22627
rect 17460 22596 17969 22624
rect 17460 22584 17466 22596
rect 17957 22593 17969 22596
rect 18003 22593 18015 22627
rect 17957 22587 18015 22593
rect 18598 22584 18604 22636
rect 18656 22624 18662 22636
rect 20165 22627 20223 22633
rect 18656 22596 20024 22624
rect 18656 22584 18662 22596
rect 14976 22528 15424 22556
rect 14976 22516 14982 22528
rect 7929 22491 7987 22497
rect 7929 22457 7941 22491
rect 7975 22488 7987 22491
rect 14826 22488 14832 22500
rect 7975 22460 14832 22488
rect 7975 22457 7987 22460
rect 7929 22451 7987 22457
rect 7944 22420 7972 22451
rect 14826 22448 14832 22460
rect 14884 22448 14890 22500
rect 6472 22392 7972 22420
rect 8018 22380 8024 22432
rect 8076 22420 8082 22432
rect 8389 22423 8447 22429
rect 8389 22420 8401 22423
rect 8076 22392 8401 22420
rect 8076 22380 8082 22392
rect 8389 22389 8401 22392
rect 8435 22389 8447 22423
rect 11882 22420 11888 22432
rect 11843 22392 11888 22420
rect 8389 22383 8447 22389
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 14185 22423 14243 22429
rect 14185 22389 14197 22423
rect 14231 22420 14243 22423
rect 14550 22420 14556 22432
rect 14231 22392 14556 22420
rect 14231 22389 14243 22392
rect 14185 22383 14243 22389
rect 14550 22380 14556 22392
rect 14608 22380 14614 22432
rect 15746 22380 15752 22432
rect 15804 22420 15810 22432
rect 16669 22423 16727 22429
rect 16669 22420 16681 22423
rect 15804 22392 16681 22420
rect 15804 22380 15810 22392
rect 16669 22389 16681 22392
rect 16715 22389 16727 22423
rect 16669 22383 16727 22389
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19996 22429 20024 22596
rect 20165 22593 20177 22627
rect 20211 22624 20223 22627
rect 20806 22624 20812 22636
rect 20211 22596 20812 22624
rect 20211 22593 20223 22596
rect 20165 22587 20223 22593
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 21174 22624 21180 22636
rect 21135 22596 21180 22624
rect 21174 22584 21180 22596
rect 21232 22584 21238 22636
rect 25038 22624 25044 22636
rect 24999 22596 25044 22624
rect 25038 22584 25044 22596
rect 25096 22584 25102 22636
rect 26804 22624 26832 22732
rect 31573 22729 31585 22763
rect 31619 22760 31631 22763
rect 32766 22760 32772 22772
rect 31619 22732 32772 22760
rect 31619 22729 31631 22732
rect 31573 22723 31631 22729
rect 32766 22720 32772 22732
rect 32824 22720 32830 22772
rect 33410 22760 33416 22772
rect 33371 22732 33416 22760
rect 33410 22720 33416 22732
rect 33468 22720 33474 22772
rect 35618 22760 35624 22772
rect 35579 22732 35624 22760
rect 35618 22720 35624 22732
rect 35676 22720 35682 22772
rect 37277 22763 37335 22769
rect 37277 22729 37289 22763
rect 37323 22760 37335 22763
rect 38194 22760 38200 22772
rect 37323 22732 38200 22760
rect 37323 22729 37335 22732
rect 37277 22723 37335 22729
rect 38194 22720 38200 22732
rect 38252 22720 38258 22772
rect 40037 22763 40095 22769
rect 40037 22729 40049 22763
rect 40083 22760 40095 22763
rect 40310 22760 40316 22772
rect 40083 22732 40316 22760
rect 40083 22729 40095 22732
rect 40037 22723 40095 22729
rect 40310 22720 40316 22732
rect 40368 22720 40374 22772
rect 27157 22695 27215 22701
rect 27157 22661 27169 22695
rect 27203 22692 27215 22695
rect 27614 22692 27620 22704
rect 27203 22664 27620 22692
rect 27203 22661 27215 22664
rect 27157 22655 27215 22661
rect 27614 22652 27620 22664
rect 27672 22652 27678 22704
rect 28442 22692 28448 22704
rect 28403 22664 28448 22692
rect 28442 22652 28448 22664
rect 28500 22652 28506 22704
rect 29914 22652 29920 22704
rect 29972 22692 29978 22704
rect 31202 22692 31208 22704
rect 29972 22664 31208 22692
rect 29972 22652 29978 22664
rect 31202 22652 31208 22664
rect 31260 22652 31266 22704
rect 31297 22695 31355 22701
rect 31297 22661 31309 22695
rect 31343 22692 31355 22695
rect 32306 22692 32312 22704
rect 31343 22664 32312 22692
rect 31343 22661 31355 22664
rect 31297 22655 31355 22661
rect 32306 22652 32312 22664
rect 32364 22652 32370 22704
rect 33870 22692 33876 22704
rect 33831 22664 33876 22692
rect 33870 22652 33876 22664
rect 33928 22652 33934 22704
rect 35894 22692 35900 22704
rect 35855 22664 35900 22692
rect 35894 22652 35900 22664
rect 35952 22652 35958 22704
rect 36078 22652 36084 22704
rect 36136 22692 36142 22704
rect 37461 22695 37519 22701
rect 37461 22692 37473 22695
rect 36136 22664 37473 22692
rect 36136 22652 36142 22664
rect 37461 22661 37473 22664
rect 37507 22661 37519 22695
rect 37461 22655 37519 22661
rect 37645 22695 37703 22701
rect 37645 22661 37657 22695
rect 37691 22692 37703 22695
rect 40126 22692 40132 22704
rect 37691 22664 40132 22692
rect 37691 22661 37703 22664
rect 37645 22655 37703 22661
rect 40126 22652 40132 22664
rect 40184 22692 40190 22704
rect 40586 22692 40592 22704
rect 40184 22664 40592 22692
rect 40184 22652 40190 22664
rect 40586 22652 40592 22664
rect 40644 22652 40650 22704
rect 27341 22627 27399 22633
rect 27341 22624 27353 22627
rect 26804 22596 27353 22624
rect 27341 22593 27353 22596
rect 27387 22593 27399 22627
rect 28626 22624 28632 22636
rect 28587 22596 28632 22624
rect 27341 22587 27399 22593
rect 28626 22584 28632 22596
rect 28684 22584 28690 22636
rect 29730 22584 29736 22636
rect 29788 22624 29794 22636
rect 31021 22627 31079 22633
rect 31021 22624 31033 22627
rect 29788 22596 31033 22624
rect 29788 22584 29794 22596
rect 31021 22593 31033 22596
rect 31067 22593 31079 22627
rect 31386 22624 31392 22636
rect 31347 22596 31392 22624
rect 31021 22587 31079 22593
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 32582 22584 32588 22636
rect 32640 22624 32646 22636
rect 32769 22627 32827 22633
rect 32769 22624 32781 22627
rect 32640 22596 32781 22624
rect 32640 22584 32646 22596
rect 32769 22593 32781 22596
rect 32815 22593 32827 22627
rect 32932 22627 32990 22633
rect 32932 22624 32944 22627
rect 32769 22587 32827 22593
rect 32876 22596 32944 22624
rect 20073 22559 20131 22565
rect 20073 22525 20085 22559
rect 20119 22525 20131 22559
rect 20073 22519 20131 22525
rect 21085 22559 21143 22565
rect 21085 22525 21097 22559
rect 21131 22556 21143 22559
rect 32490 22556 32496 22568
rect 21131 22528 32496 22556
rect 21131 22525 21143 22528
rect 21085 22519 21143 22525
rect 20088 22488 20116 22519
rect 32490 22516 32496 22528
rect 32548 22516 32554 22568
rect 31754 22488 31760 22500
rect 20088 22460 31760 22488
rect 31754 22448 31760 22460
rect 31812 22448 31818 22500
rect 32876 22488 32904 22596
rect 32932 22593 32944 22596
rect 32978 22593 32990 22627
rect 32932 22587 32990 22593
rect 33045 22627 33103 22633
rect 33045 22593 33057 22627
rect 33091 22593 33103 22627
rect 33045 22587 33103 22593
rect 33137 22627 33195 22633
rect 33137 22593 33149 22627
rect 33183 22593 33195 22627
rect 34146 22624 34152 22636
rect 34107 22596 34152 22624
rect 33137 22587 33195 22593
rect 33060 22500 33088 22587
rect 32950 22488 32956 22500
rect 32876 22460 32956 22488
rect 32950 22448 32956 22460
rect 33008 22448 33014 22500
rect 33042 22448 33048 22500
rect 33100 22448 33106 22500
rect 33152 22488 33180 22587
rect 34146 22584 34152 22596
rect 34204 22584 34210 22636
rect 35802 22624 35808 22636
rect 35763 22596 35808 22624
rect 35802 22584 35808 22596
rect 35860 22584 35866 22636
rect 35986 22584 35992 22636
rect 36044 22624 36050 22636
rect 36173 22627 36231 22633
rect 36044 22596 36137 22624
rect 36044 22584 36050 22596
rect 36173 22593 36185 22627
rect 36219 22624 36231 22627
rect 37090 22624 37096 22636
rect 36219 22596 37096 22624
rect 36219 22593 36231 22596
rect 36173 22587 36231 22593
rect 37090 22584 37096 22596
rect 37148 22584 37154 22636
rect 37366 22584 37372 22636
rect 37424 22624 37430 22636
rect 38102 22624 38108 22636
rect 37424 22596 38108 22624
rect 37424 22584 37430 22596
rect 38102 22584 38108 22596
rect 38160 22624 38166 22636
rect 38197 22627 38255 22633
rect 38197 22624 38209 22627
rect 38160 22596 38209 22624
rect 38160 22584 38166 22596
rect 38197 22593 38209 22596
rect 38243 22593 38255 22627
rect 38197 22587 38255 22593
rect 38286 22584 38292 22636
rect 38344 22624 38350 22636
rect 38381 22627 38439 22633
rect 38381 22624 38393 22627
rect 38344 22596 38393 22624
rect 38344 22584 38350 22596
rect 38381 22593 38393 22596
rect 38427 22593 38439 22627
rect 38381 22587 38439 22593
rect 33778 22516 33784 22568
rect 33836 22556 33842 22568
rect 33965 22559 34023 22565
rect 33965 22556 33977 22559
rect 33836 22528 33977 22556
rect 33836 22516 33842 22528
rect 33965 22525 33977 22528
rect 34011 22525 34023 22559
rect 36004 22556 36032 22584
rect 36262 22556 36268 22568
rect 36004 22528 36268 22556
rect 33965 22519 34023 22525
rect 36262 22516 36268 22528
rect 36320 22516 36326 22568
rect 34330 22488 34336 22500
rect 33152 22460 34192 22488
rect 34291 22460 34336 22488
rect 19797 22423 19855 22429
rect 19797 22420 19809 22423
rect 19392 22392 19809 22420
rect 19392 22380 19398 22392
rect 19797 22389 19809 22392
rect 19843 22389 19855 22423
rect 19797 22383 19855 22389
rect 19981 22423 20039 22429
rect 19981 22389 19993 22423
rect 20027 22389 20039 22423
rect 19981 22383 20039 22389
rect 20809 22423 20867 22429
rect 20809 22389 20821 22423
rect 20855 22420 20867 22423
rect 20898 22420 20904 22432
rect 20855 22392 20904 22420
rect 20855 22389 20867 22392
rect 20809 22383 20867 22389
rect 20898 22380 20904 22392
rect 20956 22380 20962 22432
rect 20990 22380 20996 22432
rect 21048 22420 21054 22432
rect 21048 22392 21093 22420
rect 21048 22380 21054 22392
rect 25682 22380 25688 22432
rect 25740 22420 25746 22432
rect 26973 22423 27031 22429
rect 26973 22420 26985 22423
rect 25740 22392 26985 22420
rect 25740 22380 25746 22392
rect 26973 22389 26985 22392
rect 27019 22389 27031 22423
rect 26973 22383 27031 22389
rect 28261 22423 28319 22429
rect 28261 22389 28273 22423
rect 28307 22420 28319 22423
rect 28350 22420 28356 22432
rect 28307 22392 28356 22420
rect 28307 22389 28319 22392
rect 28261 22383 28319 22389
rect 28350 22380 28356 22392
rect 28408 22380 28414 22432
rect 30926 22380 30932 22432
rect 30984 22420 30990 22432
rect 31478 22420 31484 22432
rect 30984 22392 31484 22420
rect 30984 22380 30990 22392
rect 31478 22380 31484 22392
rect 31536 22420 31542 22432
rect 32217 22423 32275 22429
rect 32217 22420 32229 22423
rect 31536 22392 32229 22420
rect 31536 22380 31542 22392
rect 32217 22389 32229 22392
rect 32263 22420 32275 22423
rect 33152 22420 33180 22460
rect 33870 22420 33876 22432
rect 32263 22392 33180 22420
rect 33831 22392 33876 22420
rect 32263 22389 32275 22392
rect 32217 22383 32275 22389
rect 33870 22380 33876 22392
rect 33928 22380 33934 22432
rect 34164 22420 34192 22460
rect 34330 22448 34336 22460
rect 34388 22448 34394 22500
rect 41230 22488 41236 22500
rect 38488 22460 41236 22488
rect 38488 22420 38516 22460
rect 41230 22448 41236 22460
rect 41288 22448 41294 22500
rect 58158 22488 58164 22500
rect 58119 22460 58164 22488
rect 58158 22448 58164 22460
rect 58216 22448 58222 22500
rect 34164 22392 38516 22420
rect 38565 22423 38623 22429
rect 38565 22389 38577 22423
rect 38611 22420 38623 22423
rect 38930 22420 38936 22432
rect 38611 22392 38936 22420
rect 38611 22389 38623 22392
rect 38565 22383 38623 22389
rect 38930 22380 38936 22392
rect 38988 22380 38994 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 3234 22216 3240 22228
rect 3147 22188 3240 22216
rect 3234 22176 3240 22188
rect 3292 22216 3298 22228
rect 6822 22216 6828 22228
rect 3292 22188 5120 22216
rect 6783 22188 6828 22216
rect 3292 22176 3298 22188
rect 5092 22148 5120 22188
rect 6822 22176 6828 22188
rect 6880 22176 6886 22228
rect 8110 22216 8116 22228
rect 8071 22188 8116 22216
rect 8110 22176 8116 22188
rect 8168 22176 8174 22228
rect 14918 22216 14924 22228
rect 14879 22188 14924 22216
rect 14918 22176 14924 22188
rect 14976 22176 14982 22228
rect 21177 22219 21235 22225
rect 21177 22185 21189 22219
rect 21223 22216 21235 22219
rect 21266 22216 21272 22228
rect 21223 22188 21272 22216
rect 21223 22185 21235 22188
rect 21177 22179 21235 22185
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 31110 22176 31116 22228
rect 31168 22216 31174 22228
rect 31478 22216 31484 22228
rect 31168 22188 31484 22216
rect 31168 22176 31174 22188
rect 31478 22176 31484 22188
rect 31536 22176 31542 22228
rect 33321 22219 33379 22225
rect 33321 22185 33333 22219
rect 33367 22216 33379 22219
rect 33870 22216 33876 22228
rect 33367 22188 33876 22216
rect 33367 22185 33379 22188
rect 33321 22179 33379 22185
rect 33870 22176 33876 22188
rect 33928 22176 33934 22228
rect 37553 22219 37611 22225
rect 37553 22185 37565 22219
rect 37599 22216 37611 22219
rect 37826 22216 37832 22228
rect 37599 22188 37832 22216
rect 37599 22185 37611 22188
rect 37553 22179 37611 22185
rect 37826 22176 37832 22188
rect 37884 22216 37890 22228
rect 38286 22216 38292 22228
rect 37884 22188 38292 22216
rect 37884 22176 37890 22188
rect 38286 22176 38292 22188
rect 38344 22176 38350 22228
rect 5092 22120 9674 22148
rect 9646 22080 9674 22120
rect 11882 22108 11888 22160
rect 11940 22148 11946 22160
rect 16942 22148 16948 22160
rect 11940 22120 16948 22148
rect 11940 22108 11946 22120
rect 16942 22108 16948 22120
rect 17000 22108 17006 22160
rect 18230 22108 18236 22160
rect 18288 22148 18294 22160
rect 22005 22151 22063 22157
rect 22005 22148 22017 22151
rect 18288 22120 22017 22148
rect 18288 22108 18294 22120
rect 22005 22117 22017 22120
rect 22051 22148 22063 22151
rect 22462 22148 22468 22160
rect 22051 22120 22468 22148
rect 22051 22117 22063 22120
rect 22005 22111 22063 22117
rect 22462 22108 22468 22120
rect 22520 22108 22526 22160
rect 22922 22148 22928 22160
rect 22835 22120 22928 22148
rect 10152 22080 10456 22094
rect 15746 22080 15752 22092
rect 9646 22066 10456 22080
rect 9646 22052 10180 22066
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 2682 22012 2688 22024
rect 1903 21984 2688 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 2682 21972 2688 21984
rect 2740 22012 2746 22024
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 2740 21984 3801 22012
rect 2740 21972 2746 21984
rect 3789 21981 3801 21984
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 5166 21972 5172 22024
rect 5224 22012 5230 22024
rect 6086 22012 6092 22024
rect 5224 21984 6092 22012
rect 5224 21972 5230 21984
rect 6086 21972 6092 21984
rect 6144 22012 6150 22024
rect 6181 22015 6239 22021
rect 6181 22012 6193 22015
rect 6144 21984 6193 22012
rect 6144 21972 6150 21984
rect 6181 21981 6193 21984
rect 6227 21981 6239 22015
rect 6357 22012 6363 22024
rect 6318 21984 6363 22012
rect 6181 21975 6239 21981
rect 6357 21972 6363 21984
rect 6415 21972 6421 22024
rect 6457 22015 6515 22021
rect 6457 21981 6469 22015
rect 6503 21981 6515 22015
rect 6457 21975 6515 21981
rect 6595 22015 6653 22021
rect 6595 21981 6607 22015
rect 6641 21981 6653 22015
rect 7650 22012 7656 22024
rect 7611 21984 7656 22012
rect 6595 21975 6653 21981
rect 2130 21953 2136 21956
rect 2124 21907 2136 21953
rect 2188 21944 2194 21956
rect 2188 21916 2224 21944
rect 2130 21904 2136 21907
rect 2188 21904 2194 21916
rect 3602 21904 3608 21956
rect 3660 21944 3666 21956
rect 4034 21947 4092 21953
rect 4034 21944 4046 21947
rect 3660 21916 4046 21944
rect 3660 21904 3666 21916
rect 4034 21913 4046 21916
rect 4080 21913 4092 21947
rect 4034 21907 4092 21913
rect 5994 21904 6000 21956
rect 6052 21944 6058 21956
rect 6472 21944 6500 21975
rect 6052 21916 6500 21944
rect 6625 21944 6653 21975
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 9214 21972 9220 22024
rect 9272 22012 9278 22024
rect 9861 22015 9919 22021
rect 9861 22012 9873 22015
rect 9272 21984 9873 22012
rect 9272 21972 9278 21984
rect 9861 21981 9873 21984
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 10318 22012 10324 22024
rect 10275 21984 10324 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 10318 21972 10324 21984
rect 10376 21972 10382 22024
rect 10428 22012 10456 22066
rect 15707 22052 15752 22080
rect 15746 22040 15752 22052
rect 15804 22040 15810 22092
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 10428 21984 11437 22012
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11698 22012 11704 22024
rect 11659 21984 11704 22012
rect 11425 21975 11483 21981
rect 11698 21972 11704 21984
rect 11756 21972 11762 22024
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 22012 11851 22015
rect 12434 22012 12440 22024
rect 11839 21984 12440 22012
rect 11839 21981 11851 21984
rect 11793 21975 11851 21981
rect 12434 21972 12440 21984
rect 12492 22012 12498 22024
rect 13354 22012 13360 22024
rect 12492 21984 13360 22012
rect 12492 21972 12498 21984
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13541 22015 13599 22021
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13587 21984 14105 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 14093 21981 14105 21984
rect 14139 22012 14151 22015
rect 14826 22012 14832 22024
rect 14139 21984 14832 22012
rect 14139 21981 14151 21984
rect 14093 21975 14151 21981
rect 14826 21972 14832 21984
rect 14884 22012 14890 22024
rect 15378 22012 15384 22024
rect 14884 21984 15384 22012
rect 14884 21972 14890 21984
rect 15378 21972 15384 21984
rect 15436 21972 15442 22024
rect 15565 22015 15623 22021
rect 15565 21981 15577 22015
rect 15611 21981 15623 22015
rect 15565 21975 15623 21981
rect 16761 22015 16819 22021
rect 16761 21981 16773 22015
rect 16807 21981 16819 22015
rect 16761 21975 16819 21981
rect 17037 22015 17095 22021
rect 17037 21981 17049 22015
rect 17083 22012 17095 22015
rect 17126 22012 17132 22024
rect 17083 21984 17132 22012
rect 17083 21981 17095 21984
rect 17037 21975 17095 21981
rect 7469 21947 7527 21953
rect 6625 21916 7420 21944
rect 6052 21904 6058 21916
rect 4706 21836 4712 21888
rect 4764 21876 4770 21888
rect 5169 21879 5227 21885
rect 5169 21876 5181 21879
rect 4764 21848 5181 21876
rect 4764 21836 4770 21848
rect 5169 21845 5181 21848
rect 5215 21876 5227 21879
rect 5258 21876 5264 21888
rect 5215 21848 5264 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 5902 21836 5908 21888
rect 5960 21876 5966 21888
rect 7285 21879 7343 21885
rect 7285 21876 7297 21879
rect 5960 21848 7297 21876
rect 5960 21836 5966 21848
rect 7285 21845 7297 21848
rect 7331 21845 7343 21879
rect 7392 21876 7420 21916
rect 7469 21913 7481 21947
rect 7515 21944 7527 21947
rect 7742 21944 7748 21956
rect 7515 21916 7748 21944
rect 7515 21913 7527 21916
rect 7469 21907 7527 21913
rect 7742 21904 7748 21916
rect 7800 21904 7806 21956
rect 10042 21944 10048 21956
rect 10003 21916 10048 21944
rect 10042 21904 10048 21916
rect 10100 21904 10106 21956
rect 10137 21947 10195 21953
rect 10137 21913 10149 21947
rect 10183 21944 10195 21947
rect 11606 21944 11612 21956
rect 10183 21916 10272 21944
rect 11567 21916 11612 21944
rect 10183 21913 10195 21916
rect 10137 21907 10195 21913
rect 10244 21888 10272 21916
rect 11606 21904 11612 21916
rect 11664 21944 11670 21956
rect 12158 21944 12164 21956
rect 11664 21916 12164 21944
rect 11664 21904 11670 21916
rect 12158 21904 12164 21916
rect 12216 21944 12222 21956
rect 15580 21944 15608 21975
rect 16776 21944 16804 21975
rect 17126 21972 17132 21984
rect 17184 22012 17190 22024
rect 17678 22012 17684 22024
rect 17184 21984 17684 22012
rect 17184 21972 17190 21984
rect 17678 21972 17684 21984
rect 17736 21972 17742 22024
rect 21082 22012 21088 22024
rect 21043 21984 21088 22012
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 22012 21235 22015
rect 22094 22012 22100 22024
rect 21223 21984 22100 22012
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 22094 21972 22100 21984
rect 22152 21972 22158 22024
rect 22186 21972 22192 22024
rect 22244 22012 22250 22024
rect 22557 22015 22615 22021
rect 22557 22012 22569 22015
rect 22244 21984 22569 22012
rect 22244 21972 22250 21984
rect 22557 21981 22569 21984
rect 22603 21981 22615 22015
rect 22738 22012 22744 22024
rect 22699 21984 22744 22012
rect 22557 21975 22615 21981
rect 22738 21972 22744 21984
rect 22796 21972 22802 22024
rect 22848 22021 22876 22120
rect 22922 22108 22928 22120
rect 22980 22148 22986 22160
rect 23382 22148 23388 22160
rect 22980 22120 23388 22148
rect 22980 22108 22986 22120
rect 23382 22108 23388 22120
rect 23440 22108 23446 22160
rect 31386 22108 31392 22160
rect 31444 22148 31450 22160
rect 33134 22148 33140 22160
rect 31444 22120 33140 22148
rect 31444 22108 31450 22120
rect 26878 22040 26884 22092
rect 26936 22080 26942 22092
rect 26936 22052 27752 22080
rect 26936 22040 26942 22052
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 22925 22015 22983 22021
rect 22925 21981 22937 22015
rect 22971 21981 22983 22015
rect 22925 21975 22983 21981
rect 12216 21916 16804 21944
rect 12216 21904 12222 21916
rect 22462 21904 22468 21956
rect 22520 21944 22526 21956
rect 22940 21944 22968 21975
rect 27430 21972 27436 22024
rect 27488 22012 27494 22024
rect 27617 22015 27675 22021
rect 27617 22012 27629 22015
rect 27488 21984 27629 22012
rect 27488 21972 27494 21984
rect 27617 21981 27629 21984
rect 27663 21981 27675 22015
rect 27724 22012 27752 22052
rect 31757 22015 31815 22021
rect 31757 22012 31769 22015
rect 27724 21984 31769 22012
rect 27617 21975 27675 21981
rect 31757 21981 31769 21984
rect 31803 21981 31815 22015
rect 31757 21975 31815 21981
rect 31846 21972 31852 22024
rect 31904 22012 31910 22024
rect 32025 22015 32083 22021
rect 32025 22012 32037 22015
rect 31904 21984 32037 22012
rect 31904 21972 31910 21984
rect 32025 21981 32037 21984
rect 32071 21981 32083 22015
rect 32025 21975 32083 21981
rect 32171 22015 32229 22021
rect 32171 21981 32183 22015
rect 32217 22012 32229 22015
rect 32324 22012 32352 22120
rect 33134 22108 33140 22120
rect 33192 22108 33198 22160
rect 33686 22080 33692 22092
rect 33060 22052 33692 22080
rect 32766 22012 32772 22024
rect 32217 21984 32352 22012
rect 32727 21984 32772 22012
rect 32217 21981 32229 21984
rect 32171 21975 32229 21981
rect 32766 21972 32772 21984
rect 32824 21972 32830 22024
rect 33060 22021 33088 22052
rect 33686 22040 33692 22052
rect 33744 22040 33750 22092
rect 33045 22015 33103 22021
rect 33045 21981 33057 22015
rect 33091 21981 33103 22015
rect 33045 21975 33103 21981
rect 33134 21972 33140 22024
rect 33192 22012 33198 22024
rect 33192 21984 33237 22012
rect 33192 21972 33198 21984
rect 38838 21972 38844 22024
rect 38896 22012 38902 22024
rect 38933 22015 38991 22021
rect 38933 22012 38945 22015
rect 38896 21984 38945 22012
rect 38896 21972 38902 21984
rect 38933 21981 38945 21984
rect 38979 21981 38991 22015
rect 38933 21975 38991 21981
rect 27890 21953 27896 21956
rect 22520 21916 22968 21944
rect 22520 21904 22526 21916
rect 27884 21907 27896 21953
rect 27948 21944 27954 21956
rect 27948 21916 27984 21944
rect 27890 21904 27896 21907
rect 27948 21904 27954 21916
rect 28718 21904 28724 21956
rect 28776 21944 28782 21956
rect 30834 21944 30840 21956
rect 28776 21916 30840 21944
rect 28776 21904 28782 21916
rect 30834 21904 30840 21916
rect 30892 21904 30898 21956
rect 31202 21904 31208 21956
rect 31260 21944 31266 21956
rect 31941 21947 31999 21953
rect 31941 21944 31953 21947
rect 31260 21916 31953 21944
rect 31260 21904 31266 21916
rect 31941 21913 31953 21916
rect 31987 21944 31999 21947
rect 32953 21947 33011 21953
rect 32953 21944 32965 21947
rect 31987 21916 32965 21944
rect 31987 21913 31999 21916
rect 31941 21907 31999 21913
rect 32953 21913 32965 21916
rect 32999 21913 33011 21947
rect 32953 21907 33011 21913
rect 38470 21904 38476 21956
rect 38528 21944 38534 21956
rect 38666 21947 38724 21953
rect 38666 21944 38678 21947
rect 38528 21916 38678 21944
rect 38528 21904 38534 21916
rect 38666 21913 38678 21916
rect 38712 21913 38724 21947
rect 38666 21907 38724 21913
rect 8110 21876 8116 21888
rect 7392 21848 8116 21876
rect 7285 21839 7343 21845
rect 8110 21836 8116 21848
rect 8168 21836 8174 21888
rect 9030 21876 9036 21888
rect 8991 21848 9036 21876
rect 9030 21836 9036 21848
rect 9088 21836 9094 21888
rect 10226 21836 10232 21888
rect 10284 21836 10290 21888
rect 10413 21879 10471 21885
rect 10413 21845 10425 21879
rect 10459 21876 10471 21879
rect 10962 21876 10968 21888
rect 10459 21848 10968 21876
rect 10459 21845 10471 21848
rect 10413 21839 10471 21845
rect 10962 21836 10968 21848
rect 11020 21836 11026 21888
rect 11977 21879 12035 21885
rect 11977 21845 11989 21879
rect 12023 21876 12035 21879
rect 12066 21876 12072 21888
rect 12023 21848 12072 21876
rect 12023 21845 12035 21848
rect 11977 21839 12035 21845
rect 12066 21836 12072 21848
rect 12124 21836 12130 21888
rect 13538 21836 13544 21888
rect 13596 21876 13602 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13596 21848 14289 21876
rect 13596 21836 13602 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 15378 21876 15384 21888
rect 15339 21848 15384 21876
rect 14277 21839 14335 21845
rect 15378 21836 15384 21848
rect 15436 21876 15442 21888
rect 15838 21876 15844 21888
rect 15436 21848 15844 21876
rect 15436 21836 15442 21848
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 20809 21879 20867 21885
rect 20809 21845 20821 21879
rect 20855 21876 20867 21879
rect 21174 21876 21180 21888
rect 20855 21848 21180 21876
rect 20855 21845 20867 21848
rect 20809 21839 20867 21845
rect 21174 21836 21180 21848
rect 21232 21836 21238 21888
rect 22646 21836 22652 21888
rect 22704 21876 22710 21888
rect 23106 21876 23112 21888
rect 22704 21848 23112 21876
rect 22704 21836 22710 21848
rect 23106 21836 23112 21848
rect 23164 21836 23170 21888
rect 23201 21879 23259 21885
rect 23201 21845 23213 21879
rect 23247 21876 23259 21879
rect 23290 21876 23296 21888
rect 23247 21848 23296 21876
rect 23247 21845 23259 21848
rect 23201 21839 23259 21845
rect 23290 21836 23296 21848
rect 23348 21836 23354 21888
rect 28442 21836 28448 21888
rect 28500 21876 28506 21888
rect 28997 21879 29055 21885
rect 28997 21876 29009 21879
rect 28500 21848 29009 21876
rect 28500 21836 28506 21848
rect 28997 21845 29009 21848
rect 29043 21845 29055 21879
rect 28997 21839 29055 21845
rect 32309 21879 32367 21885
rect 32309 21845 32321 21879
rect 32355 21876 32367 21879
rect 32674 21876 32680 21888
rect 32355 21848 32680 21876
rect 32355 21845 32367 21848
rect 32309 21839 32367 21845
rect 32674 21836 32680 21848
rect 32732 21836 32738 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 2130 21672 2136 21684
rect 2091 21644 2136 21672
rect 2130 21632 2136 21644
rect 2188 21632 2194 21684
rect 3602 21672 3608 21684
rect 3563 21644 3608 21672
rect 3602 21632 3608 21644
rect 3660 21632 3666 21684
rect 5994 21672 6000 21684
rect 3988 21644 6000 21672
rect 3050 21604 3056 21616
rect 2516 21576 3056 21604
rect 2516 21545 2544 21576
rect 3050 21564 3056 21576
rect 3108 21604 3114 21616
rect 3988 21604 4016 21644
rect 4614 21604 4620 21616
rect 3108 21576 4016 21604
rect 3108 21564 3114 21576
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21505 2467 21539
rect 2409 21499 2467 21505
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21505 2559 21539
rect 2501 21499 2559 21505
rect 2424 21400 2452 21499
rect 2590 21496 2596 21548
rect 2648 21536 2654 21548
rect 2777 21539 2835 21545
rect 2648 21508 2693 21536
rect 2648 21496 2654 21508
rect 2777 21505 2789 21539
rect 2823 21505 2835 21539
rect 3878 21536 3884 21548
rect 3839 21508 3884 21536
rect 2777 21499 2835 21505
rect 2792 21468 2820 21499
rect 3878 21496 3884 21508
rect 3936 21496 3942 21548
rect 3988 21545 4016 21576
rect 4080 21576 4620 21604
rect 4080 21545 4108 21576
rect 4614 21564 4620 21576
rect 4672 21564 4678 21616
rect 5414 21604 5442 21644
rect 5994 21632 6000 21644
rect 6052 21672 6058 21684
rect 7374 21672 7380 21684
rect 6052 21644 7380 21672
rect 6052 21632 6058 21644
rect 7374 21632 7380 21644
rect 7432 21632 7438 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 11606 21672 11612 21684
rect 10100 21644 11612 21672
rect 10100 21632 10106 21644
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 14366 21632 14372 21684
rect 14424 21672 14430 21684
rect 14829 21675 14887 21681
rect 14829 21672 14841 21675
rect 14424 21644 14841 21672
rect 14424 21632 14430 21644
rect 14829 21641 14841 21644
rect 14875 21641 14887 21675
rect 14829 21635 14887 21641
rect 15562 21632 15568 21684
rect 15620 21672 15626 21684
rect 15657 21675 15715 21681
rect 15657 21672 15669 21675
rect 15620 21644 15669 21672
rect 15620 21632 15626 21644
rect 15657 21641 15669 21644
rect 15703 21672 15715 21675
rect 15703 21644 21036 21672
rect 15703 21641 15715 21644
rect 15657 21635 15715 21641
rect 5813 21607 5871 21613
rect 5414 21576 5488 21604
rect 3973 21539 4031 21545
rect 3973 21505 3985 21539
rect 4019 21505 4031 21539
rect 3973 21499 4031 21505
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4249 21539 4307 21545
rect 4249 21505 4261 21539
rect 4295 21536 4307 21539
rect 5166 21536 5172 21548
rect 4295 21508 5172 21536
rect 4295 21505 4307 21508
rect 4249 21499 4307 21505
rect 2958 21468 2964 21480
rect 2792 21440 2964 21468
rect 2958 21428 2964 21440
rect 3016 21468 3022 21480
rect 4264 21468 4292 21499
rect 5166 21496 5172 21508
rect 5224 21496 5230 21548
rect 5332 21545 5390 21551
rect 5460 21545 5488 21576
rect 5813 21573 5825 21607
rect 5859 21604 5871 21607
rect 6610 21607 6668 21613
rect 6610 21604 6622 21607
rect 5859 21576 6622 21604
rect 5859 21573 5871 21576
rect 5813 21567 5871 21573
rect 6610 21573 6622 21576
rect 6656 21573 6668 21607
rect 10134 21604 10140 21616
rect 10095 21576 10140 21604
rect 6610 21567 6668 21573
rect 10134 21564 10140 21576
rect 10192 21564 10198 21616
rect 14277 21607 14335 21613
rect 14277 21573 14289 21607
rect 14323 21604 14335 21607
rect 14458 21604 14464 21616
rect 14323 21576 14464 21604
rect 14323 21573 14335 21576
rect 14277 21567 14335 21573
rect 14458 21564 14464 21576
rect 14516 21604 14522 21616
rect 20073 21607 20131 21613
rect 20073 21604 20085 21607
rect 14516 21576 20085 21604
rect 14516 21564 14522 21576
rect 20073 21573 20085 21576
rect 20119 21604 20131 21607
rect 20717 21607 20775 21613
rect 20717 21604 20729 21607
rect 20119 21576 20729 21604
rect 20119 21573 20131 21576
rect 20073 21567 20131 21573
rect 20717 21573 20729 21576
rect 20763 21573 20775 21607
rect 21008 21604 21036 21644
rect 21082 21632 21088 21684
rect 21140 21672 21146 21684
rect 33502 21672 33508 21684
rect 21140 21644 33508 21672
rect 21140 21632 21146 21644
rect 33502 21632 33508 21644
rect 33560 21632 33566 21684
rect 38470 21672 38476 21684
rect 38431 21644 38476 21672
rect 38470 21632 38476 21644
rect 38528 21632 38534 21684
rect 21634 21604 21640 21616
rect 21008 21576 21640 21604
rect 20717 21567 20775 21573
rect 21634 21564 21640 21576
rect 21692 21564 21698 21616
rect 23008 21607 23066 21613
rect 23008 21573 23020 21607
rect 23054 21604 23066 21607
rect 23106 21604 23112 21616
rect 23054 21576 23112 21604
rect 23054 21573 23066 21576
rect 23008 21567 23066 21573
rect 23106 21564 23112 21576
rect 23164 21564 23170 21616
rect 24949 21607 25007 21613
rect 24949 21573 24961 21607
rect 24995 21604 25007 21607
rect 25038 21604 25044 21616
rect 24995 21576 25044 21604
rect 24995 21573 25007 21576
rect 24949 21567 25007 21573
rect 25038 21564 25044 21576
rect 25096 21564 25102 21616
rect 27890 21604 27896 21616
rect 27851 21576 27896 21604
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 28442 21564 28448 21616
rect 28500 21564 28506 21616
rect 32858 21564 32864 21616
rect 32916 21604 32922 21616
rect 32953 21607 33011 21613
rect 32953 21604 32965 21607
rect 32916 21576 32965 21604
rect 32916 21564 32922 21576
rect 32953 21573 32965 21576
rect 32999 21573 33011 21607
rect 34790 21604 34796 21616
rect 32953 21567 33011 21573
rect 33060 21576 34796 21604
rect 5332 21542 5344 21545
rect 5276 21514 5344 21542
rect 3016 21440 4292 21468
rect 5276 21468 5304 21514
rect 5332 21511 5344 21514
rect 5378 21511 5390 21545
rect 5332 21505 5390 21511
rect 5445 21539 5503 21545
rect 5445 21505 5457 21539
rect 5491 21505 5503 21539
rect 5445 21499 5503 21505
rect 5537 21539 5595 21545
rect 5537 21505 5549 21539
rect 5583 21536 5672 21539
rect 5718 21536 5724 21548
rect 5583 21511 5724 21536
rect 5583 21505 5595 21511
rect 5644 21508 5724 21511
rect 5537 21499 5595 21505
rect 5718 21496 5724 21508
rect 5776 21496 5782 21548
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 6104 21508 9873 21536
rect 5902 21468 5908 21480
rect 5276 21440 5908 21468
rect 3016 21428 3022 21440
rect 5902 21428 5908 21440
rect 5960 21428 5966 21480
rect 2774 21400 2780 21412
rect 2424 21372 2780 21400
rect 2774 21360 2780 21372
rect 2832 21360 2838 21412
rect 5258 21360 5264 21412
rect 5316 21400 5322 21412
rect 6104 21400 6132 21508
rect 9861 21505 9873 21508
rect 9907 21505 9919 21539
rect 10042 21536 10048 21548
rect 10003 21508 10048 21536
rect 9861 21499 9919 21505
rect 10042 21496 10048 21508
rect 10100 21496 10106 21548
rect 10229 21539 10287 21545
rect 10229 21505 10241 21539
rect 10275 21536 10287 21539
rect 10318 21536 10324 21548
rect 10275 21508 10324 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 10318 21496 10324 21508
rect 10376 21536 10382 21548
rect 12434 21536 12440 21548
rect 10376 21508 12440 21536
rect 10376 21496 10382 21508
rect 12434 21496 12440 21508
rect 12492 21496 12498 21548
rect 15746 21536 15752 21548
rect 15707 21508 15752 21536
rect 15746 21496 15752 21508
rect 15804 21496 15810 21548
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16224 21508 17049 21536
rect 6362 21468 6368 21480
rect 6323 21440 6368 21468
rect 6362 21428 6368 21440
rect 6420 21428 6426 21480
rect 9030 21428 9036 21480
rect 9088 21468 9094 21480
rect 9088 21440 12434 21468
rect 9088 21428 9094 21440
rect 7742 21400 7748 21412
rect 5316 21372 6132 21400
rect 7655 21372 7748 21400
rect 5316 21360 5322 21372
rect 7742 21360 7748 21372
rect 7800 21400 7806 21412
rect 11054 21400 11060 21412
rect 7800 21372 11060 21400
rect 7800 21360 7806 21372
rect 11054 21360 11060 21372
rect 11112 21360 11118 21412
rect 12406 21400 12434 21440
rect 13538 21428 13544 21480
rect 13596 21468 13602 21480
rect 16224 21468 16252 21508
rect 17037 21505 17049 21508
rect 17083 21505 17095 21539
rect 17037 21499 17095 21505
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21505 17187 21539
rect 17129 21499 17187 21505
rect 13596 21440 16252 21468
rect 13596 21428 13602 21440
rect 15378 21400 15384 21412
rect 12406 21372 15384 21400
rect 15378 21360 15384 21372
rect 15436 21360 15442 21412
rect 16224 21400 16252 21440
rect 16942 21428 16948 21480
rect 17000 21468 17006 21480
rect 17144 21468 17172 21499
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 17405 21539 17463 21545
rect 17276 21508 17321 21536
rect 17276 21496 17282 21508
rect 17405 21505 17417 21539
rect 17451 21536 17463 21539
rect 17770 21536 17776 21548
rect 17451 21508 17776 21536
rect 17451 21505 17463 21508
rect 17405 21499 17463 21505
rect 17770 21496 17776 21508
rect 17828 21536 17834 21548
rect 20533 21539 20591 21545
rect 20533 21536 20545 21539
rect 17828 21508 20545 21536
rect 17828 21496 17834 21508
rect 20533 21505 20545 21508
rect 20579 21505 20591 21539
rect 20533 21499 20591 21505
rect 22554 21496 22560 21548
rect 22612 21536 22618 21548
rect 24581 21539 24639 21545
rect 24581 21536 24593 21539
rect 22612 21508 24593 21536
rect 22612 21496 22618 21508
rect 24581 21505 24593 21508
rect 24627 21505 24639 21539
rect 24581 21499 24639 21505
rect 24670 21496 24676 21548
rect 24728 21536 24734 21548
rect 24765 21539 24823 21545
rect 24765 21536 24777 21539
rect 24728 21508 24777 21536
rect 24728 21496 24734 21508
rect 24765 21505 24777 21508
rect 24811 21505 24823 21539
rect 24765 21499 24823 21505
rect 27433 21539 27491 21545
rect 27433 21505 27445 21539
rect 27479 21536 27491 21539
rect 27706 21536 27712 21548
rect 27479 21508 27712 21536
rect 27479 21505 27491 21508
rect 27433 21499 27491 21505
rect 27706 21496 27712 21508
rect 27764 21536 27770 21548
rect 28123 21539 28181 21545
rect 28123 21536 28135 21539
rect 27764 21508 28135 21536
rect 27764 21496 27770 21508
rect 28123 21505 28135 21508
rect 28169 21505 28181 21539
rect 28258 21536 28264 21548
rect 28219 21508 28264 21536
rect 28123 21499 28181 21505
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 28358 21545 28416 21551
rect 28358 21511 28370 21545
rect 28404 21536 28416 21545
rect 28460 21536 28488 21564
rect 28404 21511 28488 21536
rect 28358 21508 28488 21511
rect 28537 21539 28595 21545
rect 28358 21505 28416 21508
rect 28537 21505 28549 21539
rect 28583 21536 28595 21539
rect 28997 21539 29055 21545
rect 28997 21536 29009 21539
rect 28583 21508 29009 21536
rect 28583 21505 28595 21508
rect 28537 21499 28595 21505
rect 28997 21505 29009 21508
rect 29043 21505 29055 21539
rect 28997 21499 29055 21505
rect 29733 21539 29791 21545
rect 29733 21505 29745 21539
rect 29779 21505 29791 21539
rect 29733 21499 29791 21505
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 33060 21536 33088 21576
rect 34790 21564 34796 21576
rect 34848 21564 34854 21616
rect 30055 21508 33088 21536
rect 33137 21539 33195 21545
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 33137 21505 33149 21539
rect 33183 21536 33195 21539
rect 33318 21536 33324 21548
rect 33183 21508 33324 21536
rect 33183 21505 33195 21508
rect 33137 21499 33195 21505
rect 17000 21440 17172 21468
rect 17000 21428 17006 21440
rect 20070 21428 20076 21480
rect 20128 21468 20134 21480
rect 22646 21468 22652 21480
rect 20128 21440 22652 21468
rect 20128 21428 20134 21440
rect 22646 21428 22652 21440
rect 22704 21428 22710 21480
rect 22741 21471 22799 21477
rect 22741 21437 22753 21471
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 17865 21403 17923 21409
rect 17865 21400 17877 21403
rect 16224 21372 17877 21400
rect 17865 21369 17877 21372
rect 17911 21400 17923 21403
rect 21818 21400 21824 21412
rect 17911 21372 21824 21400
rect 17911 21369 17923 21372
rect 17865 21363 17923 21369
rect 21818 21360 21824 21372
rect 21876 21360 21882 21412
rect 10413 21335 10471 21341
rect 10413 21301 10425 21335
rect 10459 21332 10471 21335
rect 10594 21332 10600 21344
rect 10459 21304 10600 21332
rect 10459 21301 10471 21304
rect 10413 21295 10471 21301
rect 10594 21292 10600 21304
rect 10652 21292 10658 21344
rect 16758 21332 16764 21344
rect 16719 21304 16764 21332
rect 16758 21292 16764 21304
rect 16816 21292 16822 21344
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 22189 21335 22247 21341
rect 22189 21332 22201 21335
rect 22152 21304 22201 21332
rect 22152 21292 22158 21304
rect 22189 21301 22201 21304
rect 22235 21301 22247 21335
rect 22756 21332 22784 21431
rect 26418 21360 26424 21412
rect 26476 21400 26482 21412
rect 28552 21400 28580 21499
rect 29546 21400 29552 21412
rect 26476 21372 28580 21400
rect 29507 21372 29552 21400
rect 26476 21360 26482 21372
rect 29546 21360 29552 21372
rect 29604 21360 29610 21412
rect 29748 21400 29776 21499
rect 33318 21496 33324 21508
rect 33376 21496 33382 21548
rect 38654 21536 38660 21548
rect 37936 21508 38660 21536
rect 29917 21471 29975 21477
rect 29917 21437 29929 21471
rect 29963 21468 29975 21471
rect 30098 21468 30104 21480
rect 29963 21440 30104 21468
rect 29963 21437 29975 21440
rect 29917 21431 29975 21437
rect 30098 21428 30104 21440
rect 30156 21428 30162 21480
rect 32769 21471 32827 21477
rect 32769 21437 32781 21471
rect 32815 21468 32827 21471
rect 32950 21468 32956 21480
rect 32815 21440 32956 21468
rect 32815 21437 32827 21440
rect 32769 21431 32827 21437
rect 32950 21428 32956 21440
rect 33008 21428 33014 21480
rect 37274 21400 37280 21412
rect 29748 21372 37280 21400
rect 37274 21360 37280 21372
rect 37332 21360 37338 21412
rect 23014 21332 23020 21344
rect 22756 21304 23020 21332
rect 22189 21295 22247 21301
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 24121 21335 24179 21341
rect 24121 21301 24133 21335
rect 24167 21332 24179 21335
rect 24670 21332 24676 21344
rect 24167 21304 24676 21332
rect 24167 21301 24179 21304
rect 24121 21295 24179 21301
rect 24670 21292 24676 21304
rect 24728 21292 24734 21344
rect 29822 21332 29828 21344
rect 29783 21304 29828 21332
rect 29822 21292 29828 21304
rect 29880 21292 29886 21344
rect 32950 21292 32956 21344
rect 33008 21332 33014 21344
rect 37936 21341 37964 21508
rect 38654 21496 38660 21508
rect 38712 21536 38718 21548
rect 38749 21539 38807 21545
rect 38749 21536 38761 21539
rect 38712 21508 38761 21536
rect 38712 21496 38718 21508
rect 38749 21505 38761 21508
rect 38795 21505 38807 21539
rect 38749 21499 38807 21505
rect 38841 21539 38899 21545
rect 38841 21505 38853 21539
rect 38887 21505 38899 21539
rect 38841 21499 38899 21505
rect 38856 21468 38884 21499
rect 38930 21496 38936 21548
rect 38988 21536 38994 21548
rect 39117 21539 39175 21545
rect 38988 21508 39033 21536
rect 38988 21496 38994 21508
rect 39117 21505 39129 21539
rect 39163 21536 39175 21539
rect 39758 21536 39764 21548
rect 39163 21508 39764 21536
rect 39163 21505 39175 21508
rect 39117 21499 39175 21505
rect 39758 21496 39764 21508
rect 39816 21496 39822 21548
rect 40034 21468 40040 21480
rect 38856 21440 40040 21468
rect 40034 21428 40040 21440
rect 40092 21468 40098 21480
rect 40862 21468 40868 21480
rect 40092 21440 40868 21468
rect 40092 21428 40098 21440
rect 40862 21428 40868 21440
rect 40920 21428 40926 21480
rect 37921 21335 37979 21341
rect 37921 21332 37933 21335
rect 33008 21304 37933 21332
rect 33008 21292 33014 21304
rect 37921 21301 37933 21304
rect 37967 21301 37979 21335
rect 58158 21332 58164 21344
rect 58119 21304 58164 21332
rect 37921 21295 37979 21301
rect 58158 21292 58164 21304
rect 58216 21292 58222 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 5718 21088 5724 21140
rect 5776 21128 5782 21140
rect 5905 21131 5963 21137
rect 5905 21128 5917 21131
rect 5776 21100 5917 21128
rect 5776 21088 5782 21100
rect 5905 21097 5917 21100
rect 5951 21128 5963 21131
rect 5994 21128 6000 21140
rect 5951 21100 6000 21128
rect 5951 21097 5963 21100
rect 5905 21091 5963 21097
rect 5994 21088 6000 21100
rect 6052 21088 6058 21140
rect 8202 21088 8208 21140
rect 8260 21128 8266 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 8260 21100 10149 21128
rect 8260 21088 8266 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 14645 21131 14703 21137
rect 14645 21128 14657 21131
rect 13136 21100 14657 21128
rect 13136 21088 13142 21100
rect 14645 21097 14657 21100
rect 14691 21128 14703 21131
rect 17954 21128 17960 21140
rect 14691 21100 17960 21128
rect 14691 21097 14703 21100
rect 14645 21091 14703 21097
rect 17954 21088 17960 21100
rect 18012 21088 18018 21140
rect 18874 21088 18880 21140
rect 18932 21128 18938 21140
rect 20162 21128 20168 21140
rect 18932 21100 20168 21128
rect 18932 21088 18938 21100
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 21177 21131 21235 21137
rect 21177 21128 21189 21131
rect 20400 21100 21189 21128
rect 10965 21063 11023 21069
rect 10965 21029 10977 21063
rect 11011 21060 11023 21063
rect 11146 21060 11152 21072
rect 11011 21032 11152 21060
rect 11011 21029 11023 21032
rect 10965 21023 11023 21029
rect 11146 21020 11152 21032
rect 11204 21020 11210 21072
rect 12250 21020 12256 21072
rect 12308 21060 12314 21072
rect 15933 21063 15991 21069
rect 15933 21060 15945 21063
rect 12308 21032 15945 21060
rect 12308 21020 12314 21032
rect 15933 21029 15945 21032
rect 15979 21029 15991 21063
rect 15933 21023 15991 21029
rect 17494 21020 17500 21072
rect 17552 21060 17558 21072
rect 19889 21063 19947 21069
rect 19889 21060 19901 21063
rect 17552 21032 19901 21060
rect 17552 21020 17558 21032
rect 19889 21029 19901 21032
rect 19935 21029 19947 21063
rect 20400 21060 20428 21100
rect 21177 21097 21189 21100
rect 21223 21128 21235 21131
rect 21358 21128 21364 21140
rect 21223 21100 21364 21128
rect 21223 21097 21235 21100
rect 21177 21091 21235 21097
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 21818 21128 21824 21140
rect 21779 21100 21824 21128
rect 21818 21088 21824 21100
rect 21876 21128 21882 21140
rect 21876 21100 22784 21128
rect 21876 21088 21882 21100
rect 20530 21060 20536 21072
rect 19889 21023 19947 21029
rect 20088 21032 20428 21060
rect 20457 21032 20536 21060
rect 13630 20952 13636 21004
rect 13688 20992 13694 21004
rect 20088 20992 20116 21032
rect 13688 20964 15424 20992
rect 13688 20952 13694 20964
rect 12897 20927 12955 20933
rect 12897 20893 12909 20927
rect 12943 20924 12955 20927
rect 13648 20924 13676 20952
rect 12943 20896 13676 20924
rect 12943 20893 12955 20896
rect 12897 20887 12955 20893
rect 14458 20884 14464 20936
rect 14516 20924 14522 20936
rect 14553 20927 14611 20933
rect 14553 20924 14565 20927
rect 14516 20896 14565 20924
rect 14516 20884 14522 20896
rect 14553 20893 14565 20896
rect 14599 20893 14611 20927
rect 15286 20924 15292 20936
rect 15247 20896 15292 20924
rect 14553 20887 14611 20893
rect 15286 20884 15292 20896
rect 15344 20884 15350 20936
rect 15396 20933 15424 20964
rect 19306 20964 20116 20992
rect 15382 20927 15440 20933
rect 15382 20893 15394 20927
rect 15428 20893 15440 20927
rect 15562 20924 15568 20936
rect 15523 20896 15568 20924
rect 15382 20887 15440 20893
rect 15562 20884 15568 20896
rect 15620 20884 15626 20936
rect 15795 20927 15853 20933
rect 15795 20893 15807 20927
rect 15841 20924 15853 20927
rect 16393 20927 16451 20933
rect 15841 20896 16344 20924
rect 15841 20893 15853 20896
rect 15795 20887 15853 20893
rect 2774 20816 2780 20868
rect 2832 20856 2838 20868
rect 2961 20859 3019 20865
rect 2961 20856 2973 20859
rect 2832 20828 2973 20856
rect 2832 20816 2838 20828
rect 2961 20825 2973 20828
rect 3007 20856 3019 20859
rect 4614 20856 4620 20868
rect 3007 20828 4620 20856
rect 3007 20825 3019 20828
rect 2961 20819 3019 20825
rect 4614 20816 4620 20828
rect 4672 20816 4678 20868
rect 6178 20856 6184 20868
rect 5644 20828 6184 20856
rect 5644 20800 5672 20828
rect 6178 20816 6184 20828
rect 6236 20816 6242 20868
rect 10413 20859 10471 20865
rect 10413 20825 10425 20859
rect 10459 20825 10471 20859
rect 10413 20819 10471 20825
rect 11149 20859 11207 20865
rect 11149 20825 11161 20859
rect 11195 20825 11207 20859
rect 12710 20856 12716 20868
rect 12671 20828 12716 20856
rect 11149 20819 11207 20825
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 4433 20791 4491 20797
rect 4433 20788 4445 20791
rect 3936 20760 4445 20788
rect 3936 20748 3942 20760
rect 4433 20757 4445 20760
rect 4479 20788 4491 20791
rect 5626 20788 5632 20800
rect 4479 20760 5632 20788
rect 4479 20757 4491 20760
rect 4433 20751 4491 20757
rect 5626 20748 5632 20760
rect 5684 20748 5690 20800
rect 6546 20748 6552 20800
rect 6604 20788 6610 20800
rect 6641 20791 6699 20797
rect 6641 20788 6653 20791
rect 6604 20760 6653 20788
rect 6604 20748 6610 20760
rect 6641 20757 6653 20760
rect 6687 20757 6699 20791
rect 6641 20751 6699 20757
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 9493 20791 9551 20797
rect 9493 20788 9505 20791
rect 8536 20760 9505 20788
rect 8536 20748 8542 20760
rect 9493 20757 9505 20760
rect 9539 20788 9551 20791
rect 10428 20788 10456 20819
rect 9539 20760 10456 20788
rect 11164 20788 11192 20819
rect 12710 20816 12716 20828
rect 12768 20816 12774 20868
rect 14476 20856 14504 20884
rect 12912 20828 14504 20856
rect 11606 20788 11612 20800
rect 11164 20760 11612 20788
rect 9539 20757 9551 20760
rect 9493 20751 9551 20757
rect 11606 20748 11612 20760
rect 11664 20788 11670 20800
rect 11701 20791 11759 20797
rect 11701 20788 11713 20791
rect 11664 20760 11713 20788
rect 11664 20748 11670 20760
rect 11701 20757 11713 20760
rect 11747 20788 11759 20791
rect 12912 20788 12940 20828
rect 15654 20816 15660 20868
rect 15712 20856 15718 20868
rect 15712 20828 15757 20856
rect 15712 20816 15718 20828
rect 11747 20760 12940 20788
rect 11747 20757 11759 20760
rect 11701 20751 11759 20757
rect 12986 20748 12992 20800
rect 13044 20788 13050 20800
rect 13081 20791 13139 20797
rect 13081 20788 13093 20791
rect 13044 20760 13093 20788
rect 13044 20748 13050 20760
rect 13081 20757 13093 20760
rect 13127 20757 13139 20791
rect 16316 20788 16344 20896
rect 16393 20893 16405 20927
rect 16439 20924 16451 20927
rect 17402 20924 17408 20936
rect 16439 20896 17408 20924
rect 16439 20893 16451 20896
rect 16393 20887 16451 20893
rect 17402 20884 17408 20896
rect 17460 20884 17466 20936
rect 16660 20859 16718 20865
rect 16660 20825 16672 20859
rect 16706 20856 16718 20859
rect 16758 20856 16764 20868
rect 16706 20828 16764 20856
rect 16706 20825 16718 20828
rect 16660 20819 16718 20825
rect 16758 20816 16764 20828
rect 16816 20816 16822 20868
rect 19306 20856 19334 20964
rect 20457 20933 20485 21032
rect 20530 21020 20536 21032
rect 20588 21020 20594 21072
rect 20068 20927 20126 20933
rect 20068 20924 20080 20927
rect 17604 20828 19334 20856
rect 19996 20896 20080 20924
rect 17604 20788 17632 20828
rect 17770 20788 17776 20800
rect 16316 20760 17632 20788
rect 17731 20760 17776 20788
rect 13081 20751 13139 20757
rect 17770 20748 17776 20760
rect 17828 20748 17834 20800
rect 19996 20788 20024 20896
rect 20068 20893 20080 20896
rect 20114 20893 20126 20927
rect 20068 20887 20126 20893
rect 20257 20927 20315 20933
rect 20257 20893 20269 20927
rect 20303 20893 20315 20927
rect 20257 20887 20315 20893
rect 20440 20927 20498 20933
rect 20440 20893 20452 20927
rect 20486 20893 20498 20927
rect 20440 20887 20498 20893
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20924 20591 20927
rect 20990 20924 20996 20936
rect 20579 20896 20996 20924
rect 20579 20893 20591 20896
rect 20533 20887 20591 20893
rect 20162 20856 20168 20868
rect 20123 20828 20168 20856
rect 20162 20816 20168 20828
rect 20220 20816 20226 20868
rect 20272 20856 20300 20887
rect 20990 20884 20996 20896
rect 21048 20884 21054 20936
rect 22094 20884 22100 20936
rect 22152 20924 22158 20936
rect 22373 20927 22431 20933
rect 22373 20924 22385 20927
rect 22152 20896 22385 20924
rect 22152 20884 22158 20896
rect 22373 20893 22385 20896
rect 22419 20893 22431 20927
rect 22554 20924 22560 20936
rect 22515 20896 22560 20924
rect 22373 20887 22431 20893
rect 22554 20884 22560 20896
rect 22612 20884 22618 20936
rect 22756 20933 22784 21100
rect 22830 21088 22836 21140
rect 22888 21088 22894 21140
rect 23017 21131 23075 21137
rect 23017 21097 23029 21131
rect 23063 21128 23075 21131
rect 23106 21128 23112 21140
rect 23063 21100 23112 21128
rect 23063 21097 23075 21100
rect 23017 21091 23075 21097
rect 23106 21088 23112 21100
rect 23164 21088 23170 21140
rect 27706 21088 27712 21140
rect 27764 21128 27770 21140
rect 32950 21128 32956 21140
rect 27764 21100 32956 21128
rect 27764 21088 27770 21100
rect 32950 21088 32956 21100
rect 33008 21088 33014 21140
rect 22848 21060 22876 21088
rect 23477 21063 23535 21069
rect 23477 21060 23489 21063
rect 22848 21032 23489 21060
rect 23477 21029 23489 21032
rect 23523 21029 23535 21063
rect 23477 21023 23535 21029
rect 30190 20952 30196 21004
rect 30248 20952 30254 21004
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 22741 20927 22799 20933
rect 22741 20893 22753 20927
rect 22787 20893 22799 20927
rect 22741 20887 22799 20893
rect 20622 20856 20628 20868
rect 20272 20828 20628 20856
rect 20622 20816 20628 20828
rect 20680 20816 20686 20868
rect 21082 20856 21088 20868
rect 21043 20828 21088 20856
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 22664 20856 22692 20887
rect 23014 20884 23020 20936
rect 23072 20924 23078 20936
rect 28997 20927 29055 20933
rect 23072 20896 27476 20924
rect 23072 20884 23078 20896
rect 27448 20868 27476 20896
rect 28997 20893 29009 20927
rect 29043 20924 29055 20927
rect 29270 20924 29276 20936
rect 29043 20896 29276 20924
rect 29043 20893 29055 20896
rect 28997 20887 29055 20893
rect 29270 20884 29276 20896
rect 29328 20924 29334 20936
rect 30009 20927 30067 20933
rect 30009 20924 30021 20927
rect 29328 20896 30021 20924
rect 29328 20884 29334 20896
rect 30009 20893 30021 20896
rect 30055 20924 30067 20927
rect 30208 20924 30236 20952
rect 30055 20896 30236 20924
rect 30055 20893 30067 20896
rect 30009 20887 30067 20893
rect 40218 20884 40224 20936
rect 40276 20924 40282 20936
rect 40589 20927 40647 20933
rect 40589 20924 40601 20927
rect 40276 20896 40601 20924
rect 40276 20884 40282 20896
rect 40589 20893 40601 20896
rect 40635 20893 40647 20927
rect 40589 20887 40647 20893
rect 22922 20856 22928 20868
rect 22664 20828 22928 20856
rect 22922 20816 22928 20828
rect 22980 20816 22986 20868
rect 23661 20859 23719 20865
rect 23661 20825 23673 20859
rect 23707 20825 23719 20859
rect 23661 20819 23719 20825
rect 23845 20859 23903 20865
rect 23845 20825 23857 20859
rect 23891 20856 23903 20859
rect 23934 20856 23940 20868
rect 23891 20828 23940 20856
rect 23891 20825 23903 20828
rect 23845 20819 23903 20825
rect 20254 20788 20260 20800
rect 19996 20760 20260 20788
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 23676 20788 23704 20819
rect 23934 20816 23940 20828
rect 23992 20856 23998 20868
rect 25038 20856 25044 20868
rect 23992 20828 25044 20856
rect 23992 20816 23998 20828
rect 25038 20816 25044 20828
rect 25096 20816 25102 20868
rect 25685 20859 25743 20865
rect 25685 20825 25697 20859
rect 25731 20825 25743 20859
rect 27430 20856 27436 20868
rect 27391 20828 27436 20856
rect 25685 20819 25743 20825
rect 24394 20788 24400 20800
rect 23676 20760 24400 20788
rect 24394 20748 24400 20760
rect 24452 20748 24458 20800
rect 25700 20788 25728 20819
rect 27430 20816 27436 20828
rect 27488 20816 27494 20868
rect 30193 20859 30251 20865
rect 30193 20825 30205 20859
rect 30239 20856 30251 20859
rect 30834 20856 30840 20868
rect 30239 20828 30840 20856
rect 30239 20825 30251 20828
rect 30193 20819 30251 20825
rect 30834 20816 30840 20828
rect 30892 20816 30898 20868
rect 40405 20859 40463 20865
rect 40405 20825 40417 20859
rect 40451 20856 40463 20859
rect 40494 20856 40500 20868
rect 40451 20828 40500 20856
rect 40451 20825 40463 20828
rect 40405 20819 40463 20825
rect 40494 20816 40500 20828
rect 40552 20816 40558 20868
rect 40678 20816 40684 20868
rect 40736 20856 40742 20868
rect 41233 20859 41291 20865
rect 41233 20856 41245 20859
rect 40736 20828 41245 20856
rect 40736 20816 40742 20828
rect 41233 20825 41245 20828
rect 41279 20825 41291 20859
rect 41233 20819 41291 20825
rect 27706 20788 27712 20800
rect 25700 20760 27712 20788
rect 27706 20748 27712 20760
rect 27764 20748 27770 20800
rect 28166 20748 28172 20800
rect 28224 20788 28230 20800
rect 28445 20791 28503 20797
rect 28445 20788 28457 20791
rect 28224 20760 28457 20788
rect 28224 20748 28230 20760
rect 28445 20757 28457 20760
rect 28491 20788 28503 20791
rect 28534 20788 28540 20800
rect 28491 20760 28540 20788
rect 28491 20757 28503 20760
rect 28445 20751 28503 20757
rect 28534 20748 28540 20760
rect 28592 20748 28598 20800
rect 37458 20788 37464 20800
rect 37419 20760 37464 20788
rect 37458 20748 37464 20760
rect 37516 20748 37522 20800
rect 40773 20791 40831 20797
rect 40773 20757 40785 20791
rect 40819 20788 40831 20791
rect 41138 20788 41144 20800
rect 40819 20760 41144 20788
rect 40819 20757 40831 20760
rect 40773 20751 40831 20757
rect 41138 20748 41144 20760
rect 41196 20748 41202 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 7101 20587 7159 20593
rect 7101 20553 7113 20587
rect 7147 20584 7159 20587
rect 8021 20587 8079 20593
rect 7147 20556 7181 20584
rect 7147 20553 7159 20556
rect 7101 20547 7159 20553
rect 8021 20553 8033 20587
rect 8067 20584 8079 20587
rect 8386 20584 8392 20596
rect 8067 20556 8392 20584
rect 8067 20553 8079 20556
rect 8021 20547 8079 20553
rect 5810 20476 5816 20528
rect 5868 20516 5874 20528
rect 7116 20516 7144 20547
rect 8386 20544 8392 20556
rect 8444 20584 8450 20596
rect 12526 20584 12532 20596
rect 8444 20556 12532 20584
rect 8444 20544 8450 20556
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 13630 20584 13636 20596
rect 13591 20556 13636 20584
rect 13630 20544 13636 20556
rect 13688 20544 13694 20596
rect 17129 20587 17187 20593
rect 17129 20553 17141 20587
rect 17175 20584 17187 20587
rect 17218 20584 17224 20596
rect 17175 20556 17224 20584
rect 17175 20553 17187 20556
rect 17129 20547 17187 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 19444 20556 19784 20584
rect 11514 20516 11520 20528
rect 5868 20488 11520 20516
rect 5868 20476 5874 20488
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 17313 20519 17371 20525
rect 17313 20485 17325 20519
rect 17359 20516 17371 20519
rect 17770 20516 17776 20528
rect 17359 20488 17776 20516
rect 17359 20485 17371 20488
rect 17313 20479 17371 20485
rect 17770 20476 17776 20488
rect 17828 20516 17834 20528
rect 19444 20516 19472 20556
rect 17828 20488 19371 20516
rect 17828 20476 17834 20488
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 12526 20457 12532 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 6604 20420 7205 20448
rect 6604 20408 6610 20420
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 8113 20451 8171 20457
rect 8113 20417 8125 20451
rect 8159 20417 8171 20451
rect 8113 20411 8171 20417
rect 12520 20411 12532 20457
rect 12584 20448 12590 20460
rect 12584 20420 12620 20448
rect 4985 20383 5043 20389
rect 4985 20349 4997 20383
rect 5031 20380 5043 20383
rect 6822 20380 6828 20392
rect 5031 20352 6828 20380
rect 5031 20349 5043 20352
rect 4985 20343 5043 20349
rect 6822 20340 6828 20352
rect 6880 20380 6886 20392
rect 8128 20380 8156 20411
rect 12526 20408 12532 20411
rect 12584 20408 12590 20420
rect 12802 20408 12808 20460
rect 12860 20448 12866 20460
rect 14369 20451 14427 20457
rect 14369 20448 14381 20451
rect 12860 20420 14381 20448
rect 12860 20408 12866 20420
rect 14369 20417 14381 20420
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 15286 20408 15292 20460
rect 15344 20448 15350 20460
rect 15657 20451 15715 20457
rect 15657 20448 15669 20451
rect 15344 20420 15669 20448
rect 15344 20408 15350 20420
rect 15657 20417 15669 20420
rect 15703 20448 15715 20451
rect 15746 20448 15752 20460
rect 15703 20420 15752 20448
rect 15703 20417 15715 20420
rect 15657 20411 15715 20417
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16574 20448 16580 20460
rect 15887 20420 16580 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16574 20408 16580 20420
rect 16632 20448 16638 20460
rect 17497 20451 17555 20457
rect 17497 20448 17509 20451
rect 16632 20420 17509 20448
rect 16632 20408 16638 20420
rect 17497 20417 17509 20420
rect 17543 20448 17555 20451
rect 17586 20448 17592 20460
rect 17543 20420 17592 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 17586 20408 17592 20420
rect 17644 20408 17650 20460
rect 18325 20451 18383 20457
rect 18325 20417 18337 20451
rect 18371 20448 18383 20451
rect 18371 20420 19288 20448
rect 18371 20417 18383 20420
rect 18325 20411 18383 20417
rect 6880 20352 8156 20380
rect 12253 20383 12311 20389
rect 6880 20340 6886 20352
rect 12253 20349 12265 20383
rect 12299 20349 12311 20383
rect 14090 20380 14096 20392
rect 14051 20352 14096 20380
rect 12253 20343 12311 20349
rect 12268 20244 12296 20343
rect 14090 20340 14096 20352
rect 14148 20340 14154 20392
rect 15473 20383 15531 20389
rect 15473 20349 15485 20383
rect 15519 20380 15531 20383
rect 15930 20380 15936 20392
rect 15519 20352 15936 20380
rect 15519 20349 15531 20352
rect 15473 20343 15531 20349
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 18233 20383 18291 20389
rect 18233 20349 18245 20383
rect 18279 20349 18291 20383
rect 18233 20343 18291 20349
rect 14108 20312 14136 20340
rect 16942 20312 16948 20324
rect 14108 20284 16948 20312
rect 16942 20272 16948 20284
rect 17000 20272 17006 20324
rect 12434 20244 12440 20256
rect 12268 20216 12440 20244
rect 12434 20204 12440 20216
rect 12492 20204 12498 20256
rect 17954 20244 17960 20256
rect 17915 20216 17960 20244
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 18138 20244 18144 20256
rect 18099 20216 18144 20244
rect 18138 20204 18144 20216
rect 18196 20204 18202 20256
rect 18248 20244 18276 20343
rect 19260 20321 19288 20420
rect 19343 20380 19371 20488
rect 19439 20488 19472 20516
rect 19439 20457 19467 20488
rect 19610 20476 19616 20528
rect 19668 20516 19674 20528
rect 19756 20516 19784 20556
rect 20162 20544 20168 20596
rect 20220 20584 20226 20596
rect 27525 20587 27583 20593
rect 20220 20556 26188 20584
rect 20220 20544 20226 20556
rect 20254 20516 20260 20528
rect 19668 20488 19713 20516
rect 19756 20488 20260 20516
rect 19668 20476 19674 20488
rect 20254 20476 20260 20488
rect 20312 20476 20318 20528
rect 20530 20516 20536 20528
rect 20457 20488 20536 20516
rect 19424 20451 19482 20457
rect 19424 20417 19436 20451
rect 19470 20417 19482 20451
rect 19424 20411 19482 20417
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19794 20448 19800 20460
rect 19576 20420 19621 20448
rect 19755 20420 19800 20448
rect 19576 20408 19582 20420
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 20070 20448 20076 20460
rect 19935 20420 20076 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20346 20448 20352 20460
rect 20307 20420 20352 20448
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20457 20457 20485 20488
rect 20530 20476 20536 20488
rect 20588 20476 20594 20528
rect 20714 20516 20720 20528
rect 20675 20488 20720 20516
rect 20714 20476 20720 20488
rect 20772 20476 20778 20528
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 26160 20516 26188 20556
rect 27525 20553 27537 20587
rect 27571 20584 27583 20587
rect 27798 20584 27804 20596
rect 27571 20556 27804 20584
rect 27571 20553 27583 20556
rect 27525 20547 27583 20553
rect 27798 20544 27804 20556
rect 27856 20544 27862 20596
rect 28721 20587 28779 20593
rect 28721 20553 28733 20587
rect 28767 20584 28779 20587
rect 28810 20584 28816 20596
rect 28767 20556 28816 20584
rect 28767 20553 28779 20556
rect 28721 20547 28779 20553
rect 28810 20544 28816 20556
rect 28868 20584 28874 20596
rect 29546 20584 29552 20596
rect 28868 20556 29552 20584
rect 28868 20544 28874 20556
rect 29546 20544 29552 20556
rect 29604 20544 29610 20596
rect 29822 20584 29828 20596
rect 29783 20556 29828 20584
rect 29822 20544 29828 20556
rect 29880 20544 29886 20596
rect 30285 20587 30343 20593
rect 30285 20553 30297 20587
rect 30331 20553 30343 20587
rect 37274 20584 37280 20596
rect 30285 20547 30343 20553
rect 31726 20556 37105 20584
rect 37235 20556 37280 20584
rect 30300 20516 30328 20547
rect 30742 20516 30748 20528
rect 22152 20488 22197 20516
rect 26160 20488 30328 20516
rect 30703 20488 30748 20516
rect 22152 20476 22158 20488
rect 30742 20476 30748 20488
rect 30800 20476 30806 20528
rect 20442 20451 20500 20457
rect 20442 20417 20454 20451
rect 20488 20417 20500 20451
rect 20622 20448 20628 20460
rect 20583 20420 20628 20448
rect 20442 20411 20500 20417
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 20814 20451 20872 20457
rect 20814 20417 20826 20451
rect 20860 20448 20872 20451
rect 21082 20448 21088 20460
rect 20860 20420 21088 20448
rect 20860 20417 20872 20420
rect 20814 20411 20872 20417
rect 19343 20352 19467 20380
rect 19439 20324 19467 20352
rect 20254 20340 20260 20392
rect 20312 20380 20318 20392
rect 20829 20380 20857 20411
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 23014 20448 23020 20460
rect 22975 20420 23020 20448
rect 23014 20408 23020 20420
rect 23072 20408 23078 20460
rect 23290 20457 23296 20460
rect 23284 20448 23296 20457
rect 23251 20420 23296 20448
rect 23284 20411 23296 20420
rect 23290 20408 23296 20411
rect 23348 20408 23354 20460
rect 25774 20408 25780 20460
rect 25832 20448 25838 20460
rect 26154 20451 26212 20457
rect 26154 20448 26166 20451
rect 25832 20420 26166 20448
rect 25832 20408 25838 20420
rect 26154 20417 26166 20420
rect 26200 20417 26212 20451
rect 26154 20411 26212 20417
rect 27433 20451 27491 20457
rect 27433 20417 27445 20451
rect 27479 20448 27491 20451
rect 27522 20448 27528 20460
rect 27479 20420 27528 20448
rect 27479 20417 27491 20420
rect 27433 20411 27491 20417
rect 27522 20408 27528 20420
rect 27580 20448 27586 20460
rect 27890 20448 27896 20460
rect 27580 20420 27896 20448
rect 27580 20408 27586 20420
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 28534 20408 28540 20460
rect 28592 20448 28598 20460
rect 28629 20451 28687 20457
rect 28629 20448 28641 20451
rect 28592 20420 28641 20448
rect 28592 20408 28598 20420
rect 28629 20417 28641 20420
rect 28675 20417 28687 20451
rect 28629 20411 28687 20417
rect 28994 20408 29000 20460
rect 29052 20448 29058 20460
rect 29273 20451 29331 20457
rect 29273 20448 29285 20451
rect 29052 20420 29285 20448
rect 29052 20408 29058 20420
rect 29273 20417 29285 20420
rect 29319 20417 29331 20451
rect 29454 20448 29460 20460
rect 29415 20420 29460 20448
rect 29273 20411 29331 20417
rect 29454 20408 29460 20420
rect 29512 20408 29518 20460
rect 29549 20451 29607 20457
rect 29549 20417 29561 20451
rect 29595 20417 29607 20451
rect 29549 20411 29607 20417
rect 20312 20352 20857 20380
rect 26421 20383 26479 20389
rect 20312 20340 20318 20352
rect 26421 20349 26433 20383
rect 26467 20349 26479 20383
rect 26421 20343 26479 20349
rect 19245 20315 19303 20321
rect 19245 20281 19257 20315
rect 19291 20281 19303 20315
rect 19245 20275 19303 20281
rect 19426 20272 19432 20324
rect 19484 20272 19490 20324
rect 19518 20272 19524 20324
rect 19576 20312 19582 20324
rect 25041 20315 25099 20321
rect 25041 20312 25053 20315
rect 19576 20284 23060 20312
rect 19576 20272 19582 20284
rect 20162 20244 20168 20256
rect 18248 20216 20168 20244
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20990 20244 20996 20256
rect 20951 20216 20996 20244
rect 20990 20204 20996 20216
rect 21048 20204 21054 20256
rect 23032 20244 23060 20284
rect 23952 20284 25053 20312
rect 23952 20244 23980 20284
rect 25041 20281 25053 20284
rect 25087 20281 25099 20315
rect 26436 20312 26464 20343
rect 27430 20312 27436 20324
rect 26436 20284 27436 20312
rect 25041 20275 25099 20281
rect 24394 20244 24400 20256
rect 23032 20216 23980 20244
rect 24355 20216 24400 20244
rect 24394 20204 24400 20216
rect 24452 20204 24458 20256
rect 25056 20244 25084 20275
rect 27430 20272 27436 20284
rect 27488 20272 27494 20324
rect 29564 20312 29592 20411
rect 29638 20408 29644 20460
rect 29696 20448 29702 20460
rect 30469 20451 30527 20457
rect 29696 20420 29741 20448
rect 29696 20408 29702 20420
rect 30469 20417 30481 20451
rect 30515 20448 30527 20451
rect 31726 20448 31754 20556
rect 33134 20516 33140 20528
rect 32876 20488 33140 20516
rect 32582 20448 32588 20460
rect 30515 20420 31754 20448
rect 32543 20420 32588 20448
rect 30515 20417 30527 20420
rect 30469 20411 30527 20417
rect 32582 20408 32588 20420
rect 32640 20408 32646 20460
rect 32766 20448 32772 20460
rect 32727 20420 32772 20448
rect 32766 20408 32772 20420
rect 32824 20408 32830 20460
rect 32876 20457 32904 20488
rect 33134 20476 33140 20488
rect 33192 20476 33198 20528
rect 33229 20519 33287 20525
rect 33229 20485 33241 20519
rect 33275 20516 33287 20519
rect 34802 20519 34860 20525
rect 34802 20516 34814 20519
rect 33275 20488 34814 20516
rect 33275 20485 33287 20488
rect 33229 20479 33287 20485
rect 34802 20485 34814 20488
rect 34848 20485 34860 20519
rect 37077 20516 37105 20556
rect 37274 20544 37280 20556
rect 37332 20544 37338 20596
rect 40954 20584 40960 20596
rect 40788 20556 40960 20584
rect 37366 20516 37372 20528
rect 37077 20488 37372 20516
rect 34802 20479 34860 20485
rect 37366 20476 37372 20488
rect 37424 20476 37430 20528
rect 37642 20516 37648 20528
rect 37603 20488 37648 20516
rect 37642 20476 37648 20488
rect 37700 20476 37706 20528
rect 39108 20519 39166 20525
rect 39108 20485 39120 20519
rect 39154 20516 39166 20519
rect 40681 20519 40739 20525
rect 40681 20516 40693 20519
rect 39154 20488 40693 20516
rect 39154 20485 39166 20488
rect 39108 20479 39166 20485
rect 40681 20485 40693 20488
rect 40727 20485 40739 20519
rect 40681 20479 40739 20485
rect 32864 20451 32922 20457
rect 32864 20417 32876 20451
rect 32910 20417 32922 20451
rect 32864 20411 32922 20417
rect 32950 20408 32956 20460
rect 33008 20448 33014 20460
rect 33008 20420 33053 20448
rect 33008 20408 33014 20420
rect 37274 20408 37280 20460
rect 37332 20448 37338 20460
rect 37461 20451 37519 20457
rect 37461 20448 37473 20451
rect 37332 20420 37473 20448
rect 37332 20408 37338 20420
rect 37461 20417 37473 20420
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 37550 20408 37556 20460
rect 37608 20448 37614 20460
rect 37826 20448 37832 20460
rect 37608 20420 37653 20448
rect 37787 20420 37832 20448
rect 37608 20408 37614 20420
rect 37826 20408 37832 20420
rect 37884 20408 37890 20460
rect 30558 20380 30564 20392
rect 30519 20352 30564 20380
rect 30558 20340 30564 20352
rect 30616 20340 30622 20392
rect 35069 20383 35127 20389
rect 35069 20349 35081 20383
rect 35115 20380 35127 20383
rect 38746 20380 38752 20392
rect 35115 20352 38752 20380
rect 35115 20349 35127 20352
rect 35069 20343 35127 20349
rect 32766 20312 32772 20324
rect 29564 20284 32772 20312
rect 32766 20272 32772 20284
rect 32824 20272 32830 20324
rect 27062 20244 27068 20256
rect 25056 20216 27068 20244
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 30466 20244 30472 20256
rect 30427 20216 30472 20244
rect 30466 20204 30472 20216
rect 30524 20204 30530 20256
rect 33134 20204 33140 20256
rect 33192 20244 33198 20256
rect 33689 20247 33747 20253
rect 33689 20244 33701 20247
rect 33192 20216 33701 20244
rect 33192 20204 33198 20216
rect 33689 20213 33701 20216
rect 33735 20213 33747 20247
rect 33689 20207 33747 20213
rect 34146 20204 34152 20256
rect 34204 20244 34210 20256
rect 35084 20244 35112 20343
rect 38746 20340 38752 20352
rect 38804 20380 38810 20392
rect 38841 20383 38899 20389
rect 38841 20380 38853 20383
rect 38804 20352 38853 20380
rect 38804 20340 38810 20352
rect 38841 20349 38853 20352
rect 38887 20349 38899 20383
rect 38841 20343 38899 20349
rect 40494 20272 40500 20324
rect 40552 20312 40558 20324
rect 40788 20312 40816 20556
rect 40954 20544 40960 20556
rect 41012 20544 41018 20596
rect 40951 20457 40957 20460
rect 40911 20451 40957 20457
rect 40911 20417 40923 20451
rect 40911 20411 40957 20417
rect 40951 20408 40957 20411
rect 41009 20408 41015 20460
rect 41046 20451 41104 20457
rect 41046 20417 41058 20451
rect 41092 20417 41104 20451
rect 41046 20411 41104 20417
rect 41146 20451 41204 20457
rect 41146 20417 41158 20451
rect 41192 20417 41204 20451
rect 41146 20411 41204 20417
rect 41325 20451 41383 20457
rect 41325 20417 41337 20451
rect 41371 20417 41383 20451
rect 41325 20411 41383 20417
rect 41064 20380 41092 20411
rect 40969 20352 41092 20380
rect 41156 20380 41184 20411
rect 41230 20380 41236 20392
rect 41156 20352 41236 20380
rect 40969 20312 40997 20352
rect 41230 20340 41236 20352
rect 41288 20340 41294 20392
rect 40552 20284 40997 20312
rect 40552 20272 40558 20284
rect 41046 20272 41052 20324
rect 41104 20312 41110 20324
rect 41340 20312 41368 20411
rect 41104 20284 41368 20312
rect 41104 20272 41110 20284
rect 40218 20244 40224 20256
rect 34204 20216 35112 20244
rect 40179 20216 40224 20244
rect 34204 20204 34210 20216
rect 40218 20204 40224 20216
rect 40276 20204 40282 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 6270 20000 6276 20052
rect 6328 20040 6334 20052
rect 6365 20043 6423 20049
rect 6365 20040 6377 20043
rect 6328 20012 6377 20040
rect 6328 20000 6334 20012
rect 6365 20009 6377 20012
rect 6411 20009 6423 20043
rect 6365 20003 6423 20009
rect 8846 20000 8852 20052
rect 8904 20040 8910 20052
rect 9125 20043 9183 20049
rect 9125 20040 9137 20043
rect 8904 20012 9137 20040
rect 8904 20000 8910 20012
rect 9125 20009 9137 20012
rect 9171 20009 9183 20043
rect 9125 20003 9183 20009
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 11333 20043 11391 20049
rect 11333 20040 11345 20043
rect 11204 20012 11345 20040
rect 11204 20000 11210 20012
rect 11333 20009 11345 20012
rect 11379 20009 11391 20043
rect 11333 20003 11391 20009
rect 12437 20043 12495 20049
rect 12437 20009 12449 20043
rect 12483 20040 12495 20043
rect 12526 20040 12532 20052
rect 12483 20012 12532 20040
rect 12483 20009 12495 20012
rect 12437 20003 12495 20009
rect 12526 20000 12532 20012
rect 12584 20000 12590 20052
rect 15194 20040 15200 20052
rect 15155 20012 15200 20040
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15746 20000 15752 20052
rect 15804 20040 15810 20052
rect 19610 20040 19616 20052
rect 15804 20012 19616 20040
rect 15804 20000 15810 20012
rect 19610 20000 19616 20012
rect 19668 20040 19674 20052
rect 20622 20040 20628 20052
rect 19668 20012 20628 20040
rect 19668 20000 19674 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 21821 20043 21879 20049
rect 21821 20009 21833 20043
rect 21867 20040 21879 20043
rect 22094 20040 22100 20052
rect 21867 20012 22100 20040
rect 21867 20009 21879 20012
rect 21821 20003 21879 20009
rect 22094 20000 22100 20012
rect 22152 20040 22158 20052
rect 22922 20040 22928 20052
rect 22152 20012 22928 20040
rect 22152 20000 22158 20012
rect 22922 20000 22928 20012
rect 22980 20000 22986 20052
rect 25774 20040 25780 20052
rect 25735 20012 25780 20040
rect 25774 20000 25780 20012
rect 25832 20000 25838 20052
rect 27706 20040 27712 20052
rect 27667 20012 27712 20040
rect 27706 20000 27712 20012
rect 27764 20000 27770 20052
rect 28997 20043 29055 20049
rect 28997 20009 29009 20043
rect 29043 20040 29055 20043
rect 30466 20040 30472 20052
rect 29043 20012 30472 20040
rect 29043 20009 29055 20012
rect 28997 20003 29055 20009
rect 30466 20000 30472 20012
rect 30524 20000 30530 20052
rect 32858 20000 32864 20052
rect 32916 20040 32922 20052
rect 32953 20043 33011 20049
rect 32953 20040 32965 20043
rect 32916 20012 32965 20040
rect 32916 20000 32922 20012
rect 32953 20009 32965 20012
rect 32999 20009 33011 20043
rect 32953 20003 33011 20009
rect 38654 20000 38660 20052
rect 38712 20040 38718 20052
rect 41417 20043 41475 20049
rect 41417 20040 41429 20043
rect 38712 20012 41429 20040
rect 38712 20000 38718 20012
rect 12802 19932 12808 19984
rect 12860 19932 12866 19984
rect 16574 19972 16580 19984
rect 14476 19944 16580 19972
rect 4614 19904 4620 19916
rect 4527 19876 4620 19904
rect 4614 19864 4620 19876
rect 4672 19904 4678 19916
rect 5442 19904 5448 19916
rect 4672 19876 5448 19904
rect 4672 19864 4678 19876
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 2498 19836 2504 19848
rect 2459 19808 2504 19836
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 6546 19836 6552 19848
rect 5092 19808 6552 19836
rect 5092 19780 5120 19808
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19836 9367 19839
rect 12250 19836 12256 19848
rect 9355 19808 12256 19836
rect 9355 19805 9367 19808
rect 9309 19799 9367 19805
rect 3881 19771 3939 19777
rect 3881 19737 3893 19771
rect 3927 19768 3939 19771
rect 4433 19771 4491 19777
rect 4433 19768 4445 19771
rect 3927 19740 4445 19768
rect 3927 19737 3939 19740
rect 3881 19731 3939 19737
rect 4433 19737 4445 19740
rect 4479 19768 4491 19771
rect 5074 19768 5080 19780
rect 4479 19740 5080 19768
rect 4479 19737 4491 19740
rect 4433 19731 4491 19737
rect 5074 19728 5080 19740
rect 5132 19728 5138 19780
rect 5350 19728 5356 19780
rect 5408 19768 5414 19780
rect 5813 19771 5871 19777
rect 5813 19768 5825 19771
rect 5408 19740 5825 19768
rect 5408 19728 5414 19740
rect 5813 19737 5825 19740
rect 5859 19768 5871 19771
rect 6641 19771 6699 19777
rect 6641 19768 6653 19771
rect 5859 19740 6653 19768
rect 5859 19737 5871 19740
rect 5813 19731 5871 19737
rect 6641 19737 6653 19740
rect 6687 19737 6699 19771
rect 9232 19768 9260 19799
rect 12250 19796 12256 19808
rect 12308 19796 12314 19848
rect 12817 19845 12845 19932
rect 12667 19839 12725 19845
rect 12667 19836 12679 19839
rect 12544 19808 12679 19836
rect 9858 19768 9864 19780
rect 9232 19740 9864 19768
rect 6641 19731 6699 19737
rect 9858 19728 9864 19740
rect 9916 19728 9922 19780
rect 12544 19712 12572 19808
rect 12667 19805 12679 19808
rect 12713 19805 12725 19839
rect 12667 19799 12725 19805
rect 12802 19839 12860 19845
rect 12802 19805 12814 19839
rect 12848 19805 12860 19839
rect 12802 19799 12860 19805
rect 12897 19839 12955 19845
rect 12897 19805 12909 19839
rect 12943 19836 12955 19839
rect 12986 19836 12992 19848
rect 12943 19808 12992 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 13078 19796 13084 19848
rect 13136 19836 13142 19848
rect 14476 19845 14504 19944
rect 16574 19932 16580 19944
rect 16632 19932 16638 19984
rect 28258 19972 28264 19984
rect 26157 19944 28264 19972
rect 15194 19904 15200 19916
rect 15155 19876 15200 19904
rect 15194 19864 15200 19876
rect 15252 19864 15258 19916
rect 22373 19907 22431 19913
rect 22373 19904 22385 19907
rect 21744 19876 22385 19904
rect 14461 19839 14519 19845
rect 13136 19808 13181 19836
rect 13136 19796 13142 19808
rect 14461 19805 14473 19839
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19836 15347 19839
rect 17494 19836 17500 19848
rect 15335 19808 17500 19836
rect 15335 19805 15347 19808
rect 15289 19799 15347 19805
rect 17494 19796 17500 19808
rect 17552 19796 17558 19848
rect 21744 19845 21772 19876
rect 22373 19873 22385 19876
rect 22419 19873 22431 19907
rect 22373 19867 22431 19873
rect 21729 19839 21787 19845
rect 21729 19836 21741 19839
rect 19996 19808 21741 19836
rect 19996 19780 20024 19808
rect 21729 19805 21741 19808
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 21913 19839 21971 19845
rect 21913 19805 21925 19839
rect 21959 19836 21971 19839
rect 22186 19836 22192 19848
rect 21959 19808 22192 19836
rect 21959 19805 21971 19808
rect 21913 19799 21971 19805
rect 22186 19796 22192 19808
rect 22244 19796 22250 19848
rect 26050 19836 26056 19848
rect 26011 19808 26056 19836
rect 26050 19796 26056 19808
rect 26108 19796 26114 19848
rect 26157 19845 26185 19944
rect 28258 19932 28264 19944
rect 28316 19932 28322 19984
rect 26881 19907 26939 19913
rect 26881 19904 26893 19907
rect 26344 19876 26893 19904
rect 26142 19839 26200 19845
rect 26142 19805 26154 19839
rect 26188 19805 26200 19839
rect 26142 19799 26200 19805
rect 26237 19839 26295 19845
rect 26237 19805 26249 19839
rect 26283 19836 26295 19839
rect 26283 19805 26301 19836
rect 26237 19799 26301 19805
rect 14182 19728 14188 19780
rect 14240 19768 14246 19780
rect 19978 19768 19984 19780
rect 14240 19740 19984 19768
rect 14240 19728 14246 19740
rect 19978 19728 19984 19740
rect 20036 19728 20042 19780
rect 24578 19728 24584 19780
rect 24636 19768 24642 19780
rect 26151 19768 26179 19799
rect 24636 19740 26179 19768
rect 26273 19768 26301 19799
rect 26344 19768 26372 19876
rect 26881 19873 26893 19876
rect 26927 19873 26939 19907
rect 28626 19904 28632 19916
rect 26881 19867 26939 19873
rect 27264 19876 28632 19904
rect 26421 19839 26479 19845
rect 26421 19805 26433 19839
rect 26467 19836 26479 19839
rect 26510 19836 26516 19848
rect 26467 19808 26516 19836
rect 26467 19805 26479 19808
rect 26421 19799 26479 19805
rect 26510 19796 26516 19808
rect 26568 19796 26574 19848
rect 27062 19836 27068 19848
rect 27023 19808 27068 19836
rect 27062 19796 27068 19808
rect 27120 19796 27126 19848
rect 26273 19740 26372 19768
rect 24636 19728 24642 19740
rect 26878 19728 26884 19780
rect 26936 19768 26942 19780
rect 27264 19777 27292 19876
rect 28626 19864 28632 19876
rect 28684 19864 28690 19916
rect 36262 19904 36268 19916
rect 36223 19876 36268 19904
rect 36262 19864 36268 19876
rect 36320 19864 36326 19916
rect 27614 19796 27620 19848
rect 27672 19836 27678 19848
rect 28445 19839 28503 19845
rect 28445 19836 28457 19839
rect 27672 19808 28457 19836
rect 27672 19796 27678 19808
rect 28445 19805 28457 19808
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19836 28871 19839
rect 28902 19836 28908 19848
rect 28859 19808 28908 19836
rect 28859 19805 28871 19808
rect 28813 19799 28871 19805
rect 28902 19796 28908 19808
rect 28960 19836 28966 19848
rect 29638 19836 29644 19848
rect 28960 19808 29644 19836
rect 28960 19796 28966 19808
rect 29638 19796 29644 19808
rect 29696 19836 29702 19848
rect 29825 19839 29883 19845
rect 29825 19836 29837 19839
rect 29696 19808 29837 19836
rect 29696 19796 29702 19808
rect 29825 19805 29837 19808
rect 29871 19805 29883 19839
rect 29825 19799 29883 19805
rect 30006 19796 30012 19848
rect 30064 19836 30070 19848
rect 30101 19839 30159 19845
rect 30101 19836 30113 19839
rect 30064 19808 30113 19836
rect 30064 19796 30070 19808
rect 30101 19805 30113 19808
rect 30147 19836 30159 19839
rect 31386 19836 31392 19848
rect 30147 19808 31392 19836
rect 30147 19805 30159 19808
rect 30101 19799 30159 19805
rect 31386 19796 31392 19808
rect 31444 19796 31450 19848
rect 32766 19796 32772 19848
rect 32824 19836 32830 19848
rect 33134 19836 33140 19848
rect 32824 19808 33140 19836
rect 32824 19796 32830 19808
rect 33134 19796 33140 19808
rect 33192 19796 33198 19848
rect 33318 19836 33324 19848
rect 33279 19808 33324 19836
rect 33318 19796 33324 19808
rect 33376 19796 33382 19848
rect 35989 19839 36047 19845
rect 35989 19805 36001 19839
rect 36035 19805 36047 19839
rect 35989 19799 36047 19805
rect 27249 19771 27307 19777
rect 27249 19768 27261 19771
rect 26936 19740 27261 19768
rect 26936 19728 26942 19740
rect 27249 19737 27261 19740
rect 27295 19737 27307 19771
rect 28626 19768 28632 19780
rect 27249 19731 27307 19737
rect 27356 19740 28632 19768
rect 2222 19660 2228 19712
rect 2280 19700 2286 19712
rect 2317 19703 2375 19709
rect 2317 19700 2329 19703
rect 2280 19672 2329 19700
rect 2280 19660 2286 19672
rect 2317 19669 2329 19672
rect 2363 19669 2375 19703
rect 5166 19700 5172 19712
rect 5127 19672 5172 19700
rect 2317 19663 2375 19669
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 6822 19660 6828 19712
rect 6880 19700 6886 19712
rect 7561 19703 7619 19709
rect 7561 19700 7573 19703
rect 6880 19672 7573 19700
rect 6880 19660 6886 19672
rect 7561 19669 7573 19672
rect 7607 19669 7619 19703
rect 8938 19700 8944 19712
rect 8899 19672 8944 19700
rect 7561 19663 7619 19669
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 11977 19703 12035 19709
rect 11977 19669 11989 19703
rect 12023 19700 12035 19703
rect 12526 19700 12532 19712
rect 12023 19672 12532 19700
rect 12023 19669 12035 19672
rect 11977 19663 12035 19669
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 12768 19672 14289 19700
rect 12768 19660 12774 19672
rect 14277 19669 14289 19672
rect 14323 19669 14335 19703
rect 14918 19700 14924 19712
rect 14879 19672 14924 19700
rect 14277 19663 14335 19669
rect 14918 19660 14924 19672
rect 14976 19660 14982 19712
rect 15841 19703 15899 19709
rect 15841 19669 15853 19703
rect 15887 19700 15899 19703
rect 15930 19700 15936 19712
rect 15887 19672 15936 19700
rect 15887 19669 15899 19672
rect 15841 19663 15899 19669
rect 15930 19660 15936 19672
rect 15988 19700 15994 19712
rect 22002 19700 22008 19712
rect 15988 19672 22008 19700
rect 15988 19660 15994 19672
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 25314 19660 25320 19712
rect 25372 19700 25378 19712
rect 27356 19700 27384 19740
rect 28626 19728 28632 19740
rect 28684 19728 28690 19780
rect 28721 19771 28779 19777
rect 28721 19737 28733 19771
rect 28767 19768 28779 19771
rect 32674 19768 32680 19780
rect 28767 19740 32680 19768
rect 28767 19737 28779 19740
rect 28721 19731 28779 19737
rect 32674 19728 32680 19740
rect 32732 19728 32738 19780
rect 36004 19768 36032 19799
rect 37458 19796 37464 19848
rect 37516 19836 37522 19848
rect 37553 19839 37611 19845
rect 37553 19836 37565 19839
rect 37516 19808 37565 19836
rect 37516 19796 37522 19808
rect 37553 19805 37565 19808
rect 37599 19805 37611 19839
rect 40420 19836 40448 20012
rect 41417 20009 41429 20012
rect 41463 20009 41475 20043
rect 41417 20003 41475 20009
rect 40494 19864 40500 19916
rect 40552 19904 40558 19916
rect 40552 19876 40724 19904
rect 40552 19864 40558 19876
rect 40696 19845 40724 19876
rect 40589 19839 40647 19845
rect 40589 19836 40601 19839
rect 40420 19808 40601 19836
rect 37553 19799 37611 19805
rect 40589 19805 40601 19808
rect 40635 19805 40647 19839
rect 40589 19799 40647 19805
rect 40681 19839 40739 19845
rect 40681 19805 40693 19839
rect 40727 19805 40739 19839
rect 40681 19799 40739 19805
rect 40770 19796 40776 19848
rect 40828 19836 40834 19848
rect 40954 19836 40960 19848
rect 40828 19808 40873 19836
rect 40915 19808 40960 19836
rect 40828 19796 40834 19808
rect 40954 19796 40960 19808
rect 41012 19796 41018 19848
rect 58158 19836 58164 19848
rect 58119 19808 58164 19836
rect 58158 19796 58164 19808
rect 58216 19796 58222 19848
rect 37642 19768 37648 19780
rect 36004 19740 37648 19768
rect 37642 19728 37648 19740
rect 37700 19728 37706 19780
rect 40402 19768 40408 19780
rect 38672 19740 40408 19768
rect 25372 19672 27384 19700
rect 32493 19703 32551 19709
rect 25372 19660 25378 19672
rect 32493 19669 32505 19703
rect 32539 19700 32551 19703
rect 32950 19700 32956 19712
rect 32539 19672 32956 19700
rect 32539 19669 32551 19672
rect 32493 19663 32551 19669
rect 32950 19660 32956 19672
rect 33008 19660 33014 19712
rect 36078 19660 36084 19712
rect 36136 19700 36142 19712
rect 38672 19700 38700 19740
rect 40402 19728 40408 19740
rect 40460 19728 40466 19780
rect 36136 19672 38700 19700
rect 36136 19660 36142 19672
rect 38746 19660 38752 19712
rect 38804 19700 38810 19712
rect 38841 19703 38899 19709
rect 38841 19700 38853 19703
rect 38804 19672 38853 19700
rect 38804 19660 38810 19672
rect 38841 19669 38853 19672
rect 38887 19669 38899 19703
rect 40310 19700 40316 19712
rect 40271 19672 40316 19700
rect 38841 19663 38899 19669
rect 40310 19660 40316 19672
rect 40368 19660 40374 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 3329 19499 3387 19505
rect 3329 19465 3341 19499
rect 3375 19496 3387 19499
rect 4614 19496 4620 19508
rect 3375 19468 4620 19496
rect 3375 19465 3387 19468
rect 3329 19459 3387 19465
rect 4614 19456 4620 19468
rect 4672 19456 4678 19508
rect 10597 19499 10655 19505
rect 10597 19465 10609 19499
rect 10643 19496 10655 19499
rect 10778 19496 10784 19508
rect 10643 19468 10784 19496
rect 10643 19465 10655 19468
rect 10597 19459 10655 19465
rect 10778 19456 10784 19468
rect 10836 19456 10842 19508
rect 14090 19456 14096 19508
rect 14148 19496 14154 19508
rect 14185 19499 14243 19505
rect 14185 19496 14197 19499
rect 14148 19468 14197 19496
rect 14148 19456 14154 19468
rect 14185 19465 14197 19468
rect 14231 19465 14243 19499
rect 14185 19459 14243 19465
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 15289 19499 15347 19505
rect 15289 19496 15301 19499
rect 15252 19468 15301 19496
rect 15252 19456 15258 19468
rect 15289 19465 15301 19468
rect 15335 19465 15347 19499
rect 15289 19459 15347 19465
rect 18785 19499 18843 19505
rect 18785 19465 18797 19499
rect 18831 19496 18843 19499
rect 18966 19496 18972 19508
rect 18831 19468 18972 19496
rect 18831 19465 18843 19468
rect 18785 19459 18843 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 22373 19499 22431 19505
rect 22373 19465 22385 19499
rect 22419 19496 22431 19499
rect 23474 19496 23480 19508
rect 22419 19468 23480 19496
rect 22419 19465 22431 19468
rect 22373 19459 22431 19465
rect 23474 19456 23480 19468
rect 23532 19496 23538 19508
rect 23934 19496 23940 19508
rect 23532 19468 23940 19496
rect 23532 19456 23538 19468
rect 23934 19456 23940 19468
rect 23992 19456 23998 19508
rect 26418 19496 26424 19508
rect 26379 19468 26424 19496
rect 26418 19456 26424 19468
rect 26476 19456 26482 19508
rect 26970 19496 26976 19508
rect 26931 19468 26976 19496
rect 26970 19456 26976 19468
rect 27028 19456 27034 19508
rect 28626 19456 28632 19508
rect 28684 19496 28690 19508
rect 29181 19499 29239 19505
rect 28684 19468 29132 19496
rect 28684 19456 28690 19468
rect 2682 19428 2688 19440
rect 1964 19400 2688 19428
rect 1964 19372 1992 19400
rect 2682 19388 2688 19400
rect 2740 19428 2746 19440
rect 3789 19431 3847 19437
rect 2740 19388 2774 19428
rect 3789 19397 3801 19431
rect 3835 19428 3847 19431
rect 5166 19428 5172 19440
rect 3835 19400 5172 19428
rect 3835 19397 3847 19400
rect 3789 19391 3847 19397
rect 5166 19388 5172 19400
rect 5224 19428 5230 19440
rect 6546 19428 6552 19440
rect 5224 19400 6552 19428
rect 5224 19388 5230 19400
rect 6546 19388 6552 19400
rect 6604 19388 6610 19440
rect 9582 19428 9588 19440
rect 9232 19400 9588 19428
rect 1946 19360 1952 19372
rect 1907 19332 1952 19360
rect 1946 19320 1952 19332
rect 2004 19320 2010 19372
rect 2222 19369 2228 19372
rect 2216 19360 2228 19369
rect 2183 19332 2228 19360
rect 2216 19323 2228 19332
rect 2222 19320 2228 19323
rect 2280 19320 2286 19372
rect 2746 19360 2774 19388
rect 6914 19369 6920 19372
rect 6641 19363 6699 19369
rect 2746 19332 3556 19360
rect 3528 19292 3556 19332
rect 6641 19329 6653 19363
rect 6687 19329 6699 19363
rect 6641 19323 6699 19329
rect 6908 19323 6920 19369
rect 6972 19360 6978 19372
rect 9232 19369 9260 19400
rect 9582 19388 9588 19400
rect 9640 19428 9646 19440
rect 12434 19428 12440 19440
rect 9640 19400 12440 19428
rect 9640 19388 9646 19400
rect 12434 19388 12440 19400
rect 12492 19428 12498 19440
rect 13170 19428 13176 19440
rect 12492 19400 13176 19428
rect 12492 19388 12498 19400
rect 13170 19388 13176 19400
rect 13228 19388 13234 19440
rect 20990 19428 20996 19440
rect 15672 19400 20996 19428
rect 9217 19363 9275 19369
rect 6972 19332 7008 19360
rect 6362 19292 6368 19304
rect 3528 19264 6368 19292
rect 5092 19233 5120 19264
rect 6362 19252 6368 19264
rect 6420 19292 6426 19304
rect 6656 19292 6684 19323
rect 6914 19320 6920 19323
rect 6972 19320 6978 19332
rect 9217 19329 9229 19363
rect 9263 19329 9275 19363
rect 9217 19323 9275 19329
rect 9484 19363 9542 19369
rect 9484 19329 9496 19363
rect 9530 19360 9542 19363
rect 10410 19360 10416 19372
rect 9530 19332 10416 19360
rect 9530 19329 9542 19332
rect 9484 19323 9542 19329
rect 10410 19320 10416 19332
rect 10468 19320 10474 19372
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 10836 19332 11713 19360
rect 10836 19320 10842 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 12710 19360 12716 19372
rect 11931 19332 12716 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 14182 19360 14188 19372
rect 14143 19332 14188 19360
rect 14182 19320 14188 19332
rect 14240 19320 14246 19372
rect 14274 19320 14280 19372
rect 14332 19360 14338 19372
rect 15672 19369 15700 19400
rect 20990 19388 20996 19400
rect 21048 19388 21054 19440
rect 22094 19428 22100 19440
rect 21284 19400 22100 19428
rect 14369 19363 14427 19369
rect 14369 19360 14381 19363
rect 14332 19332 14381 19360
rect 14332 19320 14338 19332
rect 14369 19329 14381 19332
rect 14415 19329 14427 19363
rect 14369 19323 14427 19329
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19329 15715 19363
rect 17402 19360 17408 19372
rect 17363 19332 17408 19360
rect 15657 19323 15715 19329
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 17494 19320 17500 19372
rect 17552 19360 17558 19372
rect 17661 19363 17719 19369
rect 17661 19360 17673 19363
rect 17552 19332 17673 19360
rect 17552 19320 17558 19332
rect 17661 19329 17673 19332
rect 17707 19329 17719 19363
rect 17661 19323 17719 19329
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 21284 19369 21312 19400
rect 22094 19388 22100 19400
rect 22152 19388 22158 19440
rect 24762 19388 24768 19440
rect 24820 19428 24826 19440
rect 25314 19428 25320 19440
rect 24820 19400 25320 19428
rect 24820 19388 24826 19400
rect 25314 19388 25320 19400
rect 25372 19428 25378 19440
rect 25409 19431 25467 19437
rect 25409 19428 25421 19431
rect 25372 19400 25421 19428
rect 25372 19388 25378 19400
rect 25409 19397 25421 19400
rect 25455 19397 25467 19431
rect 25409 19391 25467 19397
rect 25498 19388 25504 19440
rect 25556 19428 25562 19440
rect 25556 19400 25601 19428
rect 25556 19388 25562 19400
rect 27246 19388 27252 19440
rect 27304 19428 27310 19440
rect 27433 19431 27491 19437
rect 27433 19428 27445 19431
rect 27304 19400 27445 19428
rect 27304 19388 27310 19400
rect 27433 19397 27445 19400
rect 27479 19397 27491 19431
rect 27433 19391 27491 19397
rect 28258 19388 28264 19440
rect 28316 19428 28322 19440
rect 28905 19431 28963 19437
rect 28905 19428 28917 19431
rect 28316 19400 28917 19428
rect 28316 19388 28322 19400
rect 28905 19397 28917 19400
rect 28951 19397 28963 19431
rect 29104 19428 29132 19468
rect 29181 19465 29193 19499
rect 29227 19496 29239 19499
rect 30926 19496 30932 19508
rect 29227 19468 30420 19496
rect 30887 19468 30932 19496
rect 29227 19465 29239 19468
rect 29181 19459 29239 19465
rect 29454 19428 29460 19440
rect 29104 19400 29460 19428
rect 28905 19391 28963 19397
rect 29454 19388 29460 19400
rect 29512 19428 29518 19440
rect 29512 19400 29684 19428
rect 29512 19388 29518 19400
rect 21269 19363 21327 19369
rect 20588 19332 21036 19360
rect 20588 19320 20594 19332
rect 12526 19292 12532 19304
rect 6420 19264 6684 19292
rect 10244 19264 12532 19292
rect 6420 19252 6426 19264
rect 5077 19227 5135 19233
rect 5077 19193 5089 19227
rect 5123 19193 5135 19227
rect 5077 19187 5135 19193
rect 7742 19184 7748 19236
rect 7800 19224 7806 19236
rect 8110 19224 8116 19236
rect 7800 19196 8116 19224
rect 7800 19184 7806 19196
rect 8110 19184 8116 19196
rect 8168 19224 8174 19236
rect 8168 19196 8616 19224
rect 8168 19184 8174 19196
rect 7650 19116 7656 19168
rect 7708 19156 7714 19168
rect 8021 19159 8079 19165
rect 8021 19156 8033 19159
rect 7708 19128 8033 19156
rect 7708 19116 7714 19128
rect 8021 19125 8033 19128
rect 8067 19125 8079 19159
rect 8021 19119 8079 19125
rect 8202 19116 8208 19168
rect 8260 19156 8266 19168
rect 8478 19156 8484 19168
rect 8260 19128 8484 19156
rect 8260 19116 8266 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8588 19156 8616 19196
rect 10244 19156 10272 19264
rect 12526 19252 12532 19264
rect 12584 19292 12590 19304
rect 13722 19292 13728 19304
rect 12584 19264 13728 19292
rect 12584 19252 12590 19264
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 21008 19301 21036 19332
rect 21269 19329 21281 19363
rect 21315 19329 21327 19363
rect 22186 19360 22192 19372
rect 22147 19332 22192 19360
rect 21269 19323 21327 19329
rect 22186 19320 22192 19332
rect 22244 19360 22250 19372
rect 22738 19360 22744 19372
rect 22244 19332 22744 19360
rect 22244 19320 22250 19332
rect 22738 19320 22744 19332
rect 22796 19320 22802 19372
rect 24394 19320 24400 19372
rect 24452 19360 24458 19372
rect 25225 19363 25283 19369
rect 25225 19360 25237 19363
rect 24452 19332 25237 19360
rect 24452 19320 24458 19332
rect 25225 19329 25237 19332
rect 25271 19329 25283 19363
rect 25590 19360 25596 19372
rect 25225 19323 25283 19329
rect 25424 19332 25596 19360
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19261 15623 19295
rect 15565 19255 15623 19261
rect 20993 19295 21051 19301
rect 20993 19261 21005 19295
rect 21039 19261 21051 19295
rect 22002 19292 22008 19304
rect 21963 19264 22008 19292
rect 20993 19255 21051 19261
rect 11146 19184 11152 19236
rect 11204 19224 11210 19236
rect 12158 19224 12164 19236
rect 11204 19196 12164 19224
rect 11204 19184 11210 19196
rect 12158 19184 12164 19196
rect 12216 19224 12222 19236
rect 12345 19227 12403 19233
rect 12345 19224 12357 19227
rect 12216 19196 12357 19224
rect 12216 19184 12222 19196
rect 12345 19193 12357 19196
rect 12391 19193 12403 19227
rect 12345 19187 12403 19193
rect 8588 19128 10272 19156
rect 10870 19116 10876 19168
rect 10928 19156 10934 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 10928 19128 11529 19156
rect 10928 19116 10934 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 15470 19156 15476 19168
rect 15431 19128 15476 19156
rect 11517 19119 11575 19125
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15580 19156 15608 19255
rect 22002 19252 22008 19264
rect 22060 19292 22066 19304
rect 22833 19295 22891 19301
rect 22833 19292 22845 19295
rect 22060 19264 22845 19292
rect 22060 19252 22066 19264
rect 22833 19261 22845 19264
rect 22879 19261 22891 19295
rect 22833 19255 22891 19261
rect 24946 19252 24952 19304
rect 25004 19292 25010 19304
rect 25424 19292 25452 19332
rect 25590 19320 25596 19332
rect 25648 19320 25654 19372
rect 27154 19360 27160 19372
rect 27115 19332 27160 19360
rect 27154 19320 27160 19332
rect 27212 19320 27218 19372
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 28629 19363 28687 19369
rect 28629 19360 28641 19363
rect 27396 19332 28641 19360
rect 27396 19320 27402 19332
rect 28629 19329 28641 19332
rect 28675 19329 28687 19363
rect 28629 19323 28687 19329
rect 28813 19363 28871 19369
rect 28813 19329 28825 19363
rect 28859 19360 28871 19363
rect 28997 19363 29055 19369
rect 28859 19332 28948 19360
rect 28859 19329 28871 19332
rect 28813 19323 28871 19329
rect 27246 19292 27252 19304
rect 25004 19264 25452 19292
rect 27207 19264 27252 19292
rect 25004 19252 25010 19264
rect 27246 19252 27252 19264
rect 27304 19252 27310 19304
rect 28920 19292 28948 19332
rect 28997 19329 29009 19363
rect 29043 19360 29055 19363
rect 29043 19332 29132 19360
rect 29043 19329 29055 19332
rect 28997 19323 29055 19329
rect 28920 19264 29040 19292
rect 18708 19196 18920 19224
rect 18708 19156 18736 19196
rect 15580 19128 18736 19156
rect 18892 19156 18920 19196
rect 18966 19184 18972 19236
rect 19024 19224 19030 19236
rect 25682 19224 25688 19236
rect 19024 19196 25688 19224
rect 19024 19184 19030 19196
rect 25682 19184 25688 19196
rect 25740 19184 25746 19236
rect 25777 19227 25835 19233
rect 25777 19193 25789 19227
rect 25823 19224 25835 19227
rect 25823 19196 27200 19224
rect 25823 19193 25835 19196
rect 25777 19187 25835 19193
rect 22186 19156 22192 19168
rect 18892 19128 22192 19156
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 22462 19116 22468 19168
rect 22520 19156 22526 19168
rect 26418 19156 26424 19168
rect 22520 19128 26424 19156
rect 22520 19116 22526 19128
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 27172 19165 27200 19196
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19125 27215 19159
rect 27890 19156 27896 19168
rect 27851 19128 27896 19156
rect 27157 19119 27215 19125
rect 27890 19116 27896 19128
rect 27948 19116 27954 19168
rect 29012 19156 29040 19264
rect 29104 19224 29132 19332
rect 29656 19301 29684 19400
rect 29641 19295 29699 19301
rect 29641 19261 29653 19295
rect 29687 19261 29699 19295
rect 29914 19292 29920 19304
rect 29875 19264 29920 19292
rect 29641 19255 29699 19261
rect 29914 19252 29920 19264
rect 29972 19252 29978 19304
rect 30006 19224 30012 19236
rect 29104 19196 30012 19224
rect 30006 19184 30012 19196
rect 30064 19184 30070 19236
rect 29822 19156 29828 19168
rect 29012 19128 29828 19156
rect 29822 19116 29828 19128
rect 29880 19116 29886 19168
rect 30392 19156 30420 19468
rect 30926 19456 30932 19468
rect 30984 19456 30990 19508
rect 35805 19499 35863 19505
rect 35805 19496 35817 19499
rect 31128 19468 35817 19496
rect 31128 19369 31156 19468
rect 35805 19465 35817 19468
rect 35851 19465 35863 19499
rect 35805 19459 35863 19465
rect 37550 19456 37556 19508
rect 37608 19496 37614 19508
rect 40129 19499 40187 19505
rect 40129 19496 40141 19499
rect 37608 19468 40141 19496
rect 37608 19456 37614 19468
rect 40129 19465 40141 19468
rect 40175 19496 40187 19499
rect 40175 19468 40448 19496
rect 40175 19465 40187 19468
rect 40129 19459 40187 19465
rect 31389 19431 31447 19437
rect 31389 19397 31401 19431
rect 31435 19428 31447 19431
rect 31662 19428 31668 19440
rect 31435 19400 31668 19428
rect 31435 19397 31447 19400
rect 31389 19391 31447 19397
rect 31662 19388 31668 19400
rect 31720 19388 31726 19440
rect 36078 19428 36084 19440
rect 36039 19400 36084 19428
rect 36078 19388 36084 19400
rect 36136 19388 36142 19440
rect 36173 19431 36231 19437
rect 36173 19397 36185 19431
rect 36219 19428 36231 19431
rect 36262 19428 36268 19440
rect 36219 19400 36268 19428
rect 36219 19397 36231 19400
rect 36173 19391 36231 19397
rect 36262 19388 36268 19400
rect 36320 19388 36326 19440
rect 38010 19428 38016 19440
rect 36372 19400 38016 19428
rect 31113 19363 31171 19369
rect 31113 19329 31125 19363
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 31202 19320 31208 19372
rect 31260 19360 31266 19372
rect 31260 19332 31305 19360
rect 31260 19320 31266 19332
rect 33226 19320 33232 19372
rect 33284 19360 33290 19372
rect 33790 19363 33848 19369
rect 33790 19360 33802 19363
rect 33284 19332 33802 19360
rect 33284 19320 33290 19332
rect 33790 19329 33802 19332
rect 33836 19329 33848 19363
rect 33790 19323 33848 19329
rect 34057 19363 34115 19369
rect 34057 19329 34069 19363
rect 34103 19360 34115 19363
rect 34146 19360 34152 19372
rect 34103 19332 34152 19360
rect 34103 19329 34115 19332
rect 34057 19323 34115 19329
rect 34146 19320 34152 19332
rect 34204 19320 34210 19372
rect 35802 19320 35808 19372
rect 35860 19360 35866 19372
rect 35986 19360 35992 19372
rect 35860 19332 35992 19360
rect 35860 19320 35866 19332
rect 35986 19320 35992 19332
rect 36044 19320 36050 19372
rect 36372 19369 36400 19400
rect 38010 19388 38016 19400
rect 38068 19388 38074 19440
rect 39016 19431 39074 19437
rect 39016 19397 39028 19431
rect 39062 19428 39074 19431
rect 40310 19428 40316 19440
rect 39062 19400 40316 19428
rect 39062 19397 39074 19400
rect 39016 19391 39074 19397
rect 40310 19388 40316 19400
rect 40368 19388 40374 19440
rect 40420 19428 40448 19468
rect 40770 19456 40776 19508
rect 40828 19496 40834 19508
rect 40957 19499 41015 19505
rect 40957 19496 40969 19499
rect 40828 19468 40969 19496
rect 40828 19456 40834 19468
rect 40957 19465 40969 19468
rect 41003 19465 41015 19499
rect 40957 19459 41015 19465
rect 40420 19400 40816 19428
rect 36357 19363 36415 19369
rect 36357 19329 36369 19363
rect 36403 19329 36415 19363
rect 37553 19363 37611 19369
rect 37553 19360 37565 19363
rect 36357 19323 36415 19329
rect 36464 19332 37565 19360
rect 36004 19292 36032 19320
rect 36464 19292 36492 19332
rect 37553 19329 37565 19332
rect 37599 19329 37611 19363
rect 40586 19360 40592 19372
rect 40547 19332 40592 19360
rect 37553 19323 37611 19329
rect 40586 19320 40592 19332
rect 40644 19320 40650 19372
rect 40788 19369 40816 19400
rect 40773 19363 40831 19369
rect 40773 19329 40785 19363
rect 40819 19329 40831 19363
rect 40773 19323 40831 19329
rect 37274 19292 37280 19304
rect 36004 19264 36492 19292
rect 37235 19264 37280 19292
rect 37274 19252 37280 19264
rect 37332 19252 37338 19304
rect 38746 19292 38752 19304
rect 38707 19264 38752 19292
rect 38746 19252 38752 19264
rect 38804 19252 38810 19304
rect 32674 19224 32680 19236
rect 32635 19196 32680 19224
rect 32674 19184 32680 19196
rect 32732 19184 32738 19236
rect 31113 19159 31171 19165
rect 31113 19156 31125 19159
rect 30392 19128 31125 19156
rect 31113 19125 31125 19128
rect 31159 19125 31171 19159
rect 31113 19119 31171 19125
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 2498 18952 2504 18964
rect 2459 18924 2504 18952
rect 2498 18912 2504 18924
rect 2556 18912 2562 18964
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 5445 18955 5503 18961
rect 5445 18952 5457 18955
rect 4028 18924 5457 18952
rect 4028 18912 4034 18924
rect 5445 18921 5457 18924
rect 5491 18921 5503 18955
rect 5445 18915 5503 18921
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 7742 18952 7748 18964
rect 7239 18924 7748 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 4065 18887 4123 18893
rect 4065 18884 4077 18887
rect 2746 18856 4077 18884
rect 2746 18816 2774 18856
rect 4065 18853 4077 18856
rect 4111 18853 4123 18887
rect 5460 18884 5488 18915
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 8294 18952 8300 18964
rect 8255 18924 8300 18952
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 8386 18912 8392 18964
rect 8444 18952 8450 18964
rect 10410 18952 10416 18964
rect 8444 18924 10272 18952
rect 10371 18924 10416 18952
rect 8444 18912 8450 18924
rect 8110 18884 8116 18896
rect 5460 18856 8116 18884
rect 4065 18847 4123 18853
rect 8110 18844 8116 18856
rect 8168 18844 8174 18896
rect 10244 18884 10272 18924
rect 10410 18912 10416 18924
rect 10468 18912 10474 18964
rect 13906 18952 13912 18964
rect 10520 18924 13912 18952
rect 10520 18884 10548 18924
rect 13906 18912 13912 18924
rect 13964 18912 13970 18964
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 14240 18924 14473 18952
rect 14240 18912 14246 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 17494 18952 17500 18964
rect 17455 18924 17500 18952
rect 14461 18915 14519 18921
rect 17494 18912 17500 18924
rect 17552 18912 17558 18964
rect 22002 18912 22008 18964
rect 22060 18952 22066 18964
rect 22189 18955 22247 18961
rect 22189 18952 22201 18955
rect 22060 18924 22201 18952
rect 22060 18912 22066 18924
rect 22189 18921 22201 18924
rect 22235 18952 22247 18955
rect 27338 18952 27344 18964
rect 22235 18924 27344 18952
rect 22235 18921 22247 18924
rect 22189 18915 22247 18921
rect 27338 18912 27344 18924
rect 27396 18912 27402 18964
rect 30193 18955 30251 18961
rect 30193 18921 30205 18955
rect 30239 18952 30251 18955
rect 30837 18955 30895 18961
rect 30837 18952 30849 18955
rect 30239 18924 30849 18952
rect 30239 18921 30251 18924
rect 30193 18915 30251 18921
rect 30837 18921 30849 18924
rect 30883 18921 30895 18955
rect 35897 18955 35955 18961
rect 35897 18952 35909 18955
rect 30837 18915 30895 18921
rect 30944 18924 35909 18952
rect 10244 18856 10548 18884
rect 10704 18856 12434 18884
rect 2700 18788 2774 18816
rect 4709 18819 4767 18825
rect 2700 18757 2728 18788
rect 4709 18785 4721 18819
rect 4755 18816 4767 18819
rect 4798 18816 4804 18828
rect 4755 18788 4804 18816
rect 4755 18785 4767 18788
rect 4709 18779 4767 18785
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 6822 18816 6828 18828
rect 5184 18788 6828 18816
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 2774 18708 2780 18760
rect 2832 18748 2838 18760
rect 4433 18751 4491 18757
rect 2832 18720 2877 18748
rect 2832 18708 2838 18720
rect 4433 18717 4445 18751
rect 4479 18748 4491 18751
rect 5184 18748 5212 18788
rect 6822 18776 6828 18788
rect 6880 18776 6886 18828
rect 8294 18816 8300 18828
rect 8255 18788 8300 18816
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 7006 18748 7012 18760
rect 4479 18720 5212 18748
rect 6967 18720 7012 18748
rect 4479 18717 4491 18720
rect 4433 18711 4491 18717
rect 7006 18708 7012 18720
rect 7064 18748 7070 18760
rect 8202 18748 8208 18760
rect 7064 18720 8208 18748
rect 7064 18708 7070 18720
rect 8202 18708 8208 18720
rect 8260 18708 8266 18760
rect 8386 18748 8392 18760
rect 8347 18720 8392 18748
rect 8386 18708 8392 18720
rect 8444 18708 8450 18760
rect 10704 18757 10732 18856
rect 12406 18816 12434 18856
rect 13446 18844 13452 18896
rect 13504 18884 13510 18896
rect 17954 18884 17960 18896
rect 13504 18856 17960 18884
rect 13504 18844 13510 18856
rect 17954 18844 17960 18856
rect 18012 18844 18018 18896
rect 23201 18887 23259 18893
rect 23201 18853 23213 18887
rect 23247 18884 23259 18887
rect 24578 18884 24584 18896
rect 23247 18856 24584 18884
rect 23247 18853 23259 18856
rect 23201 18847 23259 18853
rect 24578 18844 24584 18856
rect 24636 18844 24642 18896
rect 26878 18884 26884 18896
rect 24688 18856 26884 18884
rect 15010 18816 15016 18828
rect 10796 18788 11928 18816
rect 12406 18788 15016 18816
rect 10796 18757 10824 18788
rect 10689 18751 10747 18757
rect 10689 18748 10701 18751
rect 9646 18720 10701 18748
rect 4525 18683 4583 18689
rect 4525 18649 4537 18683
rect 4571 18680 4583 18683
rect 4614 18680 4620 18692
rect 4571 18652 4620 18680
rect 4571 18649 4583 18652
rect 4525 18643 4583 18649
rect 4614 18640 4620 18652
rect 4672 18640 4678 18692
rect 5350 18680 5356 18692
rect 5311 18652 5356 18680
rect 5350 18640 5356 18652
rect 5408 18640 5414 18692
rect 5902 18640 5908 18692
rect 5960 18680 5966 18692
rect 6457 18683 6515 18689
rect 6457 18680 6469 18683
rect 5960 18652 6469 18680
rect 5960 18640 5966 18652
rect 6457 18649 6469 18652
rect 6503 18649 6515 18683
rect 8570 18680 8576 18692
rect 6457 18643 6515 18649
rect 7116 18652 8576 18680
rect 6365 18615 6423 18621
rect 6365 18581 6377 18615
rect 6411 18612 6423 18615
rect 7116 18612 7144 18652
rect 8570 18640 8576 18652
rect 8628 18640 8634 18692
rect 6411 18584 7144 18612
rect 6411 18581 6423 18584
rect 6365 18575 6423 18581
rect 7374 18572 7380 18624
rect 7432 18612 7438 18624
rect 8021 18615 8079 18621
rect 8021 18612 8033 18615
rect 7432 18584 8033 18612
rect 7432 18572 7438 18584
rect 8021 18581 8033 18584
rect 8067 18581 8079 18615
rect 8021 18575 8079 18581
rect 8110 18572 8116 18624
rect 8168 18612 8174 18624
rect 9309 18615 9367 18621
rect 9309 18612 9321 18615
rect 8168 18584 9321 18612
rect 8168 18572 8174 18584
rect 9309 18581 9321 18584
rect 9355 18612 9367 18615
rect 9646 18612 9674 18720
rect 10689 18717 10701 18720
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 10781 18751 10839 18757
rect 10781 18717 10793 18751
rect 10827 18717 10839 18751
rect 10781 18711 10839 18717
rect 10870 18708 10876 18760
rect 10928 18748 10934 18760
rect 11057 18751 11115 18757
rect 10928 18720 10973 18748
rect 10928 18708 10934 18720
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11146 18748 11152 18760
rect 11103 18720 11152 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11146 18708 11152 18720
rect 11204 18708 11210 18760
rect 11790 18748 11796 18760
rect 11751 18720 11796 18748
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 11900 18757 11928 18788
rect 15010 18776 15016 18788
rect 15068 18776 15074 18828
rect 15120 18788 20668 18816
rect 11885 18751 11943 18757
rect 11885 18717 11897 18751
rect 11931 18717 11943 18751
rect 11885 18711 11943 18717
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18717 12035 18751
rect 12158 18748 12164 18760
rect 12119 18720 12164 18748
rect 11977 18711 12035 18717
rect 9861 18683 9919 18689
rect 9861 18649 9873 18683
rect 9907 18680 9919 18683
rect 11808 18680 11836 18708
rect 9907 18652 11836 18680
rect 9907 18649 9919 18652
rect 9861 18643 9919 18649
rect 11514 18612 11520 18624
rect 9355 18584 9674 18612
rect 11475 18584 11520 18612
rect 9355 18581 9367 18584
rect 9309 18575 9367 18581
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 11900 18612 11928 18711
rect 11992 18680 12020 18711
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 12250 18708 12256 18760
rect 12308 18748 12314 18760
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12308 18720 12817 18748
rect 12308 18708 12314 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 12894 18708 12900 18760
rect 12952 18748 12958 18760
rect 15120 18748 15148 18788
rect 12952 18720 15148 18748
rect 12952 18708 12958 18720
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 17037 18751 17095 18757
rect 17037 18748 17049 18751
rect 16632 18720 17049 18748
rect 16632 18708 16638 18720
rect 17037 18717 17049 18720
rect 17083 18748 17095 18751
rect 17773 18751 17831 18757
rect 17773 18748 17785 18751
rect 17083 18720 17785 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17773 18717 17785 18720
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18748 18015 18751
rect 18046 18748 18052 18760
rect 18003 18720 18052 18748
rect 18003 18717 18015 18720
rect 17957 18711 18015 18717
rect 12621 18683 12679 18689
rect 12621 18680 12633 18683
rect 11992 18652 12633 18680
rect 12621 18649 12633 18652
rect 12667 18649 12679 18683
rect 12621 18643 12679 18649
rect 12710 18640 12716 18692
rect 12768 18680 12774 18692
rect 12989 18683 13047 18689
rect 12989 18680 13001 18683
rect 12768 18652 13001 18680
rect 12768 18640 12774 18652
rect 12989 18649 13001 18652
rect 13035 18649 13047 18683
rect 12989 18643 13047 18649
rect 17880 18680 17908 18711
rect 18046 18708 18052 18720
rect 18104 18708 18110 18760
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18748 18199 18751
rect 18322 18748 18328 18760
rect 18187 18720 18328 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 18322 18708 18328 18720
rect 18380 18708 18386 18760
rect 20530 18680 20536 18692
rect 17880 18652 20536 18680
rect 12802 18612 12808 18624
rect 11900 18584 12808 18612
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 17880 18612 17908 18652
rect 20530 18640 20536 18652
rect 20588 18640 20594 18692
rect 17828 18584 17908 18612
rect 20640 18612 20668 18788
rect 22370 18776 22376 18828
rect 22428 18816 22434 18828
rect 24688 18825 24716 18856
rect 26878 18844 26884 18856
rect 26936 18844 26942 18896
rect 27154 18844 27160 18896
rect 27212 18884 27218 18896
rect 30374 18884 30380 18896
rect 27212 18856 30380 18884
rect 27212 18844 27218 18856
rect 30374 18844 30380 18856
rect 30432 18844 30438 18896
rect 30650 18884 30656 18896
rect 30611 18856 30656 18884
rect 30650 18844 30656 18856
rect 30708 18844 30714 18896
rect 30944 18884 30972 18924
rect 35897 18921 35909 18924
rect 35943 18921 35955 18955
rect 35897 18915 35955 18921
rect 37277 18955 37335 18961
rect 37277 18921 37289 18955
rect 37323 18952 37335 18955
rect 37366 18952 37372 18964
rect 37323 18924 37372 18952
rect 37323 18921 37335 18924
rect 37277 18915 37335 18921
rect 37366 18912 37372 18924
rect 37424 18912 37430 18964
rect 30852 18856 30972 18884
rect 24397 18819 24455 18825
rect 24397 18816 24409 18819
rect 22428 18788 24409 18816
rect 22428 18776 22434 18788
rect 24397 18785 24409 18788
rect 24443 18785 24455 18819
rect 24397 18779 24455 18785
rect 24673 18819 24731 18825
rect 24673 18785 24685 18819
rect 24719 18785 24731 18819
rect 24673 18779 24731 18785
rect 25682 18776 25688 18828
rect 25740 18816 25746 18828
rect 25740 18788 29684 18816
rect 25740 18776 25746 18788
rect 20806 18748 20812 18760
rect 20767 18720 20812 18748
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 25498 18708 25504 18760
rect 25556 18748 25562 18760
rect 25961 18751 26019 18757
rect 25961 18748 25973 18751
rect 25556 18720 25973 18748
rect 25556 18708 25562 18720
rect 25961 18717 25973 18720
rect 26007 18717 26019 18751
rect 25961 18711 26019 18717
rect 26602 18708 26608 18760
rect 26660 18708 26666 18760
rect 29656 18757 29684 18788
rect 29641 18751 29699 18757
rect 29641 18717 29653 18751
rect 29687 18717 29699 18751
rect 29822 18748 29828 18760
rect 29783 18720 29828 18748
rect 29641 18711 29699 18717
rect 29822 18708 29828 18720
rect 29880 18708 29886 18760
rect 30006 18748 30012 18760
rect 29967 18720 30012 18748
rect 30006 18708 30012 18720
rect 30064 18708 30070 18760
rect 30852 18757 30880 18856
rect 32030 18844 32036 18896
rect 32088 18884 32094 18896
rect 32769 18887 32827 18893
rect 32769 18884 32781 18887
rect 32088 18856 32781 18884
rect 32088 18844 32094 18856
rect 32769 18853 32781 18856
rect 32815 18884 32827 18887
rect 32858 18884 32864 18896
rect 32815 18856 32864 18884
rect 32815 18853 32827 18856
rect 32769 18847 32827 18853
rect 32858 18844 32864 18856
rect 32916 18844 32922 18896
rect 34146 18816 34152 18828
rect 34107 18788 34152 18816
rect 34146 18776 34152 18788
rect 34204 18776 34210 18828
rect 40218 18816 40224 18828
rect 37568 18788 40224 18816
rect 30837 18751 30895 18757
rect 30837 18717 30849 18751
rect 30883 18717 30895 18751
rect 30837 18711 30895 18717
rect 30929 18751 30987 18757
rect 30929 18717 30941 18751
rect 30975 18717 30987 18751
rect 31110 18748 31116 18760
rect 31071 18720 31116 18748
rect 30929 18711 30987 18717
rect 20898 18640 20904 18692
rect 20956 18680 20962 18692
rect 21054 18683 21112 18689
rect 21054 18680 21066 18683
rect 20956 18652 21066 18680
rect 20956 18640 20962 18652
rect 21054 18649 21066 18652
rect 21100 18649 21112 18683
rect 21054 18643 21112 18649
rect 21542 18640 21548 18692
rect 21600 18680 21606 18692
rect 23017 18683 23075 18689
rect 23017 18680 23029 18683
rect 21600 18652 23029 18680
rect 21600 18640 21606 18652
rect 23017 18649 23029 18652
rect 23063 18649 23075 18683
rect 23017 18643 23075 18649
rect 26145 18683 26203 18689
rect 26145 18649 26157 18683
rect 26191 18680 26203 18683
rect 26326 18680 26332 18692
rect 26191 18652 26332 18680
rect 26191 18649 26203 18652
rect 26145 18643 26203 18649
rect 26326 18640 26332 18652
rect 26384 18640 26390 18692
rect 26620 18680 26648 18708
rect 27062 18680 27068 18692
rect 26620 18652 27068 18680
rect 27062 18640 27068 18652
rect 27120 18680 27126 18692
rect 27433 18683 27491 18689
rect 27433 18680 27445 18683
rect 27120 18652 27445 18680
rect 27120 18640 27126 18652
rect 27433 18649 27445 18652
rect 27479 18649 27491 18683
rect 27433 18643 27491 18649
rect 29914 18640 29920 18692
rect 29972 18680 29978 18692
rect 29972 18652 30017 18680
rect 29972 18640 29978 18652
rect 24302 18612 24308 18624
rect 20640 18584 24308 18612
rect 17828 18572 17834 18584
rect 24302 18572 24308 18584
rect 24360 18572 24366 18624
rect 25774 18612 25780 18624
rect 25735 18584 25780 18612
rect 25774 18572 25780 18584
rect 25832 18572 25838 18624
rect 26050 18572 26056 18624
rect 26108 18612 26114 18624
rect 26605 18615 26663 18621
rect 26605 18612 26617 18615
rect 26108 18584 26617 18612
rect 26108 18572 26114 18584
rect 26605 18581 26617 18584
rect 26651 18612 26663 18615
rect 27522 18612 27528 18624
rect 26651 18584 27528 18612
rect 26651 18581 26663 18584
rect 26605 18575 26663 18581
rect 27522 18572 27528 18584
rect 27580 18572 27586 18624
rect 30006 18572 30012 18624
rect 30064 18612 30070 18624
rect 30944 18612 30972 18711
rect 31110 18708 31116 18720
rect 31168 18708 31174 18760
rect 32125 18751 32183 18757
rect 32125 18717 32137 18751
rect 32171 18748 32183 18751
rect 32674 18748 32680 18760
rect 32171 18720 32680 18748
rect 32171 18717 32183 18720
rect 32125 18711 32183 18717
rect 32674 18708 32680 18720
rect 32732 18708 32738 18760
rect 35986 18708 35992 18760
rect 36044 18748 36050 18760
rect 36081 18751 36139 18757
rect 36081 18748 36093 18751
rect 36044 18720 36093 18748
rect 36044 18708 36050 18720
rect 36081 18717 36093 18720
rect 36127 18717 36139 18751
rect 36262 18748 36268 18760
rect 36223 18720 36268 18748
rect 36081 18711 36139 18717
rect 36262 18708 36268 18720
rect 36320 18708 36326 18760
rect 36449 18751 36507 18757
rect 36449 18717 36461 18751
rect 36495 18748 36507 18751
rect 36906 18748 36912 18760
rect 36495 18720 36912 18748
rect 36495 18717 36507 18720
rect 36449 18711 36507 18717
rect 36906 18708 36912 18720
rect 36964 18708 36970 18760
rect 37274 18708 37280 18760
rect 37332 18748 37338 18760
rect 37568 18757 37596 18788
rect 40218 18776 40224 18788
rect 40276 18776 40282 18828
rect 37461 18751 37519 18757
rect 37461 18748 37473 18751
rect 37332 18720 37473 18748
rect 37332 18708 37338 18720
rect 37461 18717 37473 18720
rect 37507 18717 37519 18751
rect 37461 18711 37519 18717
rect 37553 18751 37611 18757
rect 37553 18717 37565 18751
rect 37599 18717 37611 18751
rect 37553 18711 37611 18717
rect 37829 18751 37887 18757
rect 37829 18717 37841 18751
rect 37875 18748 37887 18751
rect 40126 18748 40132 18760
rect 37875 18720 40132 18748
rect 37875 18717 37887 18720
rect 37829 18711 37887 18717
rect 40126 18708 40132 18720
rect 40184 18708 40190 18760
rect 58158 18748 58164 18760
rect 58119 18720 58164 18748
rect 58158 18708 58164 18720
rect 58216 18708 58222 18760
rect 31941 18683 31999 18689
rect 31941 18649 31953 18683
rect 31987 18680 31999 18683
rect 33318 18680 33324 18692
rect 31987 18652 33324 18680
rect 31987 18649 31999 18652
rect 31941 18643 31999 18649
rect 33318 18640 33324 18652
rect 33376 18640 33382 18692
rect 33502 18640 33508 18692
rect 33560 18680 33566 18692
rect 33882 18683 33940 18689
rect 33882 18680 33894 18683
rect 33560 18652 33894 18680
rect 33560 18640 33566 18652
rect 33882 18649 33894 18652
rect 33928 18649 33940 18683
rect 33882 18643 33940 18649
rect 36173 18683 36231 18689
rect 36173 18649 36185 18683
rect 36219 18649 36231 18683
rect 37642 18680 37648 18692
rect 37603 18652 37648 18680
rect 36173 18643 36231 18649
rect 30064 18584 30972 18612
rect 32309 18615 32367 18621
rect 30064 18572 30070 18584
rect 32309 18581 32321 18615
rect 32355 18612 32367 18615
rect 32582 18612 32588 18624
rect 32355 18584 32588 18612
rect 32355 18581 32367 18584
rect 32309 18575 32367 18581
rect 32582 18572 32588 18584
rect 32640 18572 32646 18624
rect 36188 18612 36216 18643
rect 37642 18640 37648 18652
rect 37700 18640 37706 18692
rect 38102 18640 38108 18692
rect 38160 18680 38166 18692
rect 39945 18683 40003 18689
rect 39945 18680 39957 18683
rect 38160 18652 39957 18680
rect 38160 18640 38166 18652
rect 39945 18649 39957 18652
rect 39991 18649 40003 18683
rect 39945 18643 40003 18649
rect 39390 18612 39396 18624
rect 36188 18584 39396 18612
rect 39390 18572 39396 18584
rect 39448 18572 39454 18624
rect 40313 18615 40371 18621
rect 40313 18581 40325 18615
rect 40359 18612 40371 18615
rect 40770 18612 40776 18624
rect 40359 18584 40776 18612
rect 40359 18581 40371 18584
rect 40313 18575 40371 18581
rect 40770 18572 40776 18584
rect 40828 18572 40834 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 6825 18411 6883 18417
rect 6825 18377 6837 18411
rect 6871 18408 6883 18411
rect 6914 18408 6920 18420
rect 6871 18380 6920 18408
rect 6871 18377 6883 18380
rect 6825 18371 6883 18377
rect 6914 18368 6920 18380
rect 6972 18368 6978 18420
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 8481 18411 8539 18417
rect 8481 18408 8493 18411
rect 8352 18380 8493 18408
rect 8352 18368 8358 18380
rect 8481 18377 8493 18380
rect 8527 18377 8539 18411
rect 18046 18408 18052 18420
rect 18007 18380 18052 18408
rect 8481 18371 8539 18377
rect 18046 18368 18052 18380
rect 18104 18368 18110 18420
rect 20898 18408 20904 18420
rect 18156 18380 19840 18408
rect 20859 18380 20904 18408
rect 2774 18340 2780 18352
rect 2240 18312 2780 18340
rect 2240 18281 2268 18312
rect 2774 18300 2780 18312
rect 2832 18300 2838 18352
rect 5074 18340 5080 18352
rect 4172 18312 5080 18340
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18241 2283 18275
rect 2225 18235 2283 18241
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 3145 18275 3203 18281
rect 3145 18272 3157 18275
rect 2547 18244 3157 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 3145 18241 3157 18244
rect 3191 18241 3203 18275
rect 3145 18235 3203 18241
rect 2332 18204 2360 18235
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4172 18281 4200 18312
rect 5074 18300 5080 18312
rect 5132 18300 5138 18352
rect 7650 18340 7656 18352
rect 7024 18312 7656 18340
rect 4157 18275 4215 18281
rect 4157 18272 4169 18275
rect 4120 18244 4169 18272
rect 4120 18232 4126 18244
rect 4157 18241 4169 18244
rect 4203 18241 4215 18275
rect 4157 18235 4215 18241
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18272 4307 18275
rect 4614 18272 4620 18284
rect 4295 18244 4620 18272
rect 4295 18241 4307 18244
rect 4249 18235 4307 18241
rect 4614 18232 4620 18244
rect 4672 18232 4678 18284
rect 5445 18275 5503 18281
rect 5445 18241 5457 18275
rect 5491 18272 5503 18275
rect 5902 18272 5908 18284
rect 5491 18244 5908 18272
rect 5491 18241 5503 18244
rect 5445 18235 5503 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 7024 18281 7052 18312
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 9852 18343 9910 18349
rect 9852 18309 9864 18343
rect 9898 18340 9910 18343
rect 11514 18340 11520 18352
rect 9898 18312 11520 18340
rect 9898 18309 9910 18312
rect 9852 18303 9910 18309
rect 11514 18300 11520 18312
rect 11572 18300 11578 18352
rect 13722 18300 13728 18352
rect 13780 18340 13786 18352
rect 18156 18340 18184 18380
rect 13780 18312 18184 18340
rect 18233 18343 18291 18349
rect 13780 18300 13786 18312
rect 18233 18309 18245 18343
rect 18279 18340 18291 18343
rect 18966 18340 18972 18352
rect 18279 18312 18972 18340
rect 18279 18309 18291 18312
rect 18233 18303 18291 18309
rect 18966 18300 18972 18312
rect 19024 18300 19030 18352
rect 19812 18349 19840 18380
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 22649 18411 22707 18417
rect 22649 18408 22661 18411
rect 22204 18380 22661 18408
rect 19797 18343 19855 18349
rect 19797 18309 19809 18343
rect 19843 18340 19855 18343
rect 21821 18343 21879 18349
rect 21821 18340 21833 18343
rect 19843 18312 20392 18340
rect 19843 18309 19855 18312
rect 19797 18303 19855 18309
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18241 7067 18275
rect 7374 18272 7380 18284
rect 7335 18244 7380 18272
rect 7009 18235 7067 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 7561 18275 7619 18281
rect 7561 18241 7573 18275
rect 7607 18272 7619 18275
rect 8110 18272 8116 18284
rect 7607 18244 8116 18272
rect 7607 18241 7619 18244
rect 7561 18235 7619 18241
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 9582 18272 9588 18284
rect 9543 18244 9588 18272
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 11054 18232 11060 18284
rect 11112 18272 11118 18284
rect 11885 18275 11943 18281
rect 11885 18272 11897 18275
rect 11112 18244 11897 18272
rect 11112 18232 11118 18244
rect 11885 18241 11897 18244
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18272 14335 18275
rect 14366 18272 14372 18284
rect 14323 18244 14372 18272
rect 14323 18241 14335 18244
rect 14277 18235 14335 18241
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 14461 18235 14519 18241
rect 18248 18244 18429 18272
rect 4433 18207 4491 18213
rect 2332 18176 2774 18204
rect 2746 18136 2774 18176
rect 4433 18173 4445 18207
rect 4479 18204 4491 18207
rect 4798 18204 4804 18216
rect 4479 18176 4804 18204
rect 4479 18173 4491 18176
rect 4433 18167 4491 18173
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 7190 18204 7196 18216
rect 7151 18176 7196 18204
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 7285 18207 7343 18213
rect 7285 18173 7297 18207
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 3789 18139 3847 18145
rect 3789 18136 3801 18139
rect 2746 18108 3801 18136
rect 3789 18105 3801 18108
rect 3835 18105 3847 18139
rect 3789 18099 3847 18105
rect 5534 18096 5540 18148
rect 5592 18136 5598 18148
rect 7300 18136 7328 18167
rect 12710 18164 12716 18216
rect 12768 18204 12774 18216
rect 14476 18204 14504 18235
rect 12768 18176 14504 18204
rect 12768 18164 12774 18176
rect 18248 18148 18276 18244
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 20257 18275 20315 18281
rect 20257 18241 20269 18275
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 18322 18164 18328 18216
rect 18380 18204 18386 18216
rect 20272 18204 20300 18235
rect 18380 18176 20300 18204
rect 20364 18204 20392 18312
rect 20456 18312 21833 18340
rect 20456 18281 20484 18312
rect 21821 18309 21833 18312
rect 21867 18309 21879 18343
rect 22002 18340 22008 18352
rect 21963 18312 22008 18340
rect 21821 18303 21879 18309
rect 22002 18300 22008 18312
rect 22060 18300 22066 18352
rect 22204 18349 22232 18380
rect 22649 18377 22661 18380
rect 22695 18377 22707 18411
rect 22649 18371 22707 18377
rect 27522 18368 27528 18420
rect 27580 18408 27586 18420
rect 31481 18411 31539 18417
rect 31481 18408 31493 18411
rect 27580 18380 31493 18408
rect 27580 18368 27586 18380
rect 31481 18377 31493 18380
rect 31527 18408 31539 18411
rect 31846 18408 31852 18420
rect 31527 18380 31852 18408
rect 31527 18377 31539 18380
rect 31481 18371 31539 18377
rect 31846 18368 31852 18380
rect 31904 18408 31910 18420
rect 32122 18408 32128 18420
rect 31904 18380 32128 18408
rect 31904 18368 31910 18380
rect 32122 18368 32128 18380
rect 32180 18368 32186 18420
rect 33045 18411 33103 18417
rect 33045 18377 33057 18411
rect 33091 18408 33103 18411
rect 33226 18408 33232 18420
rect 33091 18380 33232 18408
rect 33091 18377 33103 18380
rect 33045 18371 33103 18377
rect 33226 18368 33232 18380
rect 33284 18368 33290 18420
rect 33502 18408 33508 18420
rect 33463 18380 33508 18408
rect 33502 18368 33508 18380
rect 33560 18368 33566 18420
rect 34701 18411 34759 18417
rect 34701 18408 34713 18411
rect 33796 18380 34713 18408
rect 22189 18343 22247 18349
rect 22189 18309 22201 18343
rect 22235 18309 22247 18343
rect 22189 18303 22247 18309
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18241 20499 18275
rect 20441 18235 20499 18241
rect 20530 18232 20536 18284
rect 20588 18272 20594 18284
rect 20671 18275 20729 18281
rect 20588 18244 20633 18272
rect 20588 18232 20594 18244
rect 20671 18241 20683 18275
rect 20717 18272 20729 18275
rect 20717 18244 20852 18272
rect 20717 18241 20729 18244
rect 20671 18235 20729 18241
rect 20824 18204 20852 18244
rect 20364 18176 20852 18204
rect 18380 18164 18386 18176
rect 11790 18136 11796 18148
rect 5592 18108 7328 18136
rect 10520 18108 11796 18136
rect 5592 18096 5598 18108
rect 2958 18068 2964 18080
rect 2919 18040 2964 18068
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 5626 18068 5632 18080
rect 5539 18040 5632 18068
rect 5626 18028 5632 18040
rect 5684 18068 5690 18080
rect 10520 18068 10548 18108
rect 11790 18096 11796 18108
rect 11848 18136 11854 18148
rect 16298 18136 16304 18148
rect 11848 18108 16304 18136
rect 11848 18096 11854 18108
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 18230 18136 18236 18148
rect 18143 18108 18236 18136
rect 18230 18096 18236 18108
rect 18288 18136 18294 18148
rect 22204 18136 22232 18303
rect 24210 18300 24216 18352
rect 24268 18340 24274 18352
rect 24762 18340 24768 18352
rect 24268 18312 24768 18340
rect 24268 18300 24274 18312
rect 24762 18300 24768 18312
rect 24820 18300 24826 18352
rect 24857 18343 24915 18349
rect 24857 18309 24869 18343
rect 24903 18340 24915 18343
rect 26602 18340 26608 18352
rect 24903 18312 26608 18340
rect 24903 18309 24915 18312
rect 24857 18303 24915 18309
rect 26602 18300 26608 18312
rect 26660 18300 26666 18352
rect 29638 18300 29644 18352
rect 29696 18340 29702 18352
rect 33796 18340 33824 18380
rect 34701 18377 34713 18380
rect 34747 18408 34759 18411
rect 37918 18408 37924 18420
rect 34747 18380 37924 18408
rect 34747 18377 34759 18380
rect 34701 18371 34759 18377
rect 37918 18368 37924 18380
rect 37976 18368 37982 18420
rect 40126 18408 40132 18420
rect 40087 18380 40132 18408
rect 40126 18368 40132 18380
rect 40184 18368 40190 18420
rect 40236 18380 41276 18408
rect 29696 18312 33824 18340
rect 29696 18300 29702 18312
rect 22833 18275 22891 18281
rect 22833 18241 22845 18275
rect 22879 18272 22891 18275
rect 23474 18272 23480 18284
rect 22879 18244 23480 18272
rect 22879 18241 22891 18244
rect 22833 18235 22891 18241
rect 23474 18232 23480 18244
rect 23532 18232 23538 18284
rect 24581 18275 24639 18281
rect 24581 18241 24593 18275
rect 24627 18272 24639 18275
rect 24670 18272 24676 18284
rect 24627 18244 24676 18272
rect 24627 18241 24639 18244
rect 24581 18235 24639 18241
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 24946 18272 24952 18284
rect 24907 18244 24952 18272
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 25777 18275 25835 18281
rect 25777 18241 25789 18275
rect 25823 18272 25835 18275
rect 25958 18272 25964 18284
rect 25823 18244 25964 18272
rect 25823 18241 25835 18244
rect 25777 18235 25835 18241
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 26053 18275 26111 18281
rect 26053 18241 26065 18275
rect 26099 18241 26111 18275
rect 32398 18272 32404 18284
rect 32359 18244 32404 18272
rect 26053 18235 26111 18241
rect 25866 18204 25872 18216
rect 25827 18176 25872 18204
rect 25866 18164 25872 18176
rect 25924 18164 25930 18216
rect 18288 18108 22232 18136
rect 25133 18139 25191 18145
rect 18288 18096 18294 18108
rect 25133 18105 25145 18139
rect 25179 18136 25191 18139
rect 26068 18136 26096 18235
rect 32398 18232 32404 18244
rect 32456 18232 32462 18284
rect 32582 18272 32588 18284
rect 32543 18244 32588 18272
rect 32582 18232 32588 18244
rect 32640 18232 32646 18284
rect 32680 18275 32738 18281
rect 32680 18241 32692 18275
rect 32726 18241 32738 18275
rect 32680 18235 32738 18241
rect 32695 18204 32723 18235
rect 32766 18232 32772 18284
rect 32824 18272 32830 18284
rect 33796 18281 33824 18312
rect 39016 18343 39074 18349
rect 39016 18309 39028 18343
rect 39062 18340 39074 18343
rect 40236 18340 40264 18380
rect 41046 18340 41052 18352
rect 39062 18312 40264 18340
rect 40880 18312 41052 18340
rect 39062 18309 39074 18312
rect 39016 18303 39074 18309
rect 33781 18275 33839 18281
rect 32824 18244 32869 18272
rect 32824 18232 32830 18244
rect 33781 18241 33793 18275
rect 33827 18241 33839 18275
rect 33781 18235 33839 18241
rect 33870 18275 33928 18281
rect 33870 18241 33882 18275
rect 33916 18241 33928 18275
rect 33870 18235 33928 18241
rect 33970 18275 34028 18281
rect 33970 18241 33982 18275
rect 34016 18272 34028 18275
rect 34016 18244 34109 18272
rect 34016 18241 34028 18244
rect 33970 18235 34028 18241
rect 33042 18204 33048 18216
rect 32695 18176 33048 18204
rect 33042 18164 33048 18176
rect 33100 18204 33106 18216
rect 33885 18204 33913 18235
rect 33100 18176 33913 18204
rect 34081 18204 34109 18244
rect 34146 18232 34152 18284
rect 34204 18272 34210 18284
rect 37553 18275 37611 18281
rect 34204 18244 34249 18272
rect 34204 18232 34210 18244
rect 37553 18241 37565 18275
rect 37599 18272 37611 18275
rect 38102 18272 38108 18284
rect 37599 18244 38108 18272
rect 37599 18241 37611 18244
rect 37553 18235 37611 18241
rect 38102 18232 38108 18244
rect 38160 18232 38166 18284
rect 40126 18232 40132 18284
rect 40184 18272 40190 18284
rect 40589 18275 40647 18281
rect 40589 18272 40601 18275
rect 40184 18244 40601 18272
rect 40184 18232 40190 18244
rect 40589 18241 40601 18244
rect 40635 18241 40647 18275
rect 40770 18272 40776 18284
rect 40731 18244 40776 18272
rect 40589 18235 40647 18241
rect 40770 18232 40776 18244
rect 40828 18232 40834 18284
rect 40880 18281 40908 18312
rect 41046 18300 41052 18312
rect 41104 18300 41110 18352
rect 41248 18349 41276 18380
rect 41233 18343 41291 18349
rect 41233 18309 41245 18343
rect 41279 18309 41291 18343
rect 41233 18303 41291 18309
rect 40865 18275 40923 18281
rect 40865 18241 40877 18275
rect 40911 18241 40923 18275
rect 40865 18235 40923 18241
rect 40957 18275 41015 18281
rect 40957 18241 40969 18275
rect 41003 18241 41015 18275
rect 40957 18235 41015 18241
rect 34330 18204 34336 18216
rect 34081 18176 34336 18204
rect 33100 18164 33106 18176
rect 34330 18164 34336 18176
rect 34388 18164 34394 18216
rect 37182 18164 37188 18216
rect 37240 18204 37246 18216
rect 37277 18207 37335 18213
rect 37277 18204 37289 18207
rect 37240 18176 37289 18204
rect 37240 18164 37246 18176
rect 37277 18173 37289 18176
rect 37323 18173 37335 18207
rect 38746 18204 38752 18216
rect 38707 18176 38752 18204
rect 37277 18167 37335 18173
rect 38746 18164 38752 18176
rect 38804 18164 38810 18216
rect 40678 18164 40684 18216
rect 40736 18204 40742 18216
rect 40972 18204 41000 18235
rect 40736 18176 41000 18204
rect 40736 18164 40742 18176
rect 25179 18108 25820 18136
rect 26068 18108 31754 18136
rect 25179 18105 25191 18108
rect 25133 18099 25191 18105
rect 5684 18040 10548 18068
rect 10965 18071 11023 18077
rect 5684 18028 5690 18040
rect 10965 18037 10977 18071
rect 11011 18068 11023 18071
rect 11146 18068 11152 18080
rect 11011 18040 11152 18068
rect 11011 18037 11023 18040
rect 10965 18031 11023 18037
rect 11146 18028 11152 18040
rect 11204 18068 11210 18080
rect 12250 18068 12256 18080
rect 11204 18040 12256 18068
rect 11204 18028 11210 18040
rect 12250 18028 12256 18040
rect 12308 18028 12314 18080
rect 13170 18068 13176 18080
rect 13131 18040 13176 18068
rect 13170 18028 13176 18040
rect 13228 18028 13234 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14093 18071 14151 18077
rect 14093 18068 14105 18071
rect 13872 18040 14105 18068
rect 13872 18028 13878 18040
rect 14093 18037 14105 18040
rect 14139 18037 14151 18071
rect 14093 18031 14151 18037
rect 15562 18028 15568 18080
rect 15620 18068 15626 18080
rect 21174 18068 21180 18080
rect 15620 18040 21180 18068
rect 15620 18028 15626 18040
rect 21174 18028 21180 18040
rect 21232 18028 21238 18080
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 25792 18077 25820 18108
rect 25593 18071 25651 18077
rect 25593 18068 25605 18071
rect 22244 18040 25605 18068
rect 22244 18028 22250 18040
rect 25593 18037 25605 18040
rect 25639 18037 25651 18071
rect 25593 18031 25651 18037
rect 25777 18071 25835 18077
rect 25777 18037 25789 18071
rect 25823 18037 25835 18071
rect 25777 18031 25835 18037
rect 27062 18028 27068 18080
rect 27120 18068 27126 18080
rect 27157 18071 27215 18077
rect 27157 18068 27169 18071
rect 27120 18040 27169 18068
rect 27120 18028 27126 18040
rect 27157 18037 27169 18040
rect 27203 18037 27215 18071
rect 31726 18068 31754 18108
rect 32122 18096 32128 18148
rect 32180 18136 32186 18148
rect 32766 18136 32772 18148
rect 32180 18108 32772 18136
rect 32180 18096 32186 18108
rect 32766 18096 32772 18108
rect 32824 18136 32830 18148
rect 38654 18136 38660 18148
rect 32824 18108 38660 18136
rect 32824 18096 32830 18108
rect 38654 18096 38660 18108
rect 38712 18096 38718 18148
rect 33594 18068 33600 18080
rect 31726 18040 33600 18068
rect 27157 18031 27215 18037
rect 33594 18028 33600 18040
rect 33652 18028 33658 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 5353 17867 5411 17873
rect 5353 17833 5365 17867
rect 5399 17864 5411 17867
rect 5534 17864 5540 17876
rect 5399 17836 5540 17864
rect 5399 17833 5411 17836
rect 5353 17827 5411 17833
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 6052 17836 7113 17864
rect 6052 17824 6058 17836
rect 7101 17833 7113 17836
rect 7147 17864 7159 17867
rect 13262 17864 13268 17876
rect 7147 17836 13268 17864
rect 7147 17833 7159 17836
rect 7101 17827 7159 17833
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 14366 17824 14372 17876
rect 14424 17864 14430 17876
rect 15473 17867 15531 17873
rect 15473 17864 15485 17867
rect 14424 17836 15485 17864
rect 14424 17824 14430 17836
rect 15473 17833 15485 17836
rect 15519 17833 15531 17867
rect 16574 17864 16580 17876
rect 15473 17827 15531 17833
rect 15580 17836 16580 17864
rect 13170 17756 13176 17808
rect 13228 17796 13234 17808
rect 13228 17768 14136 17796
rect 13228 17756 13234 17768
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 5077 17731 5135 17737
rect 5077 17728 5089 17731
rect 4764 17700 5089 17728
rect 4764 17688 4770 17700
rect 5077 17697 5089 17700
rect 5123 17697 5135 17731
rect 12802 17728 12808 17740
rect 5077 17691 5135 17697
rect 12176 17700 12808 17728
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17660 5227 17663
rect 5534 17660 5540 17672
rect 5215 17632 5540 17660
rect 5215 17629 5227 17632
rect 5169 17623 5227 17629
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 12176 17669 12204 17700
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 13814 17728 13820 17740
rect 13096 17700 13820 17728
rect 12069 17663 12127 17669
rect 12069 17629 12081 17663
rect 12115 17629 12127 17663
rect 12069 17623 12127 17629
rect 12161 17663 12219 17669
rect 12161 17629 12173 17663
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17660 12311 17663
rect 12342 17660 12348 17672
rect 12299 17632 12348 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 7009 17595 7067 17601
rect 7009 17561 7021 17595
rect 7055 17561 7067 17595
rect 7009 17555 7067 17561
rect 3881 17527 3939 17533
rect 3881 17493 3893 17527
rect 3927 17524 3939 17527
rect 4062 17524 4068 17536
rect 3927 17496 4068 17524
rect 3927 17493 3939 17496
rect 3881 17487 3939 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 4709 17527 4767 17533
rect 4709 17493 4721 17527
rect 4755 17524 4767 17527
rect 5718 17524 5724 17536
rect 4755 17496 5724 17524
rect 4755 17493 4767 17496
rect 4709 17487 4767 17493
rect 5718 17484 5724 17496
rect 5776 17484 5782 17536
rect 5902 17524 5908 17536
rect 5863 17496 5908 17524
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 6270 17484 6276 17536
rect 6328 17524 6334 17536
rect 6365 17527 6423 17533
rect 6365 17524 6377 17527
rect 6328 17496 6377 17524
rect 6328 17484 6334 17496
rect 6365 17493 6377 17496
rect 6411 17524 6423 17527
rect 6822 17524 6828 17536
rect 6411 17496 6828 17524
rect 6411 17493 6423 17496
rect 6365 17487 6423 17493
rect 6822 17484 6828 17496
rect 6880 17524 6886 17536
rect 7024 17524 7052 17555
rect 7650 17524 7656 17536
rect 6880 17496 7052 17524
rect 7611 17496 7656 17524
rect 6880 17484 6886 17496
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 11054 17484 11060 17536
rect 11112 17524 11118 17536
rect 11241 17527 11299 17533
rect 11241 17524 11253 17527
rect 11112 17496 11253 17524
rect 11112 17484 11118 17496
rect 11241 17493 11253 17496
rect 11287 17493 11299 17527
rect 11790 17524 11796 17536
rect 11751 17496 11796 17524
rect 11241 17487 11299 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 12084 17524 12112 17623
rect 12176 17592 12204 17623
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17660 12495 17663
rect 12897 17663 12955 17669
rect 12897 17660 12909 17663
rect 12483 17632 12909 17660
rect 12483 17629 12495 17632
rect 12437 17623 12495 17629
rect 12897 17629 12909 17632
rect 12943 17660 12955 17663
rect 12986 17660 12992 17672
rect 12943 17632 12992 17660
rect 12943 17629 12955 17632
rect 12897 17623 12955 17629
rect 12986 17620 12992 17632
rect 13044 17620 13050 17672
rect 13096 17669 13124 17700
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 14108 17737 14136 17768
rect 14093 17731 14151 17737
rect 14093 17697 14105 17731
rect 14139 17697 14151 17731
rect 14093 17691 14151 17697
rect 13081 17663 13139 17669
rect 13081 17629 13093 17663
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 13173 17663 13231 17669
rect 13173 17629 13185 17663
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 13188 17592 13216 17623
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 15580 17660 15608 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 25498 17824 25504 17876
rect 25556 17864 25562 17876
rect 25869 17867 25927 17873
rect 25869 17864 25881 17867
rect 25556 17836 25881 17864
rect 25556 17824 25562 17836
rect 25869 17833 25881 17836
rect 25915 17833 25927 17867
rect 26602 17864 26608 17876
rect 26563 17836 26608 17864
rect 25869 17827 25927 17833
rect 26602 17824 26608 17836
rect 26660 17824 26666 17876
rect 33045 17867 33103 17873
rect 33045 17833 33057 17867
rect 33091 17864 33103 17867
rect 34330 17864 34336 17876
rect 33091 17836 34336 17864
rect 33091 17833 33103 17836
rect 33045 17827 33103 17833
rect 34330 17824 34336 17836
rect 34388 17824 34394 17876
rect 39117 17867 39175 17873
rect 39117 17833 39129 17867
rect 39163 17864 39175 17867
rect 40586 17864 40592 17876
rect 39163 17836 40592 17864
rect 39163 17833 39175 17836
rect 39117 17827 39175 17833
rect 40586 17824 40592 17836
rect 40644 17824 40650 17876
rect 18325 17799 18383 17805
rect 18325 17796 18337 17799
rect 13320 17632 15608 17660
rect 16224 17768 18337 17796
rect 13320 17620 13326 17632
rect 12176 17564 13216 17592
rect 13541 17595 13599 17601
rect 13541 17561 13553 17595
rect 13587 17592 13599 17595
rect 14338 17595 14396 17601
rect 14338 17592 14350 17595
rect 13587 17564 14350 17592
rect 13587 17561 13599 17564
rect 13541 17555 13599 17561
rect 14338 17561 14350 17564
rect 14384 17561 14396 17595
rect 14338 17555 14396 17561
rect 15010 17552 15016 17604
rect 15068 17592 15074 17604
rect 16224 17592 16252 17768
rect 18325 17765 18337 17768
rect 18371 17796 18383 17799
rect 18782 17796 18788 17808
rect 18371 17768 18788 17796
rect 18371 17765 18383 17768
rect 18325 17759 18383 17765
rect 18782 17756 18788 17768
rect 18840 17756 18846 17808
rect 37921 17799 37979 17805
rect 37921 17765 37933 17799
rect 37967 17796 37979 17799
rect 40034 17796 40040 17808
rect 37967 17768 40040 17796
rect 37967 17765 37979 17768
rect 37921 17759 37979 17765
rect 40034 17756 40040 17768
rect 40092 17796 40098 17808
rect 41046 17796 41052 17808
rect 40092 17768 41052 17796
rect 40092 17756 40098 17768
rect 41046 17756 41052 17768
rect 41104 17756 41110 17808
rect 20806 17688 20812 17740
rect 20864 17728 20870 17740
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 20864 17700 21373 17728
rect 20864 17688 20870 17700
rect 21361 17697 21373 17700
rect 21407 17697 21419 17731
rect 21361 17691 21419 17697
rect 33410 17688 33416 17740
rect 33468 17728 33474 17740
rect 34146 17728 34152 17740
rect 33468 17700 34152 17728
rect 33468 17688 33474 17700
rect 34146 17688 34152 17700
rect 34204 17688 34210 17740
rect 38654 17688 38660 17740
rect 38712 17728 38718 17740
rect 40405 17731 40463 17737
rect 40405 17728 40417 17731
rect 38712 17700 40417 17728
rect 38712 17688 38718 17700
rect 40405 17697 40417 17700
rect 40451 17728 40463 17731
rect 40678 17728 40684 17740
rect 40451 17700 40684 17728
rect 40451 17697 40463 17700
rect 40405 17691 40463 17697
rect 40678 17688 40684 17700
rect 40736 17688 40742 17740
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 15068 17564 16252 17592
rect 16408 17632 17141 17660
rect 15068 17552 15074 17564
rect 16301 17527 16359 17533
rect 16301 17524 16313 17527
rect 11940 17496 16313 17524
rect 11940 17484 11946 17496
rect 16301 17493 16313 17496
rect 16347 17524 16359 17527
rect 16408 17524 16436 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 17236 17592 17264 17623
rect 17310 17620 17316 17672
rect 17368 17660 17374 17672
rect 17497 17663 17555 17669
rect 17368 17632 17413 17660
rect 17368 17620 17374 17632
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 17954 17660 17960 17672
rect 17543 17632 17960 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 17954 17620 17960 17632
rect 18012 17660 18018 17672
rect 19150 17660 19156 17672
rect 18012 17632 19156 17660
rect 18012 17620 18018 17632
rect 19150 17620 19156 17632
rect 19208 17620 19214 17672
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 24118 17660 24124 17672
rect 20404 17632 24124 17660
rect 20404 17620 20410 17632
rect 24118 17620 24124 17632
rect 24176 17620 24182 17672
rect 24489 17663 24547 17669
rect 24489 17629 24501 17663
rect 24535 17660 24547 17663
rect 26510 17660 26516 17672
rect 24535 17632 26516 17660
rect 24535 17629 24547 17632
rect 24489 17623 24547 17629
rect 26510 17620 26516 17632
rect 26568 17620 26574 17672
rect 27430 17620 27436 17672
rect 27488 17660 27494 17672
rect 27985 17663 28043 17669
rect 27985 17660 27997 17663
rect 27488 17632 27997 17660
rect 27488 17620 27494 17632
rect 27985 17629 27997 17632
rect 28031 17629 28043 17663
rect 27985 17623 28043 17629
rect 28810 17620 28816 17672
rect 28868 17660 28874 17672
rect 31021 17663 31079 17669
rect 31021 17660 31033 17663
rect 28868 17632 31033 17660
rect 28868 17620 28874 17632
rect 31021 17629 31033 17632
rect 31067 17629 31079 17663
rect 32858 17660 32864 17672
rect 32819 17632 32864 17660
rect 31021 17623 31079 17629
rect 32858 17620 32864 17632
rect 32916 17620 32922 17672
rect 33686 17660 33692 17672
rect 33647 17632 33692 17660
rect 33686 17620 33692 17632
rect 33744 17620 33750 17672
rect 38930 17660 38936 17672
rect 38891 17632 38936 17660
rect 38930 17620 38936 17632
rect 38988 17620 38994 17672
rect 17770 17592 17776 17604
rect 17236 17564 17776 17592
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 21174 17552 21180 17604
rect 21232 17592 21238 17604
rect 21606 17595 21664 17601
rect 21606 17592 21618 17595
rect 21232 17564 21618 17592
rect 21232 17552 21238 17564
rect 21606 17561 21618 17564
rect 21652 17561 21664 17595
rect 21606 17555 21664 17561
rect 24756 17595 24814 17601
rect 24756 17561 24768 17595
rect 24802 17592 24814 17595
rect 25682 17592 25688 17604
rect 24802 17564 25688 17592
rect 24802 17561 24814 17564
rect 24756 17555 24814 17561
rect 25682 17552 25688 17564
rect 25740 17552 25746 17604
rect 26970 17552 26976 17604
rect 27028 17592 27034 17604
rect 27718 17595 27776 17601
rect 27718 17592 27730 17595
rect 27028 17564 27730 17592
rect 27028 17552 27034 17564
rect 27718 17561 27730 17564
rect 27764 17561 27776 17595
rect 32677 17595 32735 17601
rect 32677 17592 32689 17595
rect 27718 17555 27776 17561
rect 31726 17564 32689 17592
rect 16347 17496 16436 17524
rect 16853 17527 16911 17533
rect 16347 17493 16359 17496
rect 16301 17487 16359 17493
rect 16853 17493 16865 17527
rect 16899 17524 16911 17527
rect 16942 17524 16948 17536
rect 16899 17496 16948 17524
rect 16899 17493 16911 17496
rect 16853 17487 16911 17493
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 21818 17484 21824 17536
rect 21876 17524 21882 17536
rect 22741 17527 22799 17533
rect 22741 17524 22753 17527
rect 21876 17496 22753 17524
rect 21876 17484 21882 17496
rect 22741 17493 22753 17496
rect 22787 17493 22799 17527
rect 22741 17487 22799 17493
rect 31205 17527 31263 17533
rect 31205 17493 31217 17527
rect 31251 17524 31263 17527
rect 31726 17524 31754 17564
rect 32677 17561 32689 17564
rect 32723 17592 32735 17595
rect 33318 17592 33324 17604
rect 32723 17564 33324 17592
rect 32723 17561 32735 17564
rect 32677 17555 32735 17561
rect 33318 17552 33324 17564
rect 33376 17592 33382 17604
rect 33505 17595 33563 17601
rect 33505 17592 33517 17595
rect 33376 17564 33517 17592
rect 33376 17552 33382 17564
rect 33505 17561 33517 17564
rect 33551 17561 33563 17595
rect 36262 17592 36268 17604
rect 36223 17564 36268 17592
rect 33505 17555 33563 17561
rect 36262 17552 36268 17564
rect 36320 17552 36326 17604
rect 36449 17595 36507 17601
rect 36449 17561 36461 17595
rect 36495 17592 36507 17595
rect 37182 17592 37188 17604
rect 36495 17564 37188 17592
rect 36495 17561 36507 17564
rect 36449 17555 36507 17561
rect 37182 17552 37188 17564
rect 37240 17552 37246 17604
rect 37737 17595 37795 17601
rect 37737 17561 37749 17595
rect 37783 17592 37795 17595
rect 37826 17592 37832 17604
rect 37783 17564 37832 17592
rect 37783 17561 37795 17564
rect 37737 17555 37795 17561
rect 37826 17552 37832 17564
rect 37884 17552 37890 17604
rect 31251 17496 31754 17524
rect 31251 17493 31263 17496
rect 31205 17487 31263 17493
rect 33594 17484 33600 17536
rect 33652 17524 33658 17536
rect 33873 17527 33931 17533
rect 33873 17524 33885 17527
rect 33652 17496 33885 17524
rect 33652 17484 33658 17496
rect 33873 17493 33885 17496
rect 33919 17493 33931 17527
rect 33873 17487 33931 17493
rect 36081 17527 36139 17533
rect 36081 17493 36093 17527
rect 36127 17524 36139 17527
rect 36170 17524 36176 17536
rect 36127 17496 36176 17524
rect 36127 17493 36139 17496
rect 36081 17487 36139 17493
rect 36170 17484 36176 17496
rect 36228 17484 36234 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 11701 17323 11759 17329
rect 11701 17320 11713 17323
rect 5500 17292 11713 17320
rect 5500 17280 5506 17292
rect 11701 17289 11713 17292
rect 11747 17320 11759 17323
rect 11882 17320 11888 17332
rect 11747 17292 11888 17320
rect 11747 17289 11759 17292
rect 11701 17283 11759 17289
rect 11882 17280 11888 17292
rect 11940 17280 11946 17332
rect 12342 17320 12348 17332
rect 12303 17292 12348 17320
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 13262 17320 13268 17332
rect 13223 17292 13268 17320
rect 13262 17280 13268 17292
rect 13320 17280 13326 17332
rect 13906 17320 13912 17332
rect 13867 17292 13912 17320
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 16022 17280 16028 17332
rect 16080 17320 16086 17332
rect 16080 17292 17724 17320
rect 16080 17280 16086 17292
rect 2860 17255 2918 17261
rect 2860 17221 2872 17255
rect 2906 17252 2918 17255
rect 2958 17252 2964 17264
rect 2906 17224 2964 17252
rect 2906 17221 2918 17224
rect 2860 17215 2918 17221
rect 2958 17212 2964 17224
rect 3016 17212 3022 17264
rect 8938 17252 8944 17264
rect 7944 17224 8944 17252
rect 7006 17144 7012 17196
rect 7064 17184 7070 17196
rect 7944 17193 7972 17224
rect 8938 17212 8944 17224
rect 8996 17212 9002 17264
rect 12529 17255 12587 17261
rect 12529 17221 12541 17255
rect 12575 17252 12587 17255
rect 13078 17252 13084 17264
rect 12575 17224 13084 17252
rect 12575 17221 12587 17224
rect 12529 17215 12587 17221
rect 13078 17212 13084 17224
rect 13136 17212 13142 17264
rect 14185 17255 14243 17261
rect 14185 17221 14197 17255
rect 14231 17252 14243 17255
rect 16574 17252 16580 17264
rect 14231 17224 16580 17252
rect 14231 17221 14243 17224
rect 14185 17215 14243 17221
rect 16574 17212 16580 17224
rect 16632 17212 16638 17264
rect 7561 17187 7619 17193
rect 7561 17184 7573 17187
rect 7064 17156 7573 17184
rect 7064 17144 7070 17156
rect 7561 17153 7573 17156
rect 7607 17153 7619 17187
rect 7561 17147 7619 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 8110 17184 8116 17196
rect 8071 17156 8116 17184
rect 7929 17147 7987 17153
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 12710 17184 12716 17196
rect 12671 17156 12716 17184
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 13998 17144 14004 17196
rect 14056 17193 14062 17196
rect 14056 17187 14105 17193
rect 14056 17153 14059 17187
rect 14093 17153 14105 17187
rect 14274 17184 14280 17196
rect 14235 17156 14280 17184
rect 14056 17147 14105 17153
rect 14056 17144 14062 17147
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 14366 17144 14372 17196
rect 14424 17193 14430 17196
rect 14424 17187 14463 17193
rect 14451 17153 14463 17187
rect 14424 17147 14463 17153
rect 14424 17144 14430 17147
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 15194 17184 15200 17196
rect 14608 17156 14653 17184
rect 14752 17156 15200 17184
rect 14608 17144 14614 17156
rect 1946 17076 1952 17128
rect 2004 17116 2010 17128
rect 2593 17119 2651 17125
rect 2593 17116 2605 17119
rect 2004 17088 2605 17116
rect 2004 17076 2010 17088
rect 2593 17085 2605 17088
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 7190 17076 7196 17128
rect 7248 17116 7254 17128
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7248 17088 7757 17116
rect 7248 17076 7254 17088
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 7834 17076 7840 17128
rect 7892 17116 7898 17128
rect 14752 17116 14780 17156
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15286 17144 15292 17196
rect 15344 17184 15350 17196
rect 16669 17187 16727 17193
rect 15344 17156 15389 17184
rect 15344 17144 15350 17156
rect 16669 17153 16681 17187
rect 16715 17184 16727 17187
rect 16758 17184 16764 17196
rect 16715 17156 16764 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 16942 17193 16948 17196
rect 16936 17184 16948 17193
rect 16903 17156 16948 17184
rect 16936 17147 16948 17156
rect 16942 17144 16948 17147
rect 17000 17144 17006 17196
rect 15010 17116 15016 17128
rect 7892 17088 7937 17116
rect 8036 17088 14780 17116
rect 14971 17088 15016 17116
rect 7892 17076 7898 17088
rect 3878 17008 3884 17060
rect 3936 17048 3942 17060
rect 8036 17048 8064 17088
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 17696 17116 17724 17292
rect 18506 17280 18512 17332
rect 18564 17320 18570 17332
rect 20990 17320 20996 17332
rect 18564 17292 20996 17320
rect 18564 17280 18570 17292
rect 20990 17280 20996 17292
rect 21048 17280 21054 17332
rect 25682 17320 25688 17332
rect 25643 17292 25688 17320
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 26970 17320 26976 17332
rect 26931 17292 26976 17320
rect 26970 17280 26976 17292
rect 27028 17280 27034 17332
rect 27338 17280 27344 17332
rect 27396 17280 27402 17332
rect 32398 17320 32404 17332
rect 27632 17292 32404 17320
rect 17770 17212 17776 17264
rect 17828 17252 17834 17264
rect 17828 17224 18920 17252
rect 17828 17212 17834 17224
rect 18782 17184 18788 17196
rect 18743 17156 18788 17184
rect 18782 17144 18788 17156
rect 18840 17144 18846 17196
rect 18892 17193 18920 17224
rect 21818 17212 21824 17264
rect 21876 17252 21882 17264
rect 22005 17255 22063 17261
rect 22005 17252 22017 17255
rect 21876 17224 22017 17252
rect 21876 17212 21882 17224
rect 22005 17221 22017 17224
rect 22051 17221 22063 17255
rect 22005 17215 22063 17221
rect 22094 17212 22100 17264
rect 22152 17252 22158 17264
rect 22189 17255 22247 17261
rect 22189 17252 22201 17255
rect 22152 17224 22201 17252
rect 22152 17212 22158 17224
rect 22189 17221 22201 17224
rect 22235 17252 22247 17255
rect 22370 17252 22376 17264
rect 22235 17224 22376 17252
rect 22235 17221 22247 17224
rect 22189 17215 22247 17221
rect 22370 17212 22376 17224
rect 22428 17212 22434 17264
rect 25774 17212 25780 17264
rect 25832 17252 25838 17264
rect 27356 17252 27384 17280
rect 25832 17224 26188 17252
rect 25832 17212 25838 17224
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17153 18935 17187
rect 18877 17147 18935 17153
rect 18966 17144 18972 17196
rect 19024 17184 19030 17196
rect 19150 17184 19156 17196
rect 19024 17156 19069 17184
rect 19111 17156 19156 17184
rect 19024 17144 19030 17156
rect 19150 17144 19156 17156
rect 19208 17144 19214 17196
rect 23017 17187 23075 17193
rect 23017 17153 23029 17187
rect 23063 17184 23075 17187
rect 24210 17184 24216 17196
rect 23063 17156 24216 17184
rect 23063 17153 23075 17156
rect 23017 17147 23075 17153
rect 24210 17144 24216 17156
rect 24268 17144 24274 17196
rect 24305 17187 24363 17193
rect 24305 17153 24317 17187
rect 24351 17184 24363 17187
rect 24946 17184 24952 17196
rect 24351 17156 24952 17184
rect 24351 17153 24363 17156
rect 24305 17147 24363 17153
rect 24946 17144 24952 17156
rect 25004 17144 25010 17196
rect 25682 17144 25688 17196
rect 25740 17184 25746 17196
rect 26160 17193 26188 17224
rect 26252 17224 27384 17252
rect 25915 17187 25973 17193
rect 25915 17184 25927 17187
rect 25740 17156 25927 17184
rect 25740 17144 25746 17156
rect 25915 17153 25927 17156
rect 25961 17153 25973 17187
rect 25915 17147 25973 17153
rect 26053 17187 26111 17193
rect 26053 17153 26065 17187
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 26145 17187 26203 17193
rect 26145 17153 26157 17187
rect 26191 17153 26203 17187
rect 26145 17147 26203 17153
rect 20257 17119 20315 17125
rect 20257 17116 20269 17119
rect 17696 17088 20269 17116
rect 20257 17085 20269 17088
rect 20303 17116 20315 17119
rect 20990 17116 20996 17128
rect 20303 17088 20996 17116
rect 20303 17085 20315 17088
rect 20257 17079 20315 17085
rect 20990 17076 20996 17088
rect 21048 17076 21054 17128
rect 22741 17119 22799 17125
rect 22741 17085 22753 17119
rect 22787 17116 22799 17119
rect 22922 17116 22928 17128
rect 22787 17088 22928 17116
rect 22787 17085 22799 17088
rect 22741 17079 22799 17085
rect 22922 17076 22928 17088
rect 22980 17076 22986 17128
rect 24026 17116 24032 17128
rect 23987 17088 24032 17116
rect 24026 17076 24032 17088
rect 24084 17076 24090 17128
rect 26068 17116 26096 17147
rect 26252 17128 26280 17224
rect 27356 17196 27384 17224
rect 26329 17187 26387 17193
rect 26329 17153 26341 17187
rect 26375 17184 26387 17187
rect 26694 17184 26700 17196
rect 26375 17156 26700 17184
rect 26375 17153 26387 17156
rect 26329 17147 26387 17153
rect 26694 17144 26700 17156
rect 26752 17144 26758 17196
rect 27154 17144 27160 17196
rect 27212 17184 27218 17196
rect 27249 17187 27307 17193
rect 27249 17184 27261 17187
rect 27212 17156 27261 17184
rect 27212 17144 27218 17156
rect 27249 17153 27261 17156
rect 27295 17153 27307 17187
rect 27249 17147 27307 17153
rect 27341 17190 27399 17196
rect 27341 17156 27353 17190
rect 27387 17156 27399 17190
rect 27341 17150 27399 17156
rect 27430 17144 27436 17196
rect 27488 17184 27494 17196
rect 27632 17193 27660 17292
rect 32398 17280 32404 17292
rect 32456 17280 32462 17332
rect 36262 17280 36268 17332
rect 36320 17320 36326 17332
rect 36725 17323 36783 17329
rect 36725 17320 36737 17323
rect 36320 17292 36737 17320
rect 36320 17280 36326 17292
rect 36725 17289 36737 17292
rect 36771 17320 36783 17323
rect 37366 17320 37372 17332
rect 36771 17292 37372 17320
rect 36771 17289 36783 17292
rect 36725 17283 36783 17289
rect 37366 17280 37372 17292
rect 37424 17280 37430 17332
rect 39945 17323 40003 17329
rect 39945 17289 39957 17323
rect 39991 17320 40003 17323
rect 40494 17320 40500 17332
rect 39991 17292 40500 17320
rect 39991 17289 40003 17292
rect 39945 17283 40003 17289
rect 40494 17280 40500 17292
rect 40552 17280 40558 17332
rect 29914 17212 29920 17264
rect 29972 17252 29978 17264
rect 30193 17255 30251 17261
rect 30193 17252 30205 17255
rect 29972 17224 30205 17252
rect 29972 17212 29978 17224
rect 30193 17221 30205 17224
rect 30239 17221 30251 17255
rect 30193 17215 30251 17221
rect 33244 17224 33732 17252
rect 27617 17187 27675 17193
rect 27488 17156 27533 17184
rect 27488 17144 27494 17156
rect 27617 17153 27629 17187
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 26234 17116 26240 17128
rect 26068 17088 26240 17116
rect 26234 17076 26240 17088
rect 26292 17076 26298 17128
rect 3936 17020 8064 17048
rect 3936 17008 3942 17020
rect 10870 17008 10876 17060
rect 10928 17048 10934 17060
rect 19334 17048 19340 17060
rect 10928 17020 16160 17048
rect 10928 17008 10934 17020
rect 3973 16983 4031 16989
rect 3973 16949 3985 16983
rect 4019 16980 4031 16983
rect 4614 16980 4620 16992
rect 4019 16952 4620 16980
rect 4019 16949 4031 16952
rect 3973 16943 4031 16949
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 5077 16983 5135 16989
rect 5077 16980 5089 16983
rect 4764 16952 5089 16980
rect 4764 16940 4770 16952
rect 5077 16949 5089 16952
rect 5123 16980 5135 16983
rect 5350 16980 5356 16992
rect 5123 16952 5356 16980
rect 5123 16949 5135 16952
rect 5077 16943 5135 16949
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5721 16983 5779 16989
rect 5721 16949 5733 16983
rect 5767 16980 5779 16983
rect 5902 16980 5908 16992
rect 5767 16952 5908 16980
rect 5767 16949 5779 16952
rect 5721 16943 5779 16949
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 7374 16980 7380 16992
rect 7335 16952 7380 16980
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 16022 16980 16028 16992
rect 9732 16952 16028 16980
rect 9732 16940 9738 16952
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 16132 16980 16160 17020
rect 17604 17020 19340 17048
rect 17604 16980 17632 17020
rect 19334 17008 19340 17020
rect 19392 17008 19398 17060
rect 26712 17048 26740 17144
rect 27632 17048 27660 17147
rect 28994 17144 29000 17196
rect 29052 17184 29058 17196
rect 30009 17187 30067 17193
rect 30009 17184 30021 17187
rect 29052 17156 30021 17184
rect 29052 17144 29058 17156
rect 30009 17153 30021 17156
rect 30055 17153 30067 17187
rect 30009 17147 30067 17153
rect 32401 17187 32459 17193
rect 32401 17153 32413 17187
rect 32447 17184 32459 17187
rect 33042 17184 33048 17196
rect 32447 17156 33048 17184
rect 32447 17153 32459 17156
rect 32401 17147 32459 17153
rect 33042 17144 33048 17156
rect 33100 17184 33106 17196
rect 33244 17184 33272 17224
rect 33410 17184 33416 17196
rect 33100 17156 33272 17184
rect 33371 17156 33416 17184
rect 33100 17144 33106 17156
rect 33410 17144 33416 17156
rect 33468 17144 33474 17196
rect 33594 17184 33600 17196
rect 33555 17156 33600 17184
rect 33594 17144 33600 17156
rect 33652 17144 33658 17196
rect 33704 17193 33732 17224
rect 35618 17193 35624 17196
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17153 33747 17187
rect 33689 17147 33747 17153
rect 33781 17187 33839 17193
rect 33781 17153 33793 17187
rect 33827 17153 33839 17187
rect 33781 17147 33839 17153
rect 35612 17147 35624 17193
rect 35676 17184 35682 17196
rect 35676 17156 35712 17184
rect 32122 17116 32128 17128
rect 32083 17088 32128 17116
rect 32122 17076 32128 17088
rect 32180 17076 32186 17128
rect 26712 17020 27660 17048
rect 28074 17008 28080 17060
rect 28132 17048 28138 17060
rect 28132 17020 30604 17048
rect 28132 17008 28138 17020
rect 16132 16952 17632 16980
rect 18049 16983 18107 16989
rect 18049 16949 18061 16983
rect 18095 16980 18107 16983
rect 18138 16980 18144 16992
rect 18095 16952 18144 16980
rect 18095 16949 18107 16952
rect 18049 16943 18107 16949
rect 18138 16940 18144 16952
rect 18196 16940 18202 16992
rect 18322 16940 18328 16992
rect 18380 16980 18386 16992
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 18380 16952 18521 16980
rect 18380 16940 18386 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18509 16943 18567 16949
rect 21726 16940 21732 16992
rect 21784 16980 21790 16992
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 21784 16952 21833 16980
rect 21784 16940 21790 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 21821 16943 21879 16949
rect 25038 16940 25044 16992
rect 25096 16980 25102 16992
rect 29178 16980 29184 16992
rect 25096 16952 29184 16980
rect 25096 16940 25102 16952
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 30377 16983 30435 16989
rect 30377 16949 30389 16983
rect 30423 16980 30435 16983
rect 30466 16980 30472 16992
rect 30423 16952 30472 16980
rect 30423 16949 30435 16952
rect 30377 16943 30435 16949
rect 30466 16940 30472 16952
rect 30524 16940 30530 16992
rect 30576 16980 30604 17020
rect 31294 17008 31300 17060
rect 31352 17048 31358 17060
rect 33318 17048 33324 17060
rect 31352 17020 33324 17048
rect 31352 17008 31358 17020
rect 33318 17008 33324 17020
rect 33376 17048 33382 17060
rect 33796 17048 33824 17147
rect 35618 17144 35624 17147
rect 35676 17144 35682 17156
rect 39942 17144 39948 17196
rect 40000 17184 40006 17196
rect 40037 17187 40095 17193
rect 40037 17184 40049 17187
rect 40000 17156 40049 17184
rect 40000 17144 40006 17156
rect 40037 17153 40049 17156
rect 40083 17153 40095 17187
rect 40037 17147 40095 17153
rect 34514 17076 34520 17128
rect 34572 17116 34578 17128
rect 35345 17119 35403 17125
rect 35345 17116 35357 17119
rect 34572 17088 35357 17116
rect 34572 17076 34578 17088
rect 35345 17085 35357 17088
rect 35391 17085 35403 17119
rect 35345 17079 35403 17085
rect 58158 17048 58164 17060
rect 33376 17020 33824 17048
rect 33888 17020 35388 17048
rect 58119 17020 58164 17048
rect 33376 17008 33382 17020
rect 33888 16980 33916 17020
rect 34054 16980 34060 16992
rect 30576 16952 33916 16980
rect 34015 16952 34060 16980
rect 34054 16940 34060 16952
rect 34112 16940 34118 16992
rect 35360 16980 35388 17020
rect 58158 17008 58164 17020
rect 58216 17008 58222 17060
rect 36354 16980 36360 16992
rect 35360 16952 36360 16980
rect 36354 16940 36360 16952
rect 36412 16980 36418 16992
rect 38194 16980 38200 16992
rect 36412 16952 38200 16980
rect 36412 16940 36418 16952
rect 38194 16940 38200 16952
rect 38252 16980 38258 16992
rect 40126 16980 40132 16992
rect 38252 16952 40132 16980
rect 38252 16940 38258 16952
rect 40126 16940 40132 16952
rect 40184 16940 40190 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10045 16779 10103 16785
rect 10045 16776 10057 16779
rect 10008 16748 10057 16776
rect 10008 16736 10014 16748
rect 10045 16745 10057 16748
rect 10091 16745 10103 16779
rect 16298 16776 16304 16788
rect 16259 16748 16304 16776
rect 10045 16739 10103 16745
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 17957 16779 18015 16785
rect 17957 16776 17969 16779
rect 17368 16748 17969 16776
rect 17368 16736 17374 16748
rect 17957 16745 17969 16748
rect 18003 16745 18015 16779
rect 17957 16739 18015 16745
rect 18966 16736 18972 16788
rect 19024 16776 19030 16788
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 19024 16748 19257 16776
rect 19024 16736 19030 16748
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 21174 16776 21180 16788
rect 21135 16748 21180 16776
rect 19245 16739 19303 16745
rect 21174 16736 21180 16748
rect 21232 16736 21238 16788
rect 24578 16776 24584 16788
rect 21284 16748 24584 16776
rect 9490 16668 9496 16720
rect 9548 16708 9554 16720
rect 10318 16708 10324 16720
rect 9548 16680 10324 16708
rect 9548 16668 9554 16680
rect 10318 16668 10324 16680
rect 10376 16668 10382 16720
rect 20625 16711 20683 16717
rect 20625 16677 20637 16711
rect 20671 16708 20683 16711
rect 20898 16708 20904 16720
rect 20671 16680 20904 16708
rect 20671 16677 20683 16680
rect 20625 16671 20683 16677
rect 20898 16668 20904 16680
rect 20956 16708 20962 16720
rect 21284 16708 21312 16748
rect 24578 16736 24584 16748
rect 24636 16776 24642 16788
rect 26697 16779 26755 16785
rect 24636 16748 25636 16776
rect 24636 16736 24642 16748
rect 20956 16680 21496 16708
rect 20956 16668 20962 16680
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 5169 16643 5227 16649
rect 5169 16640 5181 16643
rect 4672 16612 5181 16640
rect 4672 16600 4678 16612
rect 5169 16609 5181 16612
rect 5215 16609 5227 16643
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5169 16603 5227 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 8389 16643 8447 16649
rect 8389 16609 8401 16643
rect 8435 16640 8447 16643
rect 9582 16640 9588 16652
rect 8435 16612 9588 16640
rect 8435 16609 8447 16612
rect 8389 16603 8447 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 11238 16640 11244 16652
rect 10244 16612 11244 16640
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 2498 16572 2504 16584
rect 2455 16544 2504 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 5261 16575 5319 16581
rect 5261 16541 5273 16575
rect 5307 16572 5319 16575
rect 5534 16572 5540 16584
rect 5307 16544 5540 16572
rect 5307 16541 5319 16544
rect 5261 16535 5319 16541
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 7374 16532 7380 16584
rect 7432 16572 7438 16584
rect 10244 16581 10272 16612
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 17770 16640 17776 16652
rect 17236 16612 17776 16640
rect 8122 16575 8180 16581
rect 8122 16572 8134 16575
rect 7432 16544 8134 16572
rect 7432 16532 7438 16544
rect 8122 16541 8134 16544
rect 8168 16541 8180 16575
rect 10045 16575 10103 16581
rect 10045 16572 10057 16575
rect 8122 16535 8180 16541
rect 9508 16544 10057 16572
rect 9508 16448 9536 16544
rect 10045 16541 10057 16544
rect 10091 16541 10103 16575
rect 10045 16535 10103 16541
rect 10229 16575 10287 16581
rect 10229 16541 10241 16575
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 10060 16504 10088 16535
rect 16298 16532 16304 16584
rect 16356 16572 16362 16584
rect 17236 16581 17264 16612
rect 17770 16600 17776 16612
rect 17828 16600 17834 16652
rect 17954 16640 17960 16652
rect 17880 16612 17960 16640
rect 17129 16575 17187 16581
rect 17129 16572 17141 16575
rect 16356 16544 17141 16572
rect 16356 16532 16362 16544
rect 17129 16541 17141 16544
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 17313 16575 17371 16581
rect 17313 16541 17325 16575
rect 17359 16572 17371 16575
rect 17402 16572 17408 16584
rect 17359 16544 17408 16572
rect 17359 16541 17371 16544
rect 17313 16535 17371 16541
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16572 17555 16575
rect 17880 16572 17908 16612
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 17543 16544 17908 16572
rect 17543 16541 17555 16544
rect 17497 16535 17555 16541
rect 18046 16532 18052 16584
rect 18104 16572 18110 16584
rect 18230 16572 18236 16584
rect 18104 16544 18236 16572
rect 18104 16532 18110 16544
rect 18230 16532 18236 16544
rect 18288 16572 18294 16584
rect 21468 16581 21496 16680
rect 21542 16668 21548 16720
rect 21600 16668 21606 16720
rect 24486 16668 24492 16720
rect 24544 16708 24550 16720
rect 25406 16708 25412 16720
rect 24544 16680 25412 16708
rect 24544 16668 24550 16680
rect 25406 16668 25412 16680
rect 25464 16668 25470 16720
rect 25608 16717 25636 16748
rect 26697 16745 26709 16779
rect 26743 16776 26755 16779
rect 27430 16776 27436 16788
rect 26743 16748 27436 16776
rect 26743 16745 26755 16748
rect 26697 16739 26755 16745
rect 27430 16736 27436 16748
rect 27488 16736 27494 16788
rect 28902 16736 28908 16788
rect 28960 16776 28966 16788
rect 30558 16776 30564 16788
rect 28960 16748 30564 16776
rect 28960 16736 28966 16748
rect 30558 16736 30564 16748
rect 30616 16736 30622 16788
rect 33318 16776 33324 16788
rect 33279 16748 33324 16776
rect 33318 16736 33324 16748
rect 33376 16736 33382 16788
rect 35618 16736 35624 16788
rect 35676 16776 35682 16788
rect 35713 16779 35771 16785
rect 35713 16776 35725 16779
rect 35676 16748 35725 16776
rect 35676 16736 35682 16748
rect 35713 16745 35725 16748
rect 35759 16745 35771 16779
rect 35713 16739 35771 16745
rect 25593 16711 25651 16717
rect 25593 16677 25605 16711
rect 25639 16708 25651 16711
rect 25682 16708 25688 16720
rect 25639 16680 25688 16708
rect 25639 16677 25651 16680
rect 25593 16671 25651 16677
rect 25682 16668 25688 16680
rect 25740 16708 25746 16720
rect 35161 16711 35219 16717
rect 35161 16708 35173 16711
rect 25740 16680 35173 16708
rect 25740 16668 25746 16680
rect 35161 16677 35173 16680
rect 35207 16677 35219 16711
rect 35161 16671 35219 16677
rect 21573 16581 21601 16668
rect 21726 16600 21732 16652
rect 21784 16600 21790 16652
rect 26050 16600 26056 16652
rect 26108 16640 26114 16652
rect 27246 16640 27252 16652
rect 26108 16612 27252 16640
rect 26108 16600 26114 16612
rect 27246 16600 27252 16612
rect 27304 16600 27310 16652
rect 27338 16600 27344 16652
rect 27396 16640 27402 16652
rect 29917 16643 29975 16649
rect 29917 16640 29929 16643
rect 27396 16612 29929 16640
rect 27396 16600 27402 16612
rect 29917 16609 29929 16612
rect 29963 16640 29975 16643
rect 32122 16640 32128 16652
rect 29963 16612 32128 16640
rect 29963 16609 29975 16612
rect 29917 16603 29975 16609
rect 32122 16600 32128 16612
rect 32180 16600 32186 16652
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 18288 16544 18337 16572
rect 18288 16532 18294 16544
rect 18325 16541 18337 16544
rect 18371 16572 18383 16575
rect 19613 16575 19671 16581
rect 19613 16572 19625 16575
rect 18371 16544 19625 16572
rect 18371 16541 18383 16544
rect 18325 16535 18383 16541
rect 19613 16541 19625 16544
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 21453 16575 21511 16581
rect 21453 16541 21465 16575
rect 21499 16541 21511 16575
rect 21453 16535 21511 16541
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16541 21603 16575
rect 21545 16535 21603 16541
rect 21637 16575 21695 16581
rect 21637 16541 21649 16575
rect 21683 16572 21695 16575
rect 21744 16572 21772 16600
rect 21683 16544 21772 16572
rect 21821 16575 21879 16581
rect 21683 16541 21695 16544
rect 21637 16535 21695 16541
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 26513 16575 26571 16581
rect 26513 16541 26525 16575
rect 26559 16572 26571 16575
rect 26602 16572 26608 16584
rect 26559 16544 26608 16572
rect 26559 16541 26571 16544
rect 26513 16535 26571 16541
rect 14550 16504 14556 16516
rect 10060 16476 14556 16504
rect 14550 16464 14556 16476
rect 14608 16464 14614 16516
rect 18138 16504 18144 16516
rect 18099 16476 18144 16504
rect 18138 16464 18144 16476
rect 18196 16464 18202 16516
rect 19426 16504 19432 16516
rect 19387 16476 19432 16504
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 21836 16504 21864 16535
rect 26602 16532 26608 16544
rect 26660 16532 26666 16584
rect 29822 16532 29828 16584
rect 29880 16572 29886 16584
rect 30193 16575 30251 16581
rect 30193 16572 30205 16575
rect 29880 16544 30205 16572
rect 29880 16532 29886 16544
rect 30193 16541 30205 16544
rect 30239 16541 30251 16575
rect 35176 16572 35204 16671
rect 37826 16640 37832 16652
rect 36832 16612 37832 16640
rect 35618 16572 35624 16584
rect 35176 16544 35624 16572
rect 30193 16535 30251 16541
rect 35618 16532 35624 16544
rect 35676 16572 35682 16584
rect 35989 16575 36047 16581
rect 35989 16572 36001 16575
rect 35676 16544 36001 16572
rect 35676 16532 35682 16544
rect 35989 16541 36001 16544
rect 36035 16541 36047 16575
rect 35989 16535 36047 16541
rect 36081 16575 36139 16581
rect 36081 16541 36093 16575
rect 36127 16541 36139 16575
rect 36081 16535 36139 16541
rect 26326 16504 26332 16516
rect 21836 16476 22416 16504
rect 26239 16476 26332 16504
rect 2222 16436 2228 16448
rect 2183 16408 2228 16436
rect 2222 16396 2228 16408
rect 2280 16396 2286 16448
rect 4801 16439 4859 16445
rect 4801 16405 4813 16439
rect 4847 16436 4859 16439
rect 5718 16436 5724 16448
rect 4847 16408 5724 16436
rect 4847 16405 4859 16408
rect 4801 16399 4859 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 7006 16436 7012 16448
rect 6967 16408 7012 16436
rect 7006 16396 7012 16408
rect 7064 16396 7070 16448
rect 8846 16396 8852 16448
rect 8904 16436 8910 16448
rect 9490 16436 9496 16448
rect 8904 16408 9496 16436
rect 8904 16396 8910 16408
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 10781 16439 10839 16445
rect 10781 16405 10793 16439
rect 10827 16436 10839 16439
rect 11238 16436 11244 16448
rect 10827 16408 11244 16436
rect 10827 16405 10839 16408
rect 10781 16399 10839 16405
rect 11238 16396 11244 16408
rect 11296 16436 11302 16448
rect 11517 16439 11575 16445
rect 11517 16436 11529 16439
rect 11296 16408 11529 16436
rect 11296 16396 11302 16408
rect 11517 16405 11529 16408
rect 11563 16436 11575 16439
rect 12158 16436 12164 16448
rect 11563 16408 12164 16436
rect 11563 16405 11575 16408
rect 11517 16399 11575 16405
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 16850 16436 16856 16448
rect 16811 16408 16856 16436
rect 16850 16396 16856 16408
rect 16908 16396 16914 16448
rect 19334 16396 19340 16448
rect 19392 16436 19398 16448
rect 22388 16445 22416 16476
rect 26326 16464 26332 16476
rect 26384 16504 26390 16516
rect 26694 16504 26700 16516
rect 26384 16476 26700 16504
rect 26384 16464 26390 16476
rect 26694 16464 26700 16476
rect 26752 16464 26758 16516
rect 27154 16464 27160 16516
rect 27212 16504 27218 16516
rect 27249 16507 27307 16513
rect 27249 16504 27261 16507
rect 27212 16476 27261 16504
rect 27212 16464 27218 16476
rect 27249 16473 27261 16476
rect 27295 16504 27307 16507
rect 30558 16504 30564 16516
rect 27295 16476 30564 16504
rect 27295 16473 27307 16476
rect 27249 16467 27307 16473
rect 30558 16464 30564 16476
rect 30616 16464 30622 16516
rect 36096 16504 36124 16535
rect 36170 16532 36176 16584
rect 36228 16572 36234 16584
rect 36228 16544 36273 16572
rect 36228 16532 36234 16544
rect 36354 16532 36360 16584
rect 36412 16572 36418 16584
rect 36412 16544 36457 16572
rect 36412 16532 36418 16544
rect 36832 16504 36860 16612
rect 37826 16600 37832 16612
rect 37884 16600 37890 16652
rect 36998 16572 37004 16584
rect 36959 16544 37004 16572
rect 36998 16532 37004 16544
rect 37056 16532 37062 16584
rect 37366 16572 37372 16584
rect 37327 16544 37372 16572
rect 37366 16532 37372 16544
rect 37424 16532 37430 16584
rect 38930 16532 38936 16584
rect 38988 16572 38994 16584
rect 39853 16575 39911 16581
rect 39853 16572 39865 16575
rect 38988 16544 39865 16572
rect 38988 16532 38994 16544
rect 39853 16541 39865 16544
rect 39899 16541 39911 16575
rect 39853 16535 39911 16541
rect 36096 16476 36860 16504
rect 37093 16507 37151 16513
rect 37093 16473 37105 16507
rect 37139 16473 37151 16507
rect 37093 16467 37151 16473
rect 37185 16507 37243 16513
rect 37185 16473 37197 16507
rect 37231 16504 37243 16507
rect 37642 16504 37648 16516
rect 37231 16476 37648 16504
rect 37231 16473 37243 16476
rect 37185 16467 37243 16473
rect 20073 16439 20131 16445
rect 20073 16436 20085 16439
rect 19392 16408 20085 16436
rect 19392 16396 19398 16408
rect 20073 16405 20085 16408
rect 20119 16405 20131 16439
rect 20073 16399 20131 16405
rect 22373 16439 22431 16445
rect 22373 16405 22385 16439
rect 22419 16436 22431 16439
rect 22462 16436 22468 16448
rect 22419 16408 22468 16436
rect 22419 16405 22431 16408
rect 22373 16399 22431 16405
rect 22462 16396 22468 16408
rect 22520 16396 22526 16448
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 22833 16439 22891 16445
rect 22833 16436 22845 16439
rect 22704 16408 22845 16436
rect 22704 16396 22710 16408
rect 22833 16405 22845 16408
rect 22879 16405 22891 16439
rect 22833 16399 22891 16405
rect 28813 16439 28871 16445
rect 28813 16405 28825 16439
rect 28859 16436 28871 16439
rect 29178 16436 29184 16448
rect 28859 16408 29184 16436
rect 28859 16405 28871 16408
rect 28813 16399 28871 16405
rect 29178 16396 29184 16408
rect 29236 16396 29242 16448
rect 30374 16396 30380 16448
rect 30432 16436 30438 16448
rect 36817 16439 36875 16445
rect 36817 16436 36829 16439
rect 30432 16408 36829 16436
rect 30432 16396 30438 16408
rect 36817 16405 36829 16408
rect 36863 16405 36875 16439
rect 37108 16436 37136 16467
rect 37642 16464 37648 16476
rect 37700 16464 37706 16516
rect 40034 16504 40040 16516
rect 39995 16476 40040 16504
rect 40034 16464 40040 16476
rect 40092 16464 40098 16516
rect 37366 16436 37372 16448
rect 37108 16408 37372 16436
rect 36817 16399 36875 16405
rect 37366 16396 37372 16408
rect 37424 16396 37430 16448
rect 40218 16436 40224 16448
rect 40179 16408 40224 16436
rect 40218 16396 40224 16408
rect 40276 16396 40282 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 3329 16235 3387 16241
rect 3329 16201 3341 16235
rect 3375 16232 3387 16235
rect 4249 16235 4307 16241
rect 4249 16232 4261 16235
rect 3375 16204 4261 16232
rect 3375 16201 3387 16204
rect 3329 16195 3387 16201
rect 4249 16201 4261 16204
rect 4295 16201 4307 16235
rect 4249 16195 4307 16201
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 7834 16232 7840 16244
rect 5675 16204 7840 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 2222 16173 2228 16176
rect 2216 16164 2228 16173
rect 2183 16136 2228 16164
rect 2216 16127 2228 16136
rect 2222 16124 2228 16127
rect 2280 16124 2286 16176
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4264 16096 4292 16195
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 10686 16232 10692 16244
rect 9815 16204 10692 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 11885 16235 11943 16241
rect 11885 16201 11897 16235
rect 11931 16232 11943 16235
rect 11974 16232 11980 16244
rect 11931 16204 11980 16232
rect 11931 16201 11943 16204
rect 11885 16195 11943 16201
rect 11974 16192 11980 16204
rect 12032 16192 12038 16244
rect 17402 16232 17408 16244
rect 17363 16204 17408 16232
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 20806 16232 20812 16244
rect 19996 16204 20812 16232
rect 4985 16167 5043 16173
rect 4985 16133 4997 16167
rect 5031 16164 5043 16167
rect 5718 16164 5724 16176
rect 5031 16136 5724 16164
rect 5031 16133 5043 16136
rect 4985 16127 5043 16133
rect 5718 16124 5724 16136
rect 5776 16124 5782 16176
rect 9490 16124 9496 16176
rect 9548 16164 9554 16176
rect 10597 16167 10655 16173
rect 9548 16136 9904 16164
rect 9548 16124 9554 16136
rect 5353 16099 5411 16105
rect 5353 16096 5365 16099
rect 4264 16068 5365 16096
rect 4157 16059 4215 16065
rect 5353 16065 5365 16068
rect 5399 16065 5411 16099
rect 5353 16059 5411 16065
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 7285 16099 7343 16105
rect 7285 16065 7297 16099
rect 7331 16096 7343 16099
rect 8110 16096 8116 16108
rect 7331 16068 8116 16096
rect 7331 16065 7343 16068
rect 7285 16059 7343 16065
rect 1946 16028 1952 16040
rect 1907 16000 1952 16028
rect 1946 15988 1952 16000
rect 2004 15988 2010 16040
rect 4172 16028 4200 16059
rect 4433 16031 4491 16037
rect 4172 16000 4292 16028
rect 3786 15892 3792 15904
rect 3747 15864 3792 15892
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 4264 15892 4292 16000
rect 4433 15997 4445 16031
rect 4479 15997 4491 16031
rect 4433 15991 4491 15997
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 16028 5503 16031
rect 5534 16028 5540 16040
rect 5491 16000 5540 16028
rect 5491 15997 5503 16000
rect 5445 15991 5503 15997
rect 4448 15960 4476 15991
rect 5534 15988 5540 16000
rect 5592 16028 5598 16040
rect 6822 16028 6828 16040
rect 5592 16000 6828 16028
rect 5592 15988 5598 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 4798 15960 4804 15972
rect 4448 15932 4804 15960
rect 4798 15920 4804 15932
rect 4856 15960 4862 15972
rect 5350 15960 5356 15972
rect 4856 15932 5356 15960
rect 4856 15920 4862 15932
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 7116 15960 7144 16059
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 9125 16099 9183 16105
rect 9125 16065 9137 16099
rect 9171 16096 9183 16099
rect 9674 16096 9680 16108
rect 9171 16068 9680 16096
rect 9171 16065 9183 16068
rect 9125 16059 9183 16065
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 9876 16105 9904 16136
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 12342 16164 12348 16176
rect 10643 16136 12348 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 12342 16124 12348 16136
rect 12400 16124 12406 16176
rect 12526 16124 12532 16176
rect 12584 16164 12590 16176
rect 12584 16136 18359 16164
rect 12584 16124 12590 16136
rect 10502 16105 10508 16108
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16065 9919 16099
rect 10500 16096 10508 16105
rect 10463 16068 10508 16096
rect 9861 16059 9919 16065
rect 10500 16059 10508 16068
rect 10502 16056 10508 16059
rect 10560 16056 10566 16108
rect 10686 16096 10692 16108
rect 10647 16068 10692 16096
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 10778 16056 10784 16108
rect 10836 16105 10842 16108
rect 10836 16099 10875 16105
rect 10863 16065 10875 16099
rect 10836 16059 10875 16065
rect 10836 16056 10842 16059
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 11793 16099 11851 16105
rect 11020 16068 11065 16096
rect 11020 16056 11026 16068
rect 11793 16065 11805 16099
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12158 16096 12164 16108
rect 12023 16068 12164 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 11808 16028 11836 16059
rect 12158 16056 12164 16068
rect 12216 16096 12222 16108
rect 14182 16096 14188 16108
rect 12216 16068 14188 16096
rect 12216 16056 12222 16068
rect 14182 16056 14188 16068
rect 14240 16056 14246 16108
rect 14458 16096 14464 16108
rect 14371 16068 14464 16096
rect 14458 16056 14464 16068
rect 14516 16096 14522 16108
rect 15010 16096 15016 16108
rect 14516 16068 15016 16096
rect 14516 16056 14522 16068
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 17589 16099 17647 16105
rect 17589 16065 17601 16099
rect 17635 16065 17647 16099
rect 17589 16059 17647 16065
rect 17773 16099 17831 16105
rect 17773 16065 17785 16099
rect 17819 16096 17831 16099
rect 18046 16096 18052 16108
rect 17819 16068 18052 16096
rect 17819 16065 17831 16068
rect 17773 16059 17831 16065
rect 12526 16028 12532 16040
rect 10612 16000 12532 16028
rect 10321 15963 10379 15969
rect 10321 15960 10333 15963
rect 7116 15932 10333 15960
rect 10321 15929 10333 15932
rect 10367 15929 10379 15963
rect 10321 15923 10379 15929
rect 4614 15892 4620 15904
rect 4264 15864 4620 15892
rect 4614 15852 4620 15864
rect 4672 15892 4678 15904
rect 6914 15892 6920 15904
rect 4672 15864 6920 15892
rect 4672 15852 4678 15864
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7466 15892 7472 15904
rect 7427 15864 7472 15892
rect 7466 15852 7472 15864
rect 7524 15852 7530 15904
rect 8021 15895 8079 15901
rect 8021 15861 8033 15895
rect 8067 15892 8079 15895
rect 8110 15892 8116 15904
rect 8067 15864 8116 15892
rect 8067 15861 8079 15864
rect 8021 15855 8079 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 8665 15895 8723 15901
rect 8665 15861 8677 15895
rect 8711 15892 8723 15895
rect 8846 15892 8852 15904
rect 8711 15864 8852 15892
rect 8711 15861 8723 15864
rect 8665 15855 8723 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 9214 15852 9220 15904
rect 9272 15892 9278 15904
rect 10612 15892 10640 16000
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 14737 16031 14795 16037
rect 14737 15997 14749 16031
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 14274 15920 14280 15972
rect 14332 15960 14338 15972
rect 14752 15960 14780 15991
rect 14332 15932 14780 15960
rect 17604 15960 17632 16059
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 18233 16099 18291 16105
rect 18233 16065 18245 16099
rect 18279 16065 18291 16099
rect 18331 16096 18359 16136
rect 19242 16124 19248 16176
rect 19300 16164 19306 16176
rect 19996 16173 20024 16204
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 28994 16232 29000 16244
rect 28368 16204 29000 16232
rect 19981 16167 20039 16173
rect 19981 16164 19993 16167
rect 19300 16136 19993 16164
rect 19300 16124 19306 16136
rect 19981 16133 19993 16136
rect 20027 16133 20039 16167
rect 19981 16127 20039 16133
rect 20717 16167 20775 16173
rect 20717 16133 20729 16167
rect 20763 16164 20775 16167
rect 26878 16164 26884 16176
rect 20763 16136 26884 16164
rect 20763 16133 20775 16136
rect 20717 16127 20775 16133
rect 26878 16124 26884 16136
rect 26936 16124 26942 16176
rect 28258 16164 28264 16176
rect 28219 16136 28264 16164
rect 28258 16124 28264 16136
rect 28316 16124 28322 16176
rect 19334 16096 19340 16108
rect 18331 16068 19340 16096
rect 18233 16059 18291 16065
rect 17954 15960 17960 15972
rect 17604 15932 17960 15960
rect 14332 15920 14338 15932
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 9272 15864 10640 15892
rect 16945 15895 17003 15901
rect 9272 15852 9278 15864
rect 16945 15861 16957 15895
rect 16991 15892 17003 15895
rect 17034 15892 17040 15904
rect 16991 15864 17040 15892
rect 16991 15861 17003 15864
rect 16945 15855 17003 15861
rect 17034 15852 17040 15864
rect 17092 15892 17098 15904
rect 18248 15892 18276 16059
rect 19334 16056 19340 16068
rect 19392 16096 19398 16108
rect 20530 16096 20536 16108
rect 19392 16068 20536 16096
rect 19392 16056 19398 16068
rect 20530 16056 20536 16068
rect 20588 16096 20594 16108
rect 20625 16099 20683 16105
rect 20625 16096 20637 16099
rect 20588 16068 20637 16096
rect 20588 16056 20594 16068
rect 20625 16065 20637 16068
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 20809 16099 20867 16105
rect 20809 16065 20821 16099
rect 20855 16096 20867 16099
rect 20990 16096 20996 16108
rect 20855 16068 20996 16096
rect 20855 16065 20867 16068
rect 20809 16059 20867 16065
rect 20990 16056 20996 16068
rect 21048 16096 21054 16108
rect 21266 16096 21272 16108
rect 21048 16068 21272 16096
rect 21048 16056 21054 16068
rect 21266 16056 21272 16068
rect 21324 16096 21330 16108
rect 21634 16096 21640 16108
rect 21324 16068 21640 16096
rect 21324 16056 21330 16068
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 22738 16096 22744 16108
rect 22699 16068 22744 16096
rect 22738 16056 22744 16068
rect 22796 16056 22802 16108
rect 22922 16056 22928 16108
rect 22980 16096 22986 16108
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 22980 16068 23029 16096
rect 22980 16056 22986 16068
rect 23017 16065 23029 16068
rect 23063 16065 23075 16099
rect 23474 16096 23480 16108
rect 23387 16068 23480 16096
rect 23017 16059 23075 16065
rect 23474 16056 23480 16068
rect 23532 16096 23538 16108
rect 24026 16096 24032 16108
rect 23532 16068 24032 16096
rect 23532 16056 23538 16068
rect 24026 16056 24032 16068
rect 24084 16056 24090 16108
rect 26418 16056 26424 16108
rect 26476 16096 26482 16108
rect 27157 16099 27215 16105
rect 27157 16096 27169 16099
rect 26476 16068 27169 16096
rect 26476 16056 26482 16068
rect 27157 16065 27169 16068
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 28077 16099 28135 16105
rect 28077 16065 28089 16099
rect 28123 16096 28135 16099
rect 28166 16096 28172 16108
rect 28123 16068 28172 16096
rect 28123 16065 28135 16068
rect 28077 16059 28135 16065
rect 28166 16056 28172 16068
rect 28224 16096 28230 16108
rect 28368 16096 28396 16204
rect 28994 16192 29000 16204
rect 29052 16192 29058 16244
rect 29914 16192 29920 16244
rect 29972 16232 29978 16244
rect 30009 16235 30067 16241
rect 30009 16232 30021 16235
rect 29972 16204 30021 16232
rect 29972 16192 29978 16204
rect 30009 16201 30021 16204
rect 30055 16201 30067 16235
rect 30009 16195 30067 16201
rect 32953 16235 33011 16241
rect 32953 16201 32965 16235
rect 32999 16232 33011 16235
rect 33686 16232 33692 16244
rect 32999 16204 33692 16232
rect 32999 16201 33011 16204
rect 32953 16195 33011 16201
rect 33686 16192 33692 16204
rect 33744 16192 33750 16244
rect 38289 16235 38347 16241
rect 38289 16232 38301 16235
rect 33980 16204 38301 16232
rect 28445 16167 28503 16173
rect 28445 16133 28457 16167
rect 28491 16164 28503 16167
rect 28491 16136 29132 16164
rect 28491 16133 28503 16136
rect 28445 16127 28503 16133
rect 29104 16105 29132 16136
rect 29196 16136 29960 16164
rect 29196 16105 29224 16136
rect 29932 16108 29960 16136
rect 30558 16124 30564 16176
rect 30616 16164 30622 16176
rect 33980 16164 34008 16204
rect 38289 16201 38301 16204
rect 38335 16232 38347 16235
rect 38562 16232 38568 16244
rect 38335 16204 38568 16232
rect 38335 16201 38347 16204
rect 38289 16195 38347 16201
rect 38562 16192 38568 16204
rect 38620 16192 38626 16244
rect 40221 16235 40279 16241
rect 40221 16201 40233 16235
rect 40267 16201 40279 16235
rect 40221 16195 40279 16201
rect 30616 16136 34008 16164
rect 30616 16124 30622 16136
rect 34054 16124 34060 16176
rect 34112 16173 34118 16176
rect 34112 16164 34124 16173
rect 37553 16167 37611 16173
rect 34112 16136 34157 16164
rect 34112 16127 34124 16136
rect 37553 16133 37565 16167
rect 37599 16164 37611 16167
rect 40034 16164 40040 16176
rect 37599 16136 40040 16164
rect 37599 16133 37611 16136
rect 37553 16127 37611 16133
rect 34112 16124 34118 16127
rect 40034 16124 40040 16136
rect 40092 16164 40098 16176
rect 40236 16164 40264 16195
rect 40092 16136 40264 16164
rect 40092 16124 40098 16136
rect 28224 16068 28396 16096
rect 28905 16099 28963 16105
rect 28224 16056 28230 16068
rect 28905 16065 28917 16099
rect 28951 16065 28963 16099
rect 28905 16059 28963 16065
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16065 29147 16099
rect 29089 16059 29147 16065
rect 29181 16099 29239 16105
rect 29181 16065 29193 16099
rect 29227 16065 29239 16099
rect 29181 16059 29239 16065
rect 23290 15988 23296 16040
rect 23348 16028 23354 16040
rect 23753 16031 23811 16037
rect 23753 16028 23765 16031
rect 23348 16000 23765 16028
rect 23348 15988 23354 16000
rect 23753 15997 23765 16000
rect 23799 16028 23811 16031
rect 26436 16028 26464 16056
rect 27341 16031 27399 16037
rect 27341 16028 27353 16031
rect 23799 16000 26464 16028
rect 26620 16000 27353 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 17092 15864 18276 15892
rect 17092 15852 17098 15864
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 22646 15892 22652 15904
rect 19944 15864 22652 15892
rect 19944 15852 19950 15864
rect 22646 15852 22652 15864
rect 22704 15852 22710 15904
rect 26326 15892 26332 15904
rect 26287 15864 26332 15892
rect 26326 15852 26332 15864
rect 26384 15892 26390 15904
rect 26620 15892 26648 16000
rect 27341 15997 27353 16000
rect 27387 16028 27399 16031
rect 27430 16028 27436 16040
rect 27387 16000 27436 16028
rect 27387 15997 27399 16000
rect 27341 15991 27399 15997
rect 27430 15988 27436 16000
rect 27488 15988 27494 16040
rect 28920 16028 28948 16059
rect 29270 16056 29276 16108
rect 29328 16096 29334 16108
rect 29328 16068 29373 16096
rect 29328 16056 29334 16068
rect 29914 16056 29920 16108
rect 29972 16056 29978 16108
rect 30374 16056 30380 16108
rect 30432 16096 30438 16108
rect 31122 16099 31180 16105
rect 31122 16096 31134 16099
rect 30432 16068 31134 16096
rect 30432 16056 30438 16068
rect 31122 16065 31134 16068
rect 31168 16065 31180 16099
rect 31122 16059 31180 16065
rect 35805 16099 35863 16105
rect 35805 16065 35817 16099
rect 35851 16096 35863 16099
rect 36998 16096 37004 16108
rect 35851 16068 37004 16096
rect 35851 16065 35863 16068
rect 35805 16059 35863 16065
rect 36998 16056 37004 16068
rect 37056 16096 37062 16108
rect 37274 16096 37280 16108
rect 37056 16068 37280 16096
rect 37056 16056 37062 16068
rect 37274 16056 37280 16068
rect 37332 16096 37338 16108
rect 37461 16099 37519 16105
rect 37461 16096 37473 16099
rect 37332 16068 37473 16096
rect 37332 16056 37338 16068
rect 37461 16065 37473 16068
rect 37507 16065 37519 16099
rect 37642 16096 37648 16108
rect 37603 16068 37648 16096
rect 37461 16059 37519 16065
rect 37642 16056 37648 16068
rect 37700 16056 37706 16108
rect 37829 16099 37887 16105
rect 37829 16065 37841 16099
rect 37875 16096 37887 16099
rect 38654 16096 38660 16108
rect 37875 16068 38660 16096
rect 37875 16065 37887 16068
rect 37829 16059 37887 16065
rect 38654 16056 38660 16068
rect 38712 16056 38718 16108
rect 38746 16056 38752 16108
rect 38804 16096 38810 16108
rect 38841 16099 38899 16105
rect 38841 16096 38853 16099
rect 38804 16068 38853 16096
rect 38804 16056 38810 16068
rect 38841 16065 38853 16068
rect 38887 16065 38899 16099
rect 38841 16059 38899 16065
rect 39108 16099 39166 16105
rect 39108 16065 39120 16099
rect 39154 16096 39166 16099
rect 39850 16096 39856 16108
rect 39154 16068 39856 16096
rect 39154 16065 39166 16068
rect 39108 16059 39166 16065
rect 39850 16056 39856 16068
rect 39908 16056 39914 16108
rect 29454 16028 29460 16040
rect 28920 16000 29460 16028
rect 29454 15988 29460 16000
rect 29512 15988 29518 16040
rect 31389 16031 31447 16037
rect 31389 15997 31401 16031
rect 31435 16028 31447 16031
rect 31754 16028 31760 16040
rect 31435 16000 31760 16028
rect 31435 15997 31447 16000
rect 31389 15991 31447 15997
rect 31754 15988 31760 16000
rect 31812 15988 31818 16040
rect 34333 16031 34391 16037
rect 34333 15997 34345 16031
rect 34379 16028 34391 16031
rect 34514 16028 34520 16040
rect 34379 16000 34520 16028
rect 34379 15997 34391 16000
rect 34333 15991 34391 15997
rect 34514 15988 34520 16000
rect 34572 15988 34578 16040
rect 35526 16028 35532 16040
rect 35487 16000 35532 16028
rect 35526 15988 35532 16000
rect 35584 15988 35590 16040
rect 40678 16028 40684 16040
rect 40639 16000 40684 16028
rect 40678 15988 40684 16000
rect 40736 15988 40742 16040
rect 40954 16028 40960 16040
rect 40915 16000 40960 16028
rect 40954 15988 40960 16000
rect 41012 15988 41018 16040
rect 26694 15920 26700 15972
rect 26752 15960 26758 15972
rect 26973 15963 27031 15969
rect 26973 15960 26985 15963
rect 26752 15932 26985 15960
rect 26752 15920 26758 15932
rect 26973 15929 26985 15932
rect 27019 15960 27031 15963
rect 28810 15960 28816 15972
rect 27019 15932 28816 15960
rect 27019 15929 27031 15932
rect 26973 15923 27031 15929
rect 28810 15920 28816 15932
rect 28868 15920 28874 15972
rect 37274 15960 37280 15972
rect 37235 15932 37280 15960
rect 37274 15920 37280 15932
rect 37332 15920 37338 15972
rect 29546 15892 29552 15904
rect 26384 15864 26648 15892
rect 29507 15864 29552 15892
rect 26384 15852 26390 15864
rect 29546 15852 29552 15864
rect 29604 15852 29610 15904
rect 58158 15892 58164 15904
rect 58119 15864 58164 15892
rect 58158 15852 58164 15864
rect 58216 15852 58222 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 9953 15691 10011 15697
rect 9953 15688 9965 15691
rect 9824 15660 9965 15688
rect 9824 15648 9830 15660
rect 9953 15657 9965 15660
rect 9999 15657 10011 15691
rect 13170 15688 13176 15700
rect 9953 15651 10011 15657
rect 11716 15660 13176 15688
rect 10594 15580 10600 15632
rect 10652 15620 10658 15632
rect 10652 15592 11192 15620
rect 10652 15580 10658 15592
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 2774 15552 2780 15564
rect 2179 15524 2780 15552
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 2774 15512 2780 15524
rect 2832 15512 2838 15564
rect 10042 15552 10048 15564
rect 10003 15524 10048 15552
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 10686 15512 10692 15564
rect 10744 15552 10750 15564
rect 11164 15552 11192 15592
rect 11716 15561 11744 15660
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 14458 15688 14464 15700
rect 14419 15660 14464 15688
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 14550 15648 14556 15700
rect 14608 15688 14614 15700
rect 14608 15660 17356 15688
rect 14608 15648 14614 15660
rect 13078 15620 13084 15632
rect 13039 15592 13084 15620
rect 13078 15580 13084 15592
rect 13136 15580 13142 15632
rect 14182 15580 14188 15632
rect 14240 15620 14246 15632
rect 17221 15623 17279 15629
rect 17221 15620 17233 15623
rect 14240 15592 17233 15620
rect 14240 15580 14246 15592
rect 17221 15589 17233 15592
rect 17267 15589 17279 15623
rect 17328 15620 17356 15660
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 18472 15660 18521 15688
rect 18472 15648 18478 15660
rect 18509 15657 18521 15660
rect 18555 15657 18567 15691
rect 19334 15688 19340 15700
rect 19295 15660 19340 15688
rect 18509 15651 18567 15657
rect 19334 15648 19340 15660
rect 19392 15648 19398 15700
rect 19886 15688 19892 15700
rect 19847 15660 19892 15688
rect 19886 15648 19892 15660
rect 19944 15648 19950 15700
rect 20346 15688 20352 15700
rect 20307 15660 20352 15688
rect 20346 15648 20352 15660
rect 20404 15648 20410 15700
rect 22741 15691 22799 15697
rect 22741 15657 22753 15691
rect 22787 15688 22799 15691
rect 22922 15688 22928 15700
rect 22787 15660 22928 15688
rect 22787 15657 22799 15660
rect 22741 15651 22799 15657
rect 22922 15648 22928 15660
rect 22980 15648 22986 15700
rect 23385 15691 23443 15697
rect 23385 15657 23397 15691
rect 23431 15688 23443 15691
rect 23474 15688 23480 15700
rect 23431 15660 23480 15688
rect 23431 15657 23443 15660
rect 23385 15651 23443 15657
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 26234 15648 26240 15700
rect 26292 15688 26298 15700
rect 26329 15691 26387 15697
rect 26329 15688 26341 15691
rect 26292 15660 26341 15688
rect 26292 15648 26298 15660
rect 26329 15657 26341 15660
rect 26375 15657 26387 15691
rect 26329 15651 26387 15657
rect 28258 15648 28264 15700
rect 28316 15688 28322 15700
rect 29549 15691 29607 15697
rect 29549 15688 29561 15691
rect 28316 15660 29561 15688
rect 28316 15648 28322 15660
rect 29549 15657 29561 15660
rect 29595 15657 29607 15691
rect 29549 15651 29607 15657
rect 36170 15648 36176 15700
rect 36228 15688 36234 15700
rect 36725 15691 36783 15697
rect 36725 15688 36737 15691
rect 36228 15660 36737 15688
rect 36228 15648 36234 15660
rect 36725 15657 36737 15660
rect 36771 15688 36783 15691
rect 37458 15688 37464 15700
rect 36771 15660 37464 15688
rect 36771 15657 36783 15660
rect 36725 15651 36783 15657
rect 37458 15648 37464 15660
rect 37516 15648 37522 15700
rect 39850 15688 39856 15700
rect 39811 15660 39856 15688
rect 39850 15648 39856 15660
rect 39908 15648 39914 15700
rect 22002 15620 22008 15632
rect 17328 15592 22008 15620
rect 17221 15583 17279 15589
rect 11701 15555 11759 15561
rect 10744 15524 11008 15552
rect 11164 15524 11284 15552
rect 10744 15512 10750 15524
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 3786 15484 3792 15496
rect 2363 15456 3792 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 8294 15484 8300 15496
rect 8255 15456 8300 15484
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 10778 15493 10784 15496
rect 10137 15487 10195 15493
rect 10137 15453 10149 15487
rect 10183 15484 10195 15487
rect 10776 15484 10784 15493
rect 10183 15456 10640 15484
rect 10739 15456 10784 15484
rect 10183 15453 10195 15456
rect 10137 15447 10195 15453
rect 7282 15376 7288 15428
rect 7340 15416 7346 15428
rect 8030 15419 8088 15425
rect 8030 15416 8042 15419
rect 7340 15388 8042 15416
rect 7340 15376 7346 15388
rect 8030 15385 8042 15388
rect 8076 15385 8088 15419
rect 8030 15379 8088 15385
rect 4614 15308 4620 15360
rect 4672 15348 4678 15360
rect 4709 15351 4767 15357
rect 4709 15348 4721 15351
rect 4672 15320 4721 15348
rect 4672 15308 4678 15320
rect 4709 15317 4721 15320
rect 4755 15348 4767 15351
rect 4798 15348 4804 15360
rect 4755 15320 4804 15348
rect 4755 15317 4767 15320
rect 4709 15311 4767 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 6914 15348 6920 15360
rect 6875 15320 6920 15348
rect 6914 15308 6920 15320
rect 6972 15308 6978 15360
rect 8478 15308 8484 15360
rect 8536 15348 8542 15360
rect 10612 15357 10640 15456
rect 10776 15447 10784 15456
rect 10778 15444 10784 15447
rect 10836 15444 10842 15496
rect 10980 15425 11008 15524
rect 11146 15484 11152 15496
rect 11107 15456 11152 15484
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11256 15493 11284 15524
rect 11701 15521 11713 15555
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 11790 15444 11796 15496
rect 11848 15484 11854 15496
rect 11957 15487 12015 15493
rect 11957 15484 11969 15487
rect 11848 15456 11969 15484
rect 11848 15444 11854 15456
rect 11957 15453 11969 15456
rect 12003 15453 12015 15487
rect 11957 15447 12015 15453
rect 13170 15444 13176 15496
rect 13228 15484 13234 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 13228 15456 14289 15484
rect 13228 15444 13234 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 14550 15484 14556 15496
rect 14507 15456 14556 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 10873 15419 10931 15425
rect 10873 15385 10885 15419
rect 10919 15385 10931 15419
rect 10873 15379 10931 15385
rect 10965 15419 11023 15425
rect 10965 15385 10977 15419
rect 11011 15416 11023 15419
rect 12618 15416 12624 15428
rect 11011 15388 12624 15416
rect 11011 15385 11023 15388
rect 10965 15379 11023 15385
rect 9769 15351 9827 15357
rect 9769 15348 9781 15351
rect 8536 15320 9781 15348
rect 8536 15308 8542 15320
rect 9769 15317 9781 15320
rect 9815 15317 9827 15351
rect 9769 15311 9827 15317
rect 10597 15351 10655 15357
rect 10597 15317 10609 15351
rect 10643 15317 10655 15351
rect 10888 15348 10916 15379
rect 12618 15376 12624 15388
rect 12676 15416 12682 15428
rect 14182 15416 14188 15428
rect 12676 15388 14188 15416
rect 12676 15376 12682 15388
rect 14182 15376 14188 15388
rect 14240 15376 14246 15428
rect 14292 15416 14320 15447
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 17236 15484 17264 15583
rect 22002 15580 22008 15592
rect 22060 15580 22066 15632
rect 22097 15623 22155 15629
rect 22097 15589 22109 15623
rect 22143 15620 22155 15623
rect 28994 15620 29000 15632
rect 22143 15592 27384 15620
rect 28955 15592 29000 15620
rect 22143 15589 22155 15592
rect 22097 15583 22155 15589
rect 22646 15552 22652 15564
rect 18340 15524 19334 15552
rect 18340 15493 18368 15524
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 17236 15456 18337 15484
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 18414 15444 18420 15496
rect 18472 15484 18478 15496
rect 18509 15487 18567 15493
rect 18509 15484 18521 15487
rect 18472 15456 18521 15484
rect 18472 15444 18478 15456
rect 18509 15453 18521 15456
rect 18555 15453 18567 15487
rect 19306 15484 19334 15524
rect 22112 15524 22652 15552
rect 19306 15474 20116 15484
rect 19306 15456 20300 15474
rect 18509 15447 18567 15453
rect 20088 15446 20300 15456
rect 14921 15419 14979 15425
rect 14921 15416 14933 15419
rect 14292 15388 14933 15416
rect 14921 15385 14933 15388
rect 14967 15416 14979 15419
rect 16022 15416 16028 15428
rect 14967 15388 16028 15416
rect 14967 15385 14979 15388
rect 14921 15379 14979 15385
rect 16022 15376 16028 15388
rect 16080 15376 16086 15428
rect 19886 15416 19892 15428
rect 16316 15388 19892 15416
rect 16316 15360 16344 15388
rect 19886 15376 19892 15388
rect 19944 15376 19950 15428
rect 20272 15416 20300 15446
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 20530 15484 20536 15496
rect 20404 15456 20449 15484
rect 20491 15456 20536 15484
rect 20404 15444 20410 15456
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 22112 15493 22140 15524
rect 22646 15512 22652 15524
rect 22704 15552 22710 15564
rect 22704 15524 23428 15552
rect 22704 15512 22710 15524
rect 21913 15487 21971 15493
rect 21913 15453 21925 15487
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 22097 15487 22155 15493
rect 22097 15453 22109 15487
rect 22143 15453 22155 15487
rect 22097 15447 22155 15453
rect 21450 15416 21456 15428
rect 20272 15388 21456 15416
rect 21450 15376 21456 15388
rect 21508 15416 21514 15428
rect 21928 15416 21956 15447
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 23400 15493 23428 15524
rect 22557 15487 22615 15493
rect 22557 15484 22569 15487
rect 22244 15456 22569 15484
rect 22244 15444 22250 15456
rect 22557 15453 22569 15456
rect 22603 15453 22615 15487
rect 22557 15447 22615 15453
rect 22741 15487 22799 15493
rect 22741 15453 22753 15487
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 23201 15487 23259 15493
rect 23201 15453 23213 15487
rect 23247 15453 23259 15487
rect 23201 15447 23259 15453
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15484 23443 15487
rect 24302 15484 24308 15496
rect 23431 15456 24308 15484
rect 23431 15453 23443 15456
rect 23385 15447 23443 15453
rect 21508 15388 21956 15416
rect 21508 15376 21514 15388
rect 22002 15376 22008 15428
rect 22060 15416 22066 15428
rect 22370 15416 22376 15428
rect 22060 15388 22376 15416
rect 22060 15376 22066 15388
rect 22370 15376 22376 15388
rect 22428 15416 22434 15428
rect 22756 15416 22784 15447
rect 22428 15388 22784 15416
rect 23216 15416 23244 15447
rect 24302 15444 24308 15456
rect 24360 15444 24366 15496
rect 25777 15487 25835 15493
rect 25777 15453 25789 15487
rect 25823 15484 25835 15487
rect 26234 15484 26240 15496
rect 25823 15456 26240 15484
rect 25823 15453 25835 15456
rect 25777 15447 25835 15453
rect 26234 15444 26240 15456
rect 26292 15444 26298 15496
rect 26418 15484 26424 15496
rect 26379 15456 26424 15484
rect 26418 15444 26424 15456
rect 26476 15444 26482 15496
rect 24397 15419 24455 15425
rect 24397 15416 24409 15419
rect 23216 15388 24409 15416
rect 22428 15376 22434 15388
rect 14090 15348 14096 15360
rect 10888 15320 14096 15348
rect 10597 15311 10655 15317
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 16298 15348 16304 15360
rect 16259 15320 16304 15348
rect 16298 15308 16304 15320
rect 16356 15308 16362 15360
rect 16666 15308 16672 15360
rect 16724 15348 16730 15360
rect 17770 15348 17776 15360
rect 16724 15320 17776 15348
rect 16724 15308 16730 15320
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 20346 15348 20352 15360
rect 19392 15320 20352 15348
rect 19392 15308 19398 15320
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 21358 15348 21364 15360
rect 21319 15320 21364 15348
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 21634 15308 21640 15360
rect 21692 15348 21698 15360
rect 23216 15348 23244 15388
rect 24397 15385 24409 15388
rect 24443 15385 24455 15419
rect 24397 15379 24455 15385
rect 26602 15376 26608 15428
rect 26660 15416 26666 15428
rect 27065 15419 27123 15425
rect 27065 15416 27077 15419
rect 26660 15388 27077 15416
rect 26660 15376 26666 15388
rect 27065 15385 27077 15388
rect 27111 15385 27123 15419
rect 27246 15416 27252 15428
rect 27207 15388 27252 15416
rect 27065 15379 27123 15385
rect 27246 15376 27252 15388
rect 27304 15376 27310 15428
rect 27356 15416 27384 15592
rect 28994 15580 29000 15592
rect 29052 15580 29058 15632
rect 37826 15580 37832 15632
rect 37884 15620 37890 15632
rect 37884 15592 38516 15620
rect 37884 15580 37890 15592
rect 35621 15555 35679 15561
rect 35621 15521 35633 15555
rect 35667 15552 35679 15555
rect 37642 15552 37648 15564
rect 35667 15524 37648 15552
rect 35667 15521 35679 15524
rect 35621 15515 35679 15521
rect 37642 15512 37648 15524
rect 37700 15512 37706 15564
rect 37737 15555 37795 15561
rect 37737 15521 37749 15555
rect 37783 15552 37795 15555
rect 37783 15524 38424 15552
rect 37783 15521 37795 15524
rect 37737 15515 37795 15521
rect 28810 15484 28816 15496
rect 28771 15456 28816 15484
rect 28810 15444 28816 15456
rect 28868 15444 28874 15496
rect 29546 15444 29552 15496
rect 29604 15484 29610 15496
rect 30662 15487 30720 15493
rect 30662 15484 30674 15487
rect 29604 15456 30674 15484
rect 29604 15444 29610 15456
rect 30662 15453 30674 15456
rect 30708 15453 30720 15487
rect 30662 15447 30720 15453
rect 30929 15487 30987 15493
rect 30929 15453 30941 15487
rect 30975 15484 30987 15487
rect 31754 15484 31760 15496
rect 30975 15456 31760 15484
rect 30975 15453 30987 15456
rect 30929 15447 30987 15453
rect 31754 15444 31760 15456
rect 31812 15444 31818 15496
rect 33318 15484 33324 15496
rect 33279 15456 33324 15484
rect 33318 15444 33324 15456
rect 33376 15444 33382 15496
rect 33597 15487 33655 15493
rect 33597 15453 33609 15487
rect 33643 15484 33655 15487
rect 33686 15484 33692 15496
rect 33643 15456 33692 15484
rect 33643 15453 33655 15456
rect 33597 15447 33655 15453
rect 33686 15444 33692 15456
rect 33744 15444 33750 15496
rect 35345 15487 35403 15493
rect 35345 15453 35357 15487
rect 35391 15453 35403 15487
rect 38194 15484 38200 15496
rect 38155 15456 38200 15484
rect 35345 15447 35403 15453
rect 35360 15416 35388 15447
rect 38194 15444 38200 15456
rect 38252 15444 38258 15496
rect 38396 15493 38424 15524
rect 38488 15493 38516 15592
rect 41049 15555 41107 15561
rect 41049 15552 41061 15555
rect 40144 15524 41061 15552
rect 38381 15487 38439 15493
rect 38381 15453 38393 15487
rect 38427 15453 38439 15487
rect 38381 15447 38439 15453
rect 38473 15487 38531 15493
rect 38473 15453 38485 15487
rect 38519 15453 38531 15487
rect 38473 15447 38531 15453
rect 38562 15444 38568 15496
rect 38620 15484 38626 15496
rect 40144 15493 40172 15524
rect 41049 15521 41061 15524
rect 41095 15521 41107 15555
rect 41049 15515 41107 15521
rect 40129 15487 40187 15493
rect 40129 15484 40141 15487
rect 38620 15456 40141 15484
rect 38620 15444 38626 15456
rect 40129 15453 40141 15456
rect 40175 15453 40187 15487
rect 40129 15447 40187 15453
rect 40218 15484 40276 15490
rect 40497 15487 40555 15493
rect 40218 15450 40230 15484
rect 40264 15450 40276 15484
rect 40218 15444 40276 15450
rect 40313 15481 40371 15487
rect 40313 15447 40325 15481
rect 40359 15447 40371 15481
rect 40497 15453 40509 15487
rect 40543 15484 40555 15487
rect 40954 15484 40960 15496
rect 40543 15456 40960 15484
rect 40543 15453 40555 15456
rect 40497 15447 40555 15453
rect 35434 15416 35440 15428
rect 27356 15388 35440 15416
rect 35434 15376 35440 15388
rect 35492 15376 35498 15428
rect 37182 15376 37188 15428
rect 37240 15416 37246 15428
rect 37369 15419 37427 15425
rect 37369 15416 37381 15419
rect 37240 15388 37381 15416
rect 37240 15376 37246 15388
rect 37369 15385 37381 15388
rect 37415 15385 37427 15419
rect 37369 15379 37427 15385
rect 37553 15419 37611 15425
rect 37553 15385 37565 15419
rect 37599 15416 37611 15419
rect 38654 15416 38660 15428
rect 37599 15388 38660 15416
rect 37599 15385 37611 15388
rect 37553 15379 37611 15385
rect 38654 15376 38660 15388
rect 38712 15376 38718 15428
rect 39942 15376 39948 15428
rect 40000 15416 40006 15428
rect 40233 15416 40261 15444
rect 40313 15441 40371 15447
rect 40954 15444 40960 15456
rect 41012 15444 41018 15496
rect 40000 15388 40261 15416
rect 40000 15376 40006 15388
rect 21692 15320 23244 15348
rect 26881 15351 26939 15357
rect 21692 15308 21698 15320
rect 26881 15317 26893 15351
rect 26927 15348 26939 15351
rect 27522 15348 27528 15360
rect 26927 15320 27528 15348
rect 26927 15317 26939 15320
rect 26881 15311 26939 15317
rect 27522 15308 27528 15320
rect 27580 15308 27586 15360
rect 32861 15351 32919 15357
rect 32861 15317 32873 15351
rect 32907 15348 32919 15351
rect 33318 15348 33324 15360
rect 32907 15320 33324 15348
rect 32907 15317 32919 15320
rect 32861 15311 32919 15317
rect 33318 15308 33324 15320
rect 33376 15348 33382 15360
rect 33594 15348 33600 15360
rect 33376 15320 33600 15348
rect 33376 15308 33382 15320
rect 33594 15308 33600 15320
rect 33652 15308 33658 15360
rect 38838 15348 38844 15360
rect 38799 15320 38844 15348
rect 38838 15308 38844 15320
rect 38896 15308 38902 15360
rect 40218 15308 40224 15360
rect 40276 15348 40282 15360
rect 40328 15348 40356 15441
rect 40276 15320 40356 15348
rect 40276 15308 40282 15320
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 4982 15104 4988 15156
rect 5040 15144 5046 15156
rect 6914 15144 6920 15156
rect 5040 15116 6920 15144
rect 5040 15104 5046 15116
rect 6914 15104 6920 15116
rect 6972 15144 6978 15156
rect 7282 15144 7288 15156
rect 6972 15116 7144 15144
rect 7243 15116 7288 15144
rect 6972 15104 6978 15116
rect 5442 15036 5448 15088
rect 5500 15076 5506 15088
rect 5500 15048 6868 15076
rect 5500 15036 5506 15048
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 3694 15017 3700 15020
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 2004 14980 3433 15008
rect 2004 14968 2010 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3688 14971 3700 15017
rect 3752 15008 3758 15020
rect 6840 15017 6868 15048
rect 7116 15017 7144 15116
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 12710 15144 12716 15156
rect 8128 15116 12716 15144
rect 8128 15017 8156 15116
rect 12710 15104 12716 15116
rect 12768 15104 12774 15156
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14550 15144 14556 15156
rect 14047 15116 14556 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 14660 15116 20484 15144
rect 13078 15076 13084 15088
rect 10060 15048 10548 15076
rect 6549 15011 6607 15017
rect 3752 14980 3788 15008
rect 3694 14968 3700 14971
rect 3752 14968 3758 14980
rect 6549 14977 6561 15011
rect 6595 15008 6607 15011
rect 6733 15011 6791 15017
rect 6595 14980 6684 15008
rect 6595 14977 6607 14980
rect 6549 14971 6607 14977
rect 4801 14807 4859 14813
rect 4801 14773 4813 14807
rect 4847 14804 4859 14807
rect 5626 14804 5632 14816
rect 4847 14776 5632 14804
rect 4847 14773 4859 14776
rect 4801 14767 4859 14773
rect 5626 14764 5632 14776
rect 5684 14764 5690 14816
rect 6656 14804 6684 14980
rect 6733 14977 6745 15011
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6825 14971 6883 14977
rect 7101 15011 7159 15017
rect 7101 14977 7113 15011
rect 7147 14977 7159 15011
rect 7101 14971 7159 14977
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 6748 14872 6776 14971
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14940 6975 14943
rect 7190 14940 7196 14952
rect 6963 14912 7196 14940
rect 6963 14909 6975 14912
rect 6917 14903 6975 14909
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 10060 14940 10088 15048
rect 10226 15008 10232 15020
rect 10187 14980 10232 15008
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 14977 10471 15011
rect 10413 14971 10471 14977
rect 10318 14940 10324 14952
rect 8067 14912 10088 14940
rect 10279 14912 10324 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 10318 14900 10324 14912
rect 10376 14900 10382 14952
rect 10428 14884 10456 14971
rect 7745 14875 7803 14881
rect 7745 14872 7757 14875
rect 6748 14844 7757 14872
rect 7745 14841 7757 14844
rect 7791 14841 7803 14875
rect 10410 14872 10416 14884
rect 7745 14835 7803 14841
rect 9692 14844 10416 14872
rect 6914 14804 6920 14816
rect 6656 14776 6920 14804
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 7926 14804 7932 14816
rect 7887 14776 7932 14804
rect 7926 14764 7932 14776
rect 7984 14764 7990 14816
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 9692 14813 9720 14844
rect 10410 14832 10416 14844
rect 10468 14832 10474 14884
rect 10520 14872 10548 15048
rect 12636 15048 13084 15076
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 12636 15017 12664 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12124 14980 12449 15008
rect 12124 14968 12130 14980
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12585 15011 12664 15017
rect 12585 14977 12597 15011
rect 12631 14980 12664 15011
rect 12713 15011 12771 15017
rect 12631 14977 12643 14980
rect 12585 14971 12643 14977
rect 12713 14977 12725 15011
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 12728 14940 12756 14971
rect 12802 14968 12808 15020
rect 12860 15008 12866 15020
rect 12986 15017 12992 15020
rect 12943 15011 12992 15017
rect 12860 14980 12905 15008
rect 12860 14968 12866 14980
rect 12943 14977 12955 15011
rect 12989 14977 12992 15011
rect 12943 14971 12992 14977
rect 12958 14968 12992 14971
rect 13044 15008 13050 15020
rect 13044 14980 13091 15008
rect 13044 14968 13050 14980
rect 12636 14912 12756 14940
rect 12958 14940 12986 14968
rect 13998 14940 14004 14952
rect 12958 14912 14004 14940
rect 12526 14872 12532 14884
rect 10520 14844 12532 14872
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 12636 14816 12664 14912
rect 13998 14900 14004 14912
rect 14056 14940 14062 14952
rect 14660 14940 14688 15116
rect 16022 15076 16028 15088
rect 15983 15048 16028 15076
rect 16022 15036 16028 15048
rect 16080 15036 16086 15088
rect 16758 15036 16764 15088
rect 16816 15076 16822 15088
rect 19242 15076 19248 15088
rect 16816 15048 19248 15076
rect 16816 15036 16822 15048
rect 16040 15008 16068 15036
rect 16666 15008 16672 15020
rect 16040 14980 16672 15008
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 18064 15017 18092 15048
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 18322 15017 18328 15020
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18316 15008 18328 15017
rect 18283 14980 18328 15008
rect 18049 14971 18107 14977
rect 18316 14971 18328 14980
rect 14056 14912 14688 14940
rect 14056 14900 14062 14912
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 16868 14940 16896 14971
rect 18322 14968 18328 14971
rect 18380 14968 18386 15020
rect 20162 14968 20168 15020
rect 20220 15008 20226 15020
rect 20456 15017 20484 15116
rect 20990 15104 20996 15156
rect 21048 15144 21054 15156
rect 21085 15147 21143 15153
rect 21085 15144 21097 15147
rect 21048 15116 21097 15144
rect 21048 15104 21054 15116
rect 21085 15113 21097 15116
rect 21131 15144 21143 15147
rect 21542 15144 21548 15156
rect 21131 15116 21548 15144
rect 21131 15113 21143 15116
rect 21085 15107 21143 15113
rect 21542 15104 21548 15116
rect 21600 15104 21606 15156
rect 26234 15144 26240 15156
rect 21652 15116 26240 15144
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 20220 14980 20269 15008
rect 20220 14968 20226 14980
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 15008 20499 15011
rect 20901 15011 20959 15017
rect 20901 15008 20913 15011
rect 20487 14980 20913 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 20901 14977 20913 14980
rect 20947 14977 20959 15011
rect 20901 14971 20959 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 15008 21143 15011
rect 21174 15008 21180 15020
rect 21131 14980 21180 15008
rect 21131 14977 21143 14980
rect 21085 14971 21143 14977
rect 21174 14968 21180 14980
rect 21232 15008 21238 15020
rect 21652 15008 21680 15116
rect 26234 15104 26240 15116
rect 26292 15144 26298 15156
rect 30009 15147 30067 15153
rect 26292 15116 28994 15144
rect 26292 15104 26298 15116
rect 21232 14980 21680 15008
rect 21744 15048 22784 15076
rect 21232 14968 21238 14980
rect 16356 14912 16896 14940
rect 16356 14900 16362 14912
rect 12710 14832 12716 14884
rect 12768 14872 12774 14884
rect 13081 14875 13139 14881
rect 13081 14872 13093 14875
rect 12768 14844 13093 14872
rect 12768 14832 12774 14844
rect 13081 14841 13093 14844
rect 13127 14841 13139 14875
rect 13081 14835 13139 14841
rect 16853 14875 16911 14881
rect 16853 14841 16865 14875
rect 16899 14872 16911 14875
rect 17126 14872 17132 14884
rect 16899 14844 17132 14872
rect 16899 14841 16911 14844
rect 16853 14835 16911 14841
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 19426 14872 19432 14884
rect 19339 14844 19432 14872
rect 19426 14832 19432 14844
rect 19484 14872 19490 14884
rect 21744 14872 21772 15048
rect 22186 14968 22192 15020
rect 22244 15008 22250 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 22244 14980 22293 15008
rect 22244 14968 22250 14980
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22281 14971 22339 14977
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 15008 22523 15011
rect 22646 15008 22652 15020
rect 22511 14980 22652 15008
rect 22511 14977 22523 14980
rect 22465 14971 22523 14977
rect 22646 14968 22652 14980
rect 22704 14968 22710 15020
rect 22756 15008 22784 15048
rect 22830 15036 22836 15088
rect 22888 15076 22894 15088
rect 23106 15076 23112 15088
rect 22888 15048 23112 15076
rect 22888 15036 22894 15048
rect 23106 15036 23112 15048
rect 23164 15036 23170 15088
rect 23201 15079 23259 15085
rect 23201 15045 23213 15079
rect 23247 15076 23259 15079
rect 26602 15076 26608 15088
rect 23247 15048 26608 15076
rect 23247 15045 23259 15048
rect 23201 15039 23259 15045
rect 26602 15036 26608 15048
rect 26660 15036 26666 15088
rect 27246 15036 27252 15088
rect 27304 15076 27310 15088
rect 27341 15079 27399 15085
rect 27341 15076 27353 15079
rect 27304 15048 27353 15076
rect 27304 15036 27310 15048
rect 27341 15045 27353 15048
rect 27387 15076 27399 15079
rect 28166 15076 28172 15088
rect 27387 15048 28172 15076
rect 27387 15045 27399 15048
rect 27341 15039 27399 15045
rect 28166 15036 28172 15048
rect 28224 15076 28230 15088
rect 28626 15076 28632 15088
rect 28224 15048 28632 15076
rect 28224 15036 28230 15048
rect 28626 15036 28632 15048
rect 28684 15036 28690 15088
rect 28966 15076 28994 15116
rect 30009 15113 30021 15147
rect 30055 15144 30067 15147
rect 30374 15144 30380 15156
rect 30055 15116 30380 15144
rect 30055 15113 30067 15116
rect 30009 15107 30067 15113
rect 30374 15104 30380 15116
rect 30432 15104 30438 15156
rect 36081 15147 36139 15153
rect 36081 15113 36093 15147
rect 36127 15144 36139 15147
rect 36127 15116 37780 15144
rect 36127 15113 36139 15116
rect 36081 15107 36139 15113
rect 37752 15076 37780 15116
rect 38654 15104 38660 15156
rect 38712 15144 38718 15156
rect 40221 15147 40279 15153
rect 40221 15144 40233 15147
rect 38712 15116 40233 15144
rect 38712 15104 38718 15116
rect 40221 15113 40233 15116
rect 40267 15113 40279 15147
rect 40221 15107 40279 15113
rect 37826 15076 37832 15088
rect 28966 15048 36124 15076
rect 37739 15048 37832 15076
rect 22925 15011 22983 15017
rect 22925 15008 22937 15011
rect 22756 14980 22937 15008
rect 22925 14977 22937 14980
rect 22971 14977 22983 15011
rect 23290 15008 23296 15020
rect 23251 14980 23296 15008
rect 22925 14971 22983 14977
rect 23290 14968 23296 14980
rect 23348 14968 23354 15020
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 15008 24271 15011
rect 24394 15008 24400 15020
rect 24259 14980 24400 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24394 14968 24400 14980
rect 24452 14968 24458 15020
rect 24489 15014 24547 15017
rect 24489 15011 24624 15014
rect 24489 14977 24501 15011
rect 24535 15008 24624 15011
rect 27525 15011 27583 15017
rect 24535 14986 25084 15008
rect 24535 14977 24547 14986
rect 24596 14980 25084 14986
rect 24489 14971 24547 14977
rect 25056 14952 25084 14980
rect 27525 14977 27537 15011
rect 27571 14977 27583 15011
rect 27525 14971 27583 14977
rect 23198 14900 23204 14952
rect 23256 14940 23262 14952
rect 24305 14943 24363 14949
rect 24305 14940 24317 14943
rect 23256 14912 24317 14940
rect 23256 14900 23262 14912
rect 24305 14909 24317 14912
rect 24351 14909 24363 14943
rect 25038 14940 25044 14952
rect 24999 14912 25044 14940
rect 24305 14903 24363 14909
rect 25038 14900 25044 14912
rect 25096 14900 25102 14952
rect 25498 14900 25504 14952
rect 25556 14940 25562 14952
rect 27540 14940 27568 14971
rect 29546 14968 29552 15020
rect 29604 15008 29610 15020
rect 30285 15011 30343 15017
rect 30285 15008 30297 15011
rect 29604 14980 30297 15008
rect 29604 14968 29610 14980
rect 30285 14977 30297 14980
rect 30331 14977 30343 15011
rect 30285 14971 30343 14977
rect 30377 15011 30435 15017
rect 30377 14977 30389 15011
rect 30423 14977 30435 15011
rect 30377 14971 30435 14977
rect 28350 14940 28356 14952
rect 25556 14912 28356 14940
rect 25556 14900 25562 14912
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 29914 14900 29920 14952
rect 29972 14940 29978 14952
rect 30392 14940 30420 14971
rect 30466 14968 30472 15020
rect 30524 15008 30530 15020
rect 30653 15011 30711 15017
rect 30524 14980 30569 15008
rect 30524 14968 30530 14980
rect 30653 14977 30665 15011
rect 30699 15008 30711 15011
rect 33321 15011 33379 15017
rect 33321 15008 33333 15011
rect 30699 14980 33333 15008
rect 30699 14977 30711 14980
rect 30653 14971 30711 14977
rect 33321 14977 33333 14980
rect 33367 15008 33379 15011
rect 33410 15008 33416 15020
rect 33367 14980 33416 15008
rect 33367 14977 33379 14980
rect 33321 14971 33379 14977
rect 29972 14912 30420 14940
rect 29972 14900 29978 14912
rect 19484 14844 21772 14872
rect 22465 14875 22523 14881
rect 19484 14832 19490 14844
rect 22465 14841 22477 14875
rect 22511 14872 22523 14875
rect 27982 14872 27988 14884
rect 22511 14844 27988 14872
rect 22511 14841 22523 14844
rect 22465 14835 22523 14841
rect 27982 14832 27988 14844
rect 28040 14832 28046 14884
rect 29454 14832 29460 14884
rect 29512 14872 29518 14884
rect 29512 14844 30236 14872
rect 29512 14832 29518 14844
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 8812 14776 9689 14804
rect 8812 14764 8818 14776
rect 9677 14773 9689 14776
rect 9723 14773 9735 14807
rect 9677 14767 9735 14773
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10873 14807 10931 14813
rect 10873 14804 10885 14807
rect 10284 14776 10885 14804
rect 10284 14764 10290 14776
rect 10873 14773 10885 14776
rect 10919 14773 10931 14807
rect 10873 14767 10931 14773
rect 12618 14764 12624 14816
rect 12676 14764 12682 14816
rect 14366 14764 14372 14816
rect 14424 14804 14430 14816
rect 17497 14807 17555 14813
rect 17497 14804 17509 14807
rect 14424 14776 17509 14804
rect 14424 14764 14430 14776
rect 17497 14773 17509 14776
rect 17543 14804 17555 14807
rect 18414 14804 18420 14816
rect 17543 14776 18420 14804
rect 17543 14773 17555 14776
rect 17497 14767 17555 14773
rect 18414 14764 18420 14776
rect 18472 14764 18478 14816
rect 21358 14764 21364 14816
rect 21416 14804 21422 14816
rect 22186 14804 22192 14816
rect 21416 14776 22192 14804
rect 21416 14764 21422 14776
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 22554 14764 22560 14816
rect 22612 14804 22618 14816
rect 23290 14804 23296 14816
rect 22612 14776 23296 14804
rect 22612 14764 22618 14776
rect 23290 14764 23296 14776
rect 23348 14764 23354 14816
rect 23474 14804 23480 14816
rect 23435 14776 23480 14804
rect 23474 14764 23480 14776
rect 23532 14764 23538 14816
rect 24026 14804 24032 14816
rect 23987 14776 24032 14804
rect 24026 14764 24032 14776
rect 24084 14764 24090 14816
rect 24210 14804 24216 14816
rect 24171 14776 24216 14804
rect 24210 14764 24216 14776
rect 24268 14764 24274 14816
rect 24302 14764 24308 14816
rect 24360 14804 24366 14816
rect 25501 14807 25559 14813
rect 25501 14804 25513 14807
rect 24360 14776 25513 14804
rect 24360 14764 24366 14776
rect 25501 14773 25513 14776
rect 25547 14773 25559 14807
rect 25501 14767 25559 14773
rect 27709 14807 27767 14813
rect 27709 14773 27721 14807
rect 27755 14804 27767 14807
rect 27798 14804 27804 14816
rect 27755 14776 27804 14804
rect 27755 14773 27767 14776
rect 27709 14767 27767 14773
rect 27798 14764 27804 14776
rect 27856 14764 27862 14816
rect 29546 14804 29552 14816
rect 29507 14776 29552 14804
rect 29546 14764 29552 14776
rect 29604 14764 29610 14816
rect 30208 14804 30236 14844
rect 30668 14804 30696 14971
rect 33410 14968 33416 14980
rect 33468 14968 33474 15020
rect 35434 15008 35440 15020
rect 35395 14980 35440 15008
rect 35434 14968 35440 14980
rect 35492 14968 35498 15020
rect 36096 15017 36124 15048
rect 37826 15036 37832 15048
rect 37884 15036 37890 15088
rect 38838 15036 38844 15088
rect 38896 15076 38902 15088
rect 39086 15079 39144 15085
rect 39086 15076 39098 15079
rect 38896 15048 39098 15076
rect 38896 15036 38902 15048
rect 39086 15045 39098 15048
rect 39132 15045 39144 15079
rect 39086 15039 39144 15045
rect 35897 15011 35955 15017
rect 35897 14977 35909 15011
rect 35943 14977 35955 15011
rect 35897 14971 35955 14977
rect 36081 15011 36139 15017
rect 36081 14977 36093 15011
rect 36127 15008 36139 15011
rect 36541 15011 36599 15017
rect 36541 15008 36553 15011
rect 36127 14980 36553 15008
rect 36127 14977 36139 14980
rect 36081 14971 36139 14977
rect 36541 14977 36553 14980
rect 36587 15008 36599 15011
rect 36722 15008 36728 15020
rect 36587 14980 36728 15008
rect 36587 14977 36599 14980
rect 36541 14971 36599 14977
rect 33597 14943 33655 14949
rect 33597 14909 33609 14943
rect 33643 14940 33655 14943
rect 33686 14940 33692 14952
rect 33643 14912 33692 14940
rect 33643 14909 33655 14912
rect 33597 14903 33655 14909
rect 30208 14776 30696 14804
rect 33612 14804 33640 14903
rect 33686 14900 33692 14912
rect 33744 14900 33750 14952
rect 35161 14943 35219 14949
rect 35161 14909 35173 14943
rect 35207 14940 35219 14943
rect 35912 14940 35940 14971
rect 36722 14968 36728 14980
rect 36780 14968 36786 15020
rect 35207 14912 35940 14940
rect 35207 14909 35219 14912
rect 35161 14903 35219 14909
rect 35452 14884 35480 14912
rect 38654 14900 38660 14952
rect 38712 14940 38718 14952
rect 38841 14943 38899 14949
rect 38841 14940 38853 14943
rect 38712 14912 38853 14940
rect 38712 14900 38718 14912
rect 38841 14909 38853 14912
rect 38887 14909 38899 14943
rect 38841 14903 38899 14909
rect 35434 14832 35440 14884
rect 35492 14832 35498 14884
rect 37642 14872 37648 14884
rect 37603 14844 37648 14872
rect 37642 14832 37648 14844
rect 37700 14832 37706 14884
rect 35986 14804 35992 14816
rect 33612 14776 35992 14804
rect 35986 14764 35992 14776
rect 36044 14764 36050 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 3053 14603 3111 14609
rect 3053 14600 3065 14603
rect 2832 14572 3065 14600
rect 2832 14560 2838 14572
rect 3053 14569 3065 14572
rect 3099 14569 3111 14603
rect 3053 14563 3111 14569
rect 3694 14560 3700 14612
rect 3752 14600 3758 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3752 14572 3801 14600
rect 3752 14560 3758 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 12860 14572 14105 14600
rect 12860 14560 12866 14572
rect 14093 14569 14105 14572
rect 14139 14600 14151 14603
rect 14458 14600 14464 14612
rect 14139 14572 14464 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 17954 14600 17960 14612
rect 17867 14572 17960 14600
rect 17954 14560 17960 14572
rect 18012 14600 18018 14612
rect 23569 14603 23627 14609
rect 18012 14572 23060 14600
rect 18012 14560 18018 14572
rect 1578 14492 1584 14544
rect 1636 14532 1642 14544
rect 7650 14532 7656 14544
rect 1636 14504 7656 14532
rect 1636 14492 1642 14504
rect 7650 14492 7656 14504
rect 7708 14492 7714 14544
rect 10410 14492 10416 14544
rect 10468 14532 10474 14544
rect 14366 14532 14372 14544
rect 10468 14504 14372 14532
rect 10468 14492 10474 14504
rect 14366 14492 14372 14504
rect 14424 14492 14430 14544
rect 18138 14492 18144 14544
rect 18196 14532 18202 14544
rect 18196 14504 22048 14532
rect 18196 14492 18202 14504
rect 18414 14424 18420 14476
rect 18472 14464 18478 14476
rect 18601 14467 18659 14473
rect 18601 14464 18613 14467
rect 18472 14436 18613 14464
rect 18472 14424 18478 14436
rect 18601 14433 18613 14436
rect 18647 14464 18659 14467
rect 20162 14464 20168 14476
rect 18647 14436 19656 14464
rect 20123 14436 20168 14464
rect 18647 14433 18659 14436
rect 18601 14427 18659 14433
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14365 3295 14399
rect 3970 14396 3976 14408
rect 3931 14368 3976 14396
rect 3237 14359 3295 14365
rect 3252 14328 3280 14359
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9646 14368 9873 14396
rect 4798 14328 4804 14340
rect 3252 14300 4804 14328
rect 4798 14288 4804 14300
rect 4856 14288 4862 14340
rect 8938 14288 8944 14340
rect 8996 14328 9002 14340
rect 9646 14328 9674 14368
rect 9861 14365 9873 14368
rect 9907 14396 9919 14399
rect 11790 14396 11796 14408
rect 9907 14368 11796 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 11790 14356 11796 14368
rect 11848 14396 11854 14408
rect 12425 14399 12483 14405
rect 12425 14396 12437 14399
rect 11848 14368 12437 14396
rect 11848 14356 11854 14368
rect 12425 14365 12437 14368
rect 12471 14365 12483 14399
rect 12425 14359 12483 14365
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 16577 14399 16635 14405
rect 16577 14396 16589 14399
rect 15519 14368 16589 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 16577 14365 16589 14368
rect 16623 14396 16635 14399
rect 16666 14396 16672 14408
rect 16623 14368 16672 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 16850 14405 16856 14408
rect 16844 14396 16856 14405
rect 16811 14368 16856 14396
rect 16844 14359 16856 14368
rect 16850 14356 16856 14359
rect 16908 14356 16914 14408
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19521 14399 19579 14405
rect 19521 14396 19533 14399
rect 19392 14368 19533 14396
rect 19392 14356 19398 14368
rect 19521 14365 19533 14368
rect 19567 14365 19579 14399
rect 19628 14396 19656 14436
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 21450 14464 21456 14476
rect 21411 14436 21456 14464
rect 21450 14424 21456 14436
rect 21508 14424 21514 14476
rect 19705 14399 19763 14405
rect 19705 14396 19717 14399
rect 19628 14368 19717 14396
rect 19521 14359 19579 14365
rect 19705 14365 19717 14368
rect 19751 14396 19763 14399
rect 19978 14396 19984 14408
rect 19751 14368 19984 14396
rect 19751 14365 19763 14368
rect 19705 14359 19763 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20070 14356 20076 14408
rect 20128 14396 20134 14408
rect 20254 14396 20260 14408
rect 20128 14368 20260 14396
rect 20128 14356 20134 14368
rect 20254 14356 20260 14368
rect 20312 14396 20318 14408
rect 22020 14405 22048 14504
rect 22738 14464 22744 14476
rect 22204 14436 22744 14464
rect 22204 14405 22232 14436
rect 22738 14424 22744 14436
rect 22796 14424 22802 14476
rect 20441 14399 20499 14405
rect 20441 14396 20453 14399
rect 20312 14368 20453 14396
rect 20312 14356 20318 14368
rect 20441 14365 20453 14368
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22189 14399 22247 14405
rect 22189 14365 22201 14399
rect 22235 14365 22247 14399
rect 22189 14359 22247 14365
rect 22373 14399 22431 14405
rect 22373 14365 22385 14399
rect 22419 14396 22431 14399
rect 22554 14396 22560 14408
rect 22419 14368 22560 14396
rect 22419 14365 22431 14368
rect 22373 14359 22431 14365
rect 22554 14356 22560 14368
rect 22612 14356 22618 14408
rect 23032 14405 23060 14572
rect 23569 14569 23581 14603
rect 23615 14600 23627 14603
rect 24210 14600 24216 14612
rect 23615 14572 24216 14600
rect 23615 14569 23627 14572
rect 23569 14563 23627 14569
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 24486 14600 24492 14612
rect 24447 14572 24492 14600
rect 24486 14560 24492 14572
rect 24544 14560 24550 14612
rect 25133 14603 25191 14609
rect 25133 14569 25145 14603
rect 25179 14600 25191 14603
rect 26602 14600 26608 14612
rect 25179 14572 26608 14600
rect 25179 14569 25191 14572
rect 25133 14563 25191 14569
rect 26602 14560 26608 14572
rect 26660 14560 26666 14612
rect 27706 14560 27712 14612
rect 27764 14600 27770 14612
rect 30374 14600 30380 14612
rect 27764 14572 30380 14600
rect 27764 14560 27770 14572
rect 30374 14560 30380 14572
rect 30432 14600 30438 14612
rect 30561 14603 30619 14609
rect 30561 14600 30573 14603
rect 30432 14572 30573 14600
rect 30432 14560 30438 14572
rect 30561 14569 30573 14572
rect 30607 14569 30619 14603
rect 30561 14563 30619 14569
rect 31726 14572 37044 14600
rect 23658 14492 23664 14544
rect 23716 14532 23722 14544
rect 24504 14532 24532 14560
rect 28350 14532 28356 14544
rect 23716 14504 24532 14532
rect 28311 14504 28356 14532
rect 23716 14492 23722 14504
rect 28350 14492 28356 14504
rect 28408 14492 28414 14544
rect 29178 14492 29184 14544
rect 29236 14532 29242 14544
rect 31726 14532 31754 14572
rect 29236 14504 31754 14532
rect 29236 14492 29242 14504
rect 25498 14464 25504 14476
rect 23308 14436 25504 14464
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 23106 14356 23112 14408
rect 23164 14396 23170 14408
rect 23308 14405 23336 14436
rect 25498 14424 25504 14436
rect 25556 14424 25562 14476
rect 26510 14464 26516 14476
rect 26471 14436 26516 14464
rect 26510 14424 26516 14436
rect 26568 14464 26574 14476
rect 26973 14467 27031 14473
rect 26973 14464 26985 14467
rect 26568 14436 26985 14464
rect 26568 14424 26574 14436
rect 26973 14433 26985 14436
rect 27019 14433 27031 14467
rect 26973 14427 27031 14433
rect 27982 14424 27988 14476
rect 28040 14464 28046 14476
rect 35526 14464 35532 14476
rect 28040 14436 35532 14464
rect 28040 14424 28046 14436
rect 35526 14424 35532 14436
rect 35584 14464 35590 14476
rect 35621 14467 35679 14473
rect 35621 14464 35633 14467
rect 35584 14436 35633 14464
rect 35584 14424 35590 14436
rect 35621 14433 35633 14436
rect 35667 14433 35679 14467
rect 37016 14464 37044 14572
rect 37734 14560 37740 14612
rect 37792 14600 37798 14612
rect 38930 14600 38936 14612
rect 37792 14572 38936 14600
rect 37792 14560 37798 14572
rect 38930 14560 38936 14572
rect 38988 14560 38994 14612
rect 40126 14560 40132 14612
rect 40184 14600 40190 14612
rect 40405 14603 40463 14609
rect 40405 14600 40417 14603
rect 40184 14572 40417 14600
rect 40184 14560 40190 14572
rect 40405 14569 40417 14572
rect 40451 14569 40463 14603
rect 40405 14563 40463 14569
rect 38381 14467 38439 14473
rect 38381 14464 38393 14467
rect 37016 14436 38393 14464
rect 35621 14427 35679 14433
rect 38381 14433 38393 14436
rect 38427 14464 38439 14467
rect 38930 14464 38936 14476
rect 38427 14436 38936 14464
rect 38427 14433 38439 14436
rect 38381 14427 38439 14433
rect 38930 14424 38936 14436
rect 38988 14424 38994 14476
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 23164 14368 23213 14396
rect 23164 14356 23170 14368
rect 23201 14365 23213 14368
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 23293 14399 23351 14405
rect 23293 14365 23305 14399
rect 23339 14365 23351 14399
rect 23293 14359 23351 14365
rect 23382 14356 23388 14408
rect 23440 14396 23446 14408
rect 23440 14368 23485 14396
rect 23440 14356 23446 14368
rect 24854 14356 24860 14408
rect 24912 14396 24918 14408
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 24912 14368 29561 14396
rect 24912 14356 24918 14368
rect 29549 14365 29561 14368
rect 29595 14396 29607 14399
rect 29822 14396 29828 14408
rect 29595 14368 29828 14396
rect 29595 14365 29607 14368
rect 29549 14359 29607 14365
rect 29822 14356 29828 14368
rect 29880 14356 29886 14408
rect 35158 14396 35164 14408
rect 29932 14368 35164 14396
rect 15194 14328 15200 14340
rect 15252 14337 15258 14340
rect 8996 14300 9674 14328
rect 12544 14300 15056 14328
rect 15164 14300 15200 14328
rect 8996 14288 9002 14300
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 7282 14260 7288 14272
rect 6972 14232 7288 14260
rect 6972 14220 6978 14232
rect 7282 14220 7288 14232
rect 7340 14260 7346 14272
rect 7469 14263 7527 14269
rect 7469 14260 7481 14263
rect 7340 14232 7481 14260
rect 7340 14220 7346 14232
rect 7469 14229 7481 14232
rect 7515 14260 7527 14263
rect 9953 14263 10011 14269
rect 9953 14260 9965 14263
rect 7515 14232 9965 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 9953 14229 9965 14232
rect 9999 14229 10011 14263
rect 9953 14223 10011 14229
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 12544 14260 12572 14300
rect 10284 14232 12572 14260
rect 12621 14263 12679 14269
rect 10284 14220 10290 14232
rect 12621 14229 12633 14263
rect 12667 14260 12679 14263
rect 12894 14260 12900 14272
rect 12667 14232 12900 14260
rect 12667 14229 12679 14232
rect 12621 14223 12679 14229
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 15028 14260 15056 14300
rect 15194 14288 15200 14300
rect 15252 14291 15264 14337
rect 21358 14328 21364 14340
rect 18524 14300 21364 14328
rect 15252 14288 15258 14291
rect 18524 14260 18552 14300
rect 21358 14288 21364 14300
rect 21416 14288 21422 14340
rect 22281 14331 22339 14337
rect 22281 14297 22293 14331
rect 22327 14328 22339 14331
rect 26268 14331 26326 14337
rect 22327 14300 23244 14328
rect 22327 14297 22339 14300
rect 22281 14291 22339 14297
rect 15028 14232 18552 14260
rect 19613 14263 19671 14269
rect 19613 14229 19625 14263
rect 19659 14260 19671 14263
rect 20162 14260 20168 14272
rect 19659 14232 20168 14260
rect 19659 14229 19671 14232
rect 19613 14223 19671 14229
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 22557 14263 22615 14269
rect 22557 14229 22569 14263
rect 22603 14260 22615 14263
rect 23106 14260 23112 14272
rect 22603 14232 23112 14260
rect 22603 14229 22615 14232
rect 22557 14223 22615 14229
rect 23106 14220 23112 14232
rect 23164 14220 23170 14272
rect 23216 14260 23244 14300
rect 24320 14300 26188 14328
rect 24320 14260 24348 14300
rect 23216 14232 24348 14260
rect 26160 14260 26188 14300
rect 26268 14297 26280 14331
rect 26314 14328 26326 14331
rect 27062 14328 27068 14340
rect 26314 14300 27068 14328
rect 26314 14297 26326 14300
rect 26268 14291 26326 14297
rect 27062 14288 27068 14300
rect 27120 14288 27126 14340
rect 27246 14337 27252 14340
rect 27240 14291 27252 14337
rect 27304 14328 27310 14340
rect 27304 14300 27340 14328
rect 27246 14288 27252 14291
rect 27304 14288 27310 14300
rect 27430 14288 27436 14340
rect 27488 14328 27494 14340
rect 29932 14328 29960 14368
rect 35158 14356 35164 14368
rect 35216 14356 35222 14408
rect 35342 14396 35348 14408
rect 35303 14368 35348 14396
rect 35342 14356 35348 14368
rect 35400 14356 35406 14408
rect 36170 14396 36176 14408
rect 36131 14368 36176 14396
rect 36170 14356 36176 14368
rect 36228 14356 36234 14408
rect 40313 14399 40371 14405
rect 40313 14365 40325 14399
rect 40359 14396 40371 14399
rect 40678 14396 40684 14408
rect 40359 14368 40684 14396
rect 40359 14365 40371 14368
rect 40313 14359 40371 14365
rect 40678 14356 40684 14368
rect 40736 14356 40742 14408
rect 58158 14396 58164 14408
rect 58119 14368 58164 14396
rect 58158 14356 58164 14368
rect 58216 14356 58222 14408
rect 27488 14300 29960 14328
rect 27488 14288 27494 14300
rect 30374 14288 30380 14340
rect 30432 14328 30438 14340
rect 32861 14331 32919 14337
rect 32861 14328 32873 14331
rect 30432 14300 32873 14328
rect 30432 14288 30438 14300
rect 32861 14297 32873 14300
rect 32907 14328 32919 14331
rect 36188 14328 36216 14356
rect 32907 14300 36216 14328
rect 32907 14297 32919 14300
rect 32861 14291 32919 14297
rect 28810 14260 28816 14272
rect 26160 14232 28816 14260
rect 28810 14220 28816 14232
rect 28868 14220 28874 14272
rect 31573 14263 31631 14269
rect 31573 14229 31585 14263
rect 31619 14260 31631 14263
rect 31754 14260 31760 14272
rect 31619 14232 31760 14260
rect 31619 14229 31631 14232
rect 31573 14223 31631 14229
rect 31754 14220 31760 14232
rect 31812 14220 31818 14272
rect 34514 14220 34520 14272
rect 34572 14260 34578 14272
rect 37461 14263 37519 14269
rect 37461 14260 37473 14263
rect 34572 14232 37473 14260
rect 34572 14220 34578 14232
rect 37461 14229 37473 14232
rect 37507 14260 37519 14263
rect 38654 14260 38660 14272
rect 37507 14232 38660 14260
rect 37507 14229 37519 14232
rect 37461 14223 37519 14229
rect 38654 14220 38660 14232
rect 38712 14220 38718 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 3145 14059 3203 14065
rect 3145 14025 3157 14059
rect 3191 14056 3203 14059
rect 3970 14056 3976 14068
rect 3191 14028 3976 14056
rect 3191 14025 3203 14028
rect 3145 14019 3203 14025
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 6604 14028 8493 14056
rect 6604 14016 6610 14028
rect 8481 14025 8493 14028
rect 8527 14056 8539 14059
rect 11054 14056 11060 14068
rect 8527 14028 11060 14056
rect 8527 14025 8539 14028
rect 8481 14019 8539 14025
rect 11054 14016 11060 14028
rect 11112 14016 11118 14068
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 23017 14059 23075 14065
rect 23017 14056 23029 14059
rect 12584 14028 23029 14056
rect 12584 14016 12590 14028
rect 23017 14025 23029 14028
rect 23063 14025 23075 14059
rect 23658 14056 23664 14068
rect 23017 14019 23075 14025
rect 23492 14028 23664 14056
rect 4798 13948 4804 14000
rect 4856 13988 4862 14000
rect 8938 13988 8944 14000
rect 4856 13960 8944 13988
rect 4856 13948 4862 13960
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 14458 13988 14464 14000
rect 14419 13960 14464 13988
rect 14458 13948 14464 13960
rect 14516 13948 14522 14000
rect 15838 13948 15844 14000
rect 15896 13988 15902 14000
rect 15896 13960 17724 13988
rect 15896 13948 15902 13960
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 2961 13923 3019 13929
rect 2832 13892 2877 13920
rect 2832 13880 2838 13892
rect 2961 13889 2973 13923
rect 3007 13920 3019 13923
rect 5166 13920 5172 13932
rect 3007 13892 5172 13920
rect 3007 13889 3019 13892
rect 2961 13883 3019 13889
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 5626 13880 5632 13932
rect 5684 13920 5690 13932
rect 6733 13923 6791 13929
rect 6733 13920 6745 13923
rect 5684 13892 6745 13920
rect 5684 13880 5690 13892
rect 6733 13889 6745 13892
rect 6779 13889 6791 13923
rect 6733 13883 6791 13889
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13964 13892 14289 13920
rect 13964 13880 13970 13892
rect 14277 13889 14289 13892
rect 14323 13920 14335 13923
rect 17696 13920 17724 13960
rect 17770 13948 17776 14000
rect 17828 13988 17834 14000
rect 19334 13988 19340 14000
rect 17828 13960 19340 13988
rect 17828 13948 17834 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 22281 13991 22339 13997
rect 19904 13960 22232 13988
rect 19904 13929 19932 13960
rect 18785 13923 18843 13929
rect 18785 13920 18797 13923
rect 14323 13892 17540 13920
rect 17696 13892 18797 13920
rect 14323 13889 14335 13892
rect 14277 13883 14335 13889
rect 17512 13864 17540 13892
rect 18785 13889 18797 13892
rect 18831 13920 18843 13923
rect 19889 13923 19947 13929
rect 19889 13920 19901 13923
rect 18831 13892 19901 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 19889 13889 19901 13892
rect 19935 13889 19947 13923
rect 20070 13920 20076 13932
rect 20031 13892 20076 13920
rect 19889 13883 19947 13889
rect 20070 13880 20076 13892
rect 20128 13880 20134 13932
rect 20901 13923 20959 13929
rect 20901 13889 20913 13923
rect 20947 13920 20959 13923
rect 22094 13920 22100 13932
rect 20947 13892 22100 13920
rect 20947 13889 20959 13892
rect 20901 13883 20959 13889
rect 5718 13812 5724 13864
rect 5776 13852 5782 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 5776 13824 6377 13852
rect 5776 13812 5782 13824
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 6822 13852 6828 13864
rect 6783 13824 6828 13852
rect 6365 13815 6423 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13852 7067 13855
rect 8018 13852 8024 13864
rect 7055 13824 8024 13852
rect 7055 13821 7067 13824
rect 7009 13815 7067 13821
rect 8018 13812 8024 13824
rect 8076 13812 8082 13864
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 16298 13852 16304 13864
rect 8628 13824 16304 13852
rect 8628 13812 8634 13824
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 17494 13812 17500 13864
rect 17552 13852 17558 13864
rect 17552 13824 19840 13852
rect 17552 13812 17558 13824
rect 12066 13744 12072 13796
rect 12124 13784 12130 13796
rect 15562 13784 15568 13796
rect 12124 13756 15568 13784
rect 12124 13744 12130 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 19812 13784 19840 13824
rect 20162 13812 20168 13864
rect 20220 13852 20226 13864
rect 20257 13855 20315 13861
rect 20257 13852 20269 13855
rect 20220 13824 20269 13852
rect 20220 13812 20226 13824
rect 20257 13821 20269 13824
rect 20303 13852 20315 13855
rect 20916 13852 20944 13883
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 20303 13824 20944 13852
rect 22204 13852 22232 13960
rect 22281 13957 22293 13991
rect 22327 13988 22339 13991
rect 22370 13988 22376 14000
rect 22327 13960 22376 13988
rect 22327 13957 22339 13960
rect 22281 13951 22339 13957
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 23492 13929 23520 14028
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 23934 14056 23940 14068
rect 23895 14028 23940 14056
rect 23934 14016 23940 14028
rect 23992 14016 23998 14068
rect 24949 14059 25007 14065
rect 24949 14025 24961 14059
rect 24995 14056 25007 14059
rect 25130 14056 25136 14068
rect 24995 14028 25136 14056
rect 24995 14025 25007 14028
rect 24949 14019 25007 14025
rect 24397 13991 24455 13997
rect 24397 13957 24409 13991
rect 24443 13988 24455 13991
rect 24964 13988 24992 14019
rect 25130 14016 25136 14028
rect 25188 14016 25194 14068
rect 27246 14056 27252 14068
rect 27207 14028 27252 14056
rect 27246 14016 27252 14028
rect 27304 14016 27310 14068
rect 29822 14016 29828 14068
rect 29880 14016 29886 14068
rect 31389 14059 31447 14065
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 31478 14056 31484 14068
rect 31435 14028 31484 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 26326 13988 26332 14000
rect 24443 13960 24992 13988
rect 26160 13960 26332 13988
rect 24443 13957 24455 13960
rect 24397 13951 24455 13957
rect 23201 13923 23259 13929
rect 23201 13889 23213 13923
rect 23247 13920 23259 13923
rect 23477 13923 23535 13929
rect 23247 13892 23428 13920
rect 23247 13889 23259 13892
rect 23201 13883 23259 13889
rect 23290 13852 23296 13864
rect 22204 13824 23152 13852
rect 23251 13824 23296 13852
rect 20303 13821 20315 13824
rect 20257 13815 20315 13821
rect 20717 13787 20775 13793
rect 20717 13784 20729 13787
rect 19812 13756 20729 13784
rect 20717 13753 20729 13756
rect 20763 13753 20775 13787
rect 23124 13784 23152 13824
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 23400 13852 23428 13892
rect 23477 13889 23489 13923
rect 23523 13889 23535 13923
rect 24026 13920 24032 13932
rect 23477 13883 23535 13889
rect 23584 13892 24032 13920
rect 23584 13852 23612 13892
rect 24026 13880 24032 13892
rect 24084 13880 24090 13932
rect 24118 13880 24124 13932
rect 24176 13920 24182 13932
rect 24176 13892 24221 13920
rect 24176 13880 24182 13892
rect 23400 13824 23612 13852
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 24213 13855 24271 13861
rect 24213 13852 24225 13855
rect 23716 13824 24225 13852
rect 23716 13812 23722 13824
rect 24213 13821 24225 13824
rect 24259 13821 24271 13855
rect 26160 13852 26188 13960
rect 26326 13948 26332 13960
rect 26384 13948 26390 14000
rect 28626 13988 28632 14000
rect 28587 13960 28632 13988
rect 28626 13948 28632 13960
rect 28684 13948 28690 14000
rect 28810 13988 28816 14000
rect 28771 13960 28816 13988
rect 28810 13948 28816 13960
rect 28868 13948 28874 14000
rect 28997 13991 29055 13997
rect 28997 13957 29009 13991
rect 29043 13988 29055 13991
rect 29043 13960 29592 13988
rect 29043 13957 29055 13960
rect 28997 13951 29055 13957
rect 26418 13920 26424 13932
rect 26331 13892 26424 13920
rect 26418 13880 26424 13892
rect 26476 13920 26482 13932
rect 27709 13929 27767 13935
rect 27479 13923 27537 13929
rect 27479 13920 27491 13923
rect 26476 13892 27491 13920
rect 26476 13880 26482 13892
rect 27479 13889 27491 13892
rect 27525 13889 27537 13923
rect 27479 13883 27537 13889
rect 27598 13923 27656 13929
rect 27598 13889 27610 13923
rect 27644 13920 27656 13923
rect 27644 13889 27657 13920
rect 27709 13895 27721 13929
rect 27755 13920 27767 13929
rect 27798 13920 27804 13932
rect 27755 13895 27804 13920
rect 27709 13892 27804 13895
rect 27709 13889 27767 13892
rect 27598 13883 27657 13889
rect 27629 13852 27657 13883
rect 27798 13880 27804 13892
rect 27856 13880 27862 13932
rect 27893 13923 27951 13929
rect 27893 13889 27905 13923
rect 27939 13920 27951 13923
rect 28074 13920 28080 13932
rect 27939 13892 28080 13920
rect 27939 13889 27951 13892
rect 27893 13883 27951 13889
rect 28074 13880 28080 13892
rect 28132 13880 28138 13932
rect 29454 13920 29460 13932
rect 29415 13892 29460 13920
rect 29454 13880 29460 13892
rect 29512 13880 29518 13932
rect 29564 13926 29592 13960
rect 29620 13929 29678 13935
rect 29840 13929 29868 14016
rect 30650 13988 30656 14000
rect 30563 13960 30656 13988
rect 30650 13948 30656 13960
rect 30708 13988 30714 14000
rect 31404 13988 31432 14019
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 35986 14016 35992 14068
rect 36044 14056 36050 14068
rect 39758 14056 39764 14068
rect 36044 14028 38976 14056
rect 39719 14028 39764 14056
rect 36044 14016 36050 14028
rect 30708 13960 31432 13988
rect 35529 13991 35587 13997
rect 30708 13948 30714 13960
rect 35529 13957 35541 13991
rect 35575 13988 35587 13991
rect 37182 13988 37188 14000
rect 35575 13960 37188 13988
rect 35575 13957 35587 13960
rect 35529 13951 35587 13957
rect 37182 13948 37188 13960
rect 37240 13948 37246 14000
rect 37642 13948 37648 14000
rect 37700 13988 37706 14000
rect 38948 13988 38976 14028
rect 39758 14016 39764 14028
rect 39816 14016 39822 14068
rect 39853 13991 39911 13997
rect 39853 13988 39865 13991
rect 37700 13960 38884 13988
rect 38948 13960 39865 13988
rect 37700 13948 37706 13960
rect 29620 13926 29632 13929
rect 29564 13898 29632 13926
rect 29620 13895 29632 13898
rect 29666 13895 29678 13929
rect 29620 13889 29678 13895
rect 29733 13923 29791 13929
rect 29733 13889 29745 13923
rect 29779 13889 29791 13923
rect 29733 13883 29791 13889
rect 29825 13923 29883 13929
rect 29825 13889 29837 13923
rect 29871 13889 29883 13923
rect 29825 13883 29883 13889
rect 30837 13923 30895 13929
rect 30837 13889 30849 13923
rect 30883 13920 30895 13923
rect 31294 13920 31300 13932
rect 30883 13892 31300 13920
rect 30883 13889 30895 13892
rect 30837 13883 30895 13889
rect 29748 13852 29776 13883
rect 31294 13880 31300 13892
rect 31352 13880 31358 13932
rect 33134 13880 33140 13932
rect 33192 13920 33198 13932
rect 34434 13923 34492 13929
rect 34434 13920 34446 13923
rect 33192 13892 34446 13920
rect 33192 13880 33198 13892
rect 34434 13889 34446 13892
rect 34480 13889 34492 13923
rect 34434 13883 34492 13889
rect 34606 13880 34612 13932
rect 34664 13920 34670 13932
rect 34701 13923 34759 13929
rect 34701 13920 34713 13923
rect 34664 13892 34713 13920
rect 34664 13880 34670 13892
rect 34701 13889 34713 13892
rect 34747 13889 34759 13923
rect 35158 13920 35164 13932
rect 35119 13892 35164 13920
rect 34701 13883 34759 13889
rect 35158 13880 35164 13892
rect 35216 13880 35222 13932
rect 35345 13923 35403 13929
rect 35345 13889 35357 13923
rect 35391 13920 35403 13923
rect 35434 13920 35440 13932
rect 35391 13892 35440 13920
rect 35391 13889 35403 13892
rect 35345 13883 35403 13889
rect 35434 13880 35440 13892
rect 35492 13880 35498 13932
rect 36265 13923 36323 13929
rect 36265 13889 36277 13923
rect 36311 13889 36323 13923
rect 36265 13883 36323 13889
rect 38565 13923 38623 13929
rect 38565 13889 38577 13923
rect 38611 13889 38623 13923
rect 38746 13920 38752 13932
rect 38707 13892 38752 13920
rect 38565 13883 38623 13889
rect 29914 13852 29920 13864
rect 24213 13815 24271 13821
rect 24320 13824 26188 13852
rect 27448 13824 29920 13852
rect 24320 13784 24348 13824
rect 27448 13796 27476 13824
rect 29914 13812 29920 13824
rect 29972 13812 29978 13864
rect 30101 13855 30159 13861
rect 30101 13821 30113 13855
rect 30147 13852 30159 13855
rect 30558 13852 30564 13864
rect 30147 13824 30564 13852
rect 30147 13821 30159 13824
rect 30101 13815 30159 13821
rect 30558 13812 30564 13824
rect 30616 13812 30622 13864
rect 35176 13852 35204 13880
rect 35894 13852 35900 13864
rect 35176 13824 35900 13852
rect 35894 13812 35900 13824
rect 35952 13852 35958 13864
rect 36081 13855 36139 13861
rect 36081 13852 36093 13855
rect 35952 13824 36093 13852
rect 35952 13812 35958 13824
rect 36081 13821 36093 13824
rect 36127 13821 36139 13855
rect 36081 13815 36139 13821
rect 23124 13756 24348 13784
rect 20717 13747 20775 13753
rect 27430 13744 27436 13796
rect 27488 13744 27494 13796
rect 35342 13744 35348 13796
rect 35400 13784 35406 13796
rect 36280 13784 36308 13883
rect 37274 13852 37280 13864
rect 37235 13824 37280 13852
rect 37274 13812 37280 13824
rect 37332 13812 37338 13864
rect 37550 13852 37556 13864
rect 37511 13824 37556 13852
rect 37550 13812 37556 13824
rect 37608 13812 37614 13864
rect 38580 13852 38608 13883
rect 38746 13880 38752 13892
rect 38804 13880 38810 13932
rect 38856 13929 38884 13960
rect 39853 13957 39865 13960
rect 39899 13988 39911 13991
rect 40678 13988 40684 14000
rect 39899 13960 40684 13988
rect 39899 13957 39911 13960
rect 39853 13951 39911 13957
rect 40678 13948 40684 13960
rect 40736 13948 40742 14000
rect 38841 13923 38899 13929
rect 38841 13889 38853 13923
rect 38887 13889 38899 13923
rect 38841 13883 38899 13889
rect 38930 13880 38936 13932
rect 38988 13920 38994 13932
rect 38988 13892 39033 13920
rect 38988 13880 38994 13892
rect 39758 13852 39764 13864
rect 38580 13824 39764 13852
rect 39758 13812 39764 13824
rect 39816 13812 39822 13864
rect 35400 13756 36308 13784
rect 35400 13744 35406 13756
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 7006 13716 7012 13728
rect 4948 13688 7012 13716
rect 4948 13676 4954 13688
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 14645 13719 14703 13725
rect 14645 13685 14657 13719
rect 14691 13716 14703 13719
rect 15010 13716 15016 13728
rect 14691 13688 15016 13716
rect 14691 13685 14703 13688
rect 14645 13679 14703 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 21818 13716 21824 13728
rect 19208 13688 21824 13716
rect 19208 13676 19214 13688
rect 21818 13676 21824 13688
rect 21876 13676 21882 13728
rect 23106 13676 23112 13728
rect 23164 13716 23170 13728
rect 23201 13719 23259 13725
rect 23201 13716 23213 13719
rect 23164 13688 23213 13716
rect 23164 13676 23170 13688
rect 23201 13685 23213 13688
rect 23247 13685 23259 13719
rect 23201 13679 23259 13685
rect 23474 13676 23480 13728
rect 23532 13716 23538 13728
rect 24121 13719 24179 13725
rect 24121 13716 24133 13719
rect 23532 13688 24133 13716
rect 23532 13676 23538 13688
rect 24121 13685 24133 13688
rect 24167 13685 24179 13719
rect 33318 13716 33324 13728
rect 33279 13688 33324 13716
rect 24121 13679 24179 13685
rect 33318 13676 33324 13688
rect 33376 13676 33382 13728
rect 36449 13719 36507 13725
rect 36449 13685 36461 13719
rect 36495 13716 36507 13719
rect 37734 13716 37740 13728
rect 36495 13688 37740 13716
rect 36495 13685 36507 13688
rect 36449 13679 36507 13685
rect 37734 13676 37740 13688
rect 37792 13676 37798 13728
rect 39206 13716 39212 13728
rect 39167 13688 39212 13716
rect 39206 13676 39212 13688
rect 39264 13676 39270 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 5166 13512 5172 13524
rect 5127 13484 5172 13512
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 11977 13515 12035 13521
rect 11977 13481 11989 13515
rect 12023 13512 12035 13515
rect 12250 13512 12256 13524
rect 12023 13484 12256 13512
rect 12023 13481 12035 13484
rect 11977 13475 12035 13481
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 14461 13515 14519 13521
rect 14461 13481 14473 13515
rect 14507 13512 14519 13515
rect 15194 13512 15200 13524
rect 14507 13484 15200 13512
rect 14507 13481 14519 13484
rect 14461 13475 14519 13481
rect 15194 13472 15200 13484
rect 15252 13472 15258 13524
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 21269 13515 21327 13521
rect 21269 13512 21281 13515
rect 21232 13484 21281 13512
rect 21232 13472 21238 13484
rect 21269 13481 21281 13484
rect 21315 13481 21327 13515
rect 22186 13512 22192 13524
rect 22147 13484 22192 13512
rect 21269 13475 21327 13481
rect 22186 13472 22192 13484
rect 22244 13472 22250 13524
rect 27062 13512 27068 13524
rect 27023 13484 27068 13512
rect 27062 13472 27068 13484
rect 27120 13472 27126 13524
rect 27706 13472 27712 13524
rect 27764 13512 27770 13524
rect 28169 13515 28227 13521
rect 28169 13512 28181 13515
rect 27764 13484 28181 13512
rect 27764 13472 27770 13484
rect 28169 13481 28181 13484
rect 28215 13481 28227 13515
rect 28169 13475 28227 13481
rect 28810 13472 28816 13524
rect 28868 13512 28874 13524
rect 29549 13515 29607 13521
rect 29549 13512 29561 13515
rect 28868 13484 29561 13512
rect 28868 13472 28874 13484
rect 29549 13481 29561 13484
rect 29595 13481 29607 13515
rect 29549 13475 29607 13481
rect 31294 13472 31300 13524
rect 31352 13512 31358 13524
rect 33134 13512 33140 13524
rect 31352 13484 32076 13512
rect 33095 13484 33140 13512
rect 31352 13472 31358 13484
rect 14826 13404 14832 13456
rect 14884 13444 14890 13456
rect 17954 13444 17960 13456
rect 14884 13416 17960 13444
rect 14884 13404 14890 13416
rect 17954 13404 17960 13416
rect 18012 13444 18018 13456
rect 18601 13447 18659 13453
rect 18601 13444 18613 13447
rect 18012 13416 18613 13444
rect 18012 13404 18018 13416
rect 18601 13413 18613 13416
rect 18647 13413 18659 13447
rect 18601 13407 18659 13413
rect 20809 13447 20867 13453
rect 20809 13413 20821 13447
rect 20855 13444 20867 13447
rect 20898 13444 20904 13456
rect 20855 13416 20904 13444
rect 20855 13413 20867 13416
rect 20809 13407 20867 13413
rect 2501 13379 2559 13385
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2774 13376 2780 13388
rect 2547 13348 2780 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 5626 13376 5632 13388
rect 5587 13348 5632 13376
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 5813 13379 5871 13385
rect 5813 13345 5825 13379
rect 5859 13376 5871 13379
rect 6178 13376 6184 13388
rect 5859 13348 6184 13376
rect 5859 13345 5871 13348
rect 5813 13339 5871 13345
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8938 13376 8944 13388
rect 8899 13348 8944 13376
rect 8938 13336 8944 13348
rect 8996 13336 9002 13388
rect 14568 13348 14872 13376
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 6604 13280 6653 13308
rect 6604 13268 6610 13280
rect 6641 13277 6653 13280
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8386 13308 8392 13320
rect 8260 13280 8392 13308
rect 8260 13268 8266 13280
rect 8386 13268 8392 13280
rect 8444 13308 8450 13320
rect 9217 13311 9275 13317
rect 9217 13308 9229 13311
rect 8444 13280 9229 13308
rect 8444 13268 8450 13280
rect 9217 13277 9229 13280
rect 9263 13308 9275 13311
rect 10042 13308 10048 13320
rect 9263 13280 10048 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 11480 13280 11805 13308
rect 11480 13268 11486 13280
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 2038 13132 2044 13184
rect 2096 13172 2102 13184
rect 2133 13175 2191 13181
rect 2133 13172 2145 13175
rect 2096 13144 2145 13172
rect 2096 13132 2102 13144
rect 2133 13141 2145 13144
rect 2179 13141 2191 13175
rect 4614 13172 4620 13184
rect 4575 13144 4620 13172
rect 2133 13135 2191 13141
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 5534 13172 5540 13184
rect 5495 13144 5540 13172
rect 5534 13132 5540 13144
rect 5592 13132 5598 13184
rect 14568 13172 14596 13348
rect 14734 13308 14740 13320
rect 14695 13280 14740 13308
rect 14734 13268 14740 13280
rect 14792 13268 14798 13320
rect 14844 13317 14872 13348
rect 15010 13336 15016 13388
rect 15068 13336 15074 13388
rect 14826 13311 14884 13317
rect 14826 13277 14838 13311
rect 14872 13277 14884 13311
rect 14826 13271 14884 13277
rect 14921 13305 14979 13311
rect 14921 13271 14933 13305
rect 14967 13302 14979 13305
rect 15028 13302 15056 13336
rect 14967 13274 15056 13302
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15378 13308 15384 13320
rect 15151 13280 15384 13308
rect 15151 13277 15163 13280
rect 14967 13271 14979 13274
rect 15105 13271 15163 13277
rect 14921 13265 14979 13271
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15654 13268 15660 13320
rect 15712 13308 15718 13320
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 15712 13280 17693 13308
rect 15712 13268 15718 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 15562 13240 15568 13252
rect 15523 13212 15568 13240
rect 15562 13200 15568 13212
rect 15620 13200 15626 13252
rect 17494 13240 17500 13252
rect 17455 13212 17500 13240
rect 17494 13200 17500 13212
rect 17552 13200 17558 13252
rect 18616 13240 18644 13407
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 27724 13444 27752 13472
rect 24780 13416 27752 13444
rect 23842 13376 23848 13388
rect 23803 13348 23848 13376
rect 23842 13336 23848 13348
rect 23900 13336 23906 13388
rect 19337 13311 19395 13317
rect 19337 13277 19349 13311
rect 19383 13308 19395 13311
rect 19426 13308 19432 13320
rect 19383 13280 19432 13308
rect 19383 13277 19395 13280
rect 19337 13271 19395 13277
rect 19426 13268 19432 13280
rect 19484 13308 19490 13320
rect 24780 13317 24808 13416
rect 26234 13336 26240 13388
rect 26292 13376 26298 13388
rect 26510 13376 26516 13388
rect 26292 13348 26516 13376
rect 26292 13336 26298 13348
rect 26510 13336 26516 13348
rect 26568 13336 26574 13388
rect 30929 13379 30987 13385
rect 30929 13345 30941 13379
rect 30975 13376 30987 13379
rect 31754 13376 31760 13388
rect 30975 13348 31760 13376
rect 30975 13345 30987 13348
rect 30929 13339 30987 13345
rect 31754 13336 31760 13348
rect 31812 13336 31818 13388
rect 32048 13385 32076 13484
rect 33134 13472 33140 13484
rect 33192 13472 33198 13524
rect 35894 13472 35900 13524
rect 35952 13512 35958 13524
rect 37277 13515 37335 13521
rect 37277 13512 37289 13515
rect 35952 13484 37289 13512
rect 35952 13472 35958 13484
rect 37277 13481 37289 13484
rect 37323 13481 37335 13515
rect 37277 13475 37335 13481
rect 38197 13515 38255 13521
rect 38197 13481 38209 13515
rect 38243 13512 38255 13515
rect 38746 13512 38752 13524
rect 38243 13484 38752 13512
rect 38243 13481 38255 13484
rect 38197 13475 38255 13481
rect 38746 13472 38752 13484
rect 38804 13472 38810 13524
rect 32033 13379 32091 13385
rect 32033 13345 32045 13379
rect 32079 13376 32091 13379
rect 32079 13348 32904 13376
rect 32079 13345 32091 13348
rect 32033 13339 32091 13345
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 19484 13280 20637 13308
rect 19484 13268 19490 13280
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 20625 13271 20683 13277
rect 23569 13311 23627 13317
rect 23569 13277 23581 13311
rect 23615 13277 23627 13311
rect 23569 13271 23627 13277
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 19889 13243 19947 13249
rect 19889 13240 19901 13243
rect 18616 13212 19901 13240
rect 19889 13209 19901 13212
rect 19935 13209 19947 13243
rect 19889 13203 19947 13209
rect 20073 13243 20131 13249
rect 20073 13209 20085 13243
rect 20119 13240 20131 13243
rect 20714 13240 20720 13252
rect 20119 13212 20720 13240
rect 20119 13209 20131 13212
rect 20073 13203 20131 13209
rect 20714 13200 20720 13212
rect 20772 13200 20778 13252
rect 23584 13240 23612 13271
rect 27246 13268 27252 13320
rect 27304 13317 27310 13320
rect 27304 13311 27353 13317
rect 27304 13277 27307 13311
rect 27341 13277 27353 13311
rect 27430 13308 27436 13320
rect 27391 13280 27436 13308
rect 27304 13271 27353 13277
rect 27304 13268 27310 13271
rect 27430 13268 27436 13280
rect 27488 13268 27494 13320
rect 27522 13268 27528 13320
rect 27580 13308 27586 13320
rect 27709 13311 27767 13317
rect 27580 13280 27625 13308
rect 27580 13268 27586 13280
rect 27709 13277 27721 13311
rect 27755 13308 27767 13311
rect 28074 13308 28080 13320
rect 27755 13280 28080 13308
rect 27755 13277 27767 13280
rect 27709 13271 27767 13277
rect 28074 13268 28080 13280
rect 28132 13268 28138 13320
rect 32490 13308 32496 13320
rect 32451 13280 32496 13308
rect 32490 13268 32496 13280
rect 32548 13268 32554 13320
rect 32674 13308 32680 13320
rect 32635 13280 32680 13308
rect 32674 13268 32680 13280
rect 32732 13268 32738 13320
rect 32876 13317 32904 13348
rect 35342 13336 35348 13388
rect 35400 13376 35406 13388
rect 35400 13348 36584 13376
rect 35400 13336 35406 13348
rect 32769 13311 32827 13317
rect 32769 13277 32781 13311
rect 32815 13277 32827 13311
rect 32769 13271 32827 13277
rect 32861 13311 32919 13317
rect 32861 13277 32873 13311
rect 32907 13277 32919 13311
rect 35710 13308 35716 13320
rect 35671 13280 35716 13308
rect 32861 13271 32919 13277
rect 25222 13240 25228 13252
rect 23584 13212 25228 13240
rect 25222 13200 25228 13212
rect 25280 13200 25286 13252
rect 30558 13200 30564 13252
rect 30616 13240 30622 13252
rect 30662 13243 30720 13249
rect 30662 13240 30674 13243
rect 30616 13212 30674 13240
rect 30616 13200 30622 13212
rect 30662 13209 30674 13212
rect 30708 13209 30720 13243
rect 30662 13203 30720 13209
rect 31018 13200 31024 13252
rect 31076 13240 31082 13252
rect 32784 13240 32812 13271
rect 35710 13268 35716 13280
rect 35768 13268 35774 13320
rect 35986 13308 35992 13320
rect 35947 13280 35992 13308
rect 35986 13268 35992 13280
rect 36044 13268 36050 13320
rect 36556 13317 36584 13348
rect 36541 13311 36599 13317
rect 36541 13277 36553 13311
rect 36587 13277 36599 13311
rect 36722 13308 36728 13320
rect 36683 13280 36728 13308
rect 36541 13271 36599 13277
rect 36722 13268 36728 13280
rect 36780 13268 36786 13320
rect 38010 13308 38016 13320
rect 37971 13280 38016 13308
rect 38010 13268 38016 13280
rect 38068 13268 38074 13320
rect 58158 13308 58164 13320
rect 58119 13280 58164 13308
rect 58158 13268 58164 13280
rect 58216 13268 58222 13320
rect 34698 13240 34704 13252
rect 31076 13212 32812 13240
rect 33244 13212 34704 13240
rect 31076 13200 31082 13212
rect 15286 13172 15292 13184
rect 14568 13144 15292 13172
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 17865 13175 17923 13181
rect 17865 13141 17877 13175
rect 17911 13172 17923 13175
rect 19150 13172 19156 13184
rect 17911 13144 19156 13172
rect 17911 13141 17923 13144
rect 17865 13135 17923 13141
rect 19150 13132 19156 13144
rect 19208 13132 19214 13184
rect 24394 13132 24400 13184
rect 24452 13172 24458 13184
rect 33244 13172 33272 13212
rect 34698 13200 34704 13212
rect 34756 13200 34762 13252
rect 37274 13200 37280 13252
rect 37332 13240 37338 13252
rect 37550 13240 37556 13252
rect 37332 13212 37556 13240
rect 37332 13200 37338 13212
rect 37550 13200 37556 13212
rect 37608 13240 37614 13252
rect 37829 13243 37887 13249
rect 37829 13240 37841 13243
rect 37608 13212 37841 13240
rect 37608 13200 37614 13212
rect 37829 13209 37841 13212
rect 37875 13209 37887 13243
rect 37829 13203 37887 13209
rect 33594 13172 33600 13184
rect 24452 13144 33272 13172
rect 33555 13144 33600 13172
rect 24452 13132 24458 13144
rect 33594 13132 33600 13144
rect 33652 13132 33658 13184
rect 36354 13132 36360 13184
rect 36412 13172 36418 13184
rect 36725 13175 36783 13181
rect 36725 13172 36737 13175
rect 36412 13144 36737 13172
rect 36412 13132 36418 13144
rect 36725 13141 36737 13144
rect 36771 13172 36783 13175
rect 39482 13172 39488 13184
rect 36771 13144 39488 13172
rect 36771 13141 36783 13144
rect 36725 13135 36783 13141
rect 39482 13132 39488 13144
rect 39540 13172 39546 13184
rect 39942 13172 39948 13184
rect 39540 13144 39948 13172
rect 39540 13132 39546 13144
rect 39942 13132 39948 13144
rect 40000 13132 40006 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 2372 12940 4813 12968
rect 2372 12928 2378 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 4801 12931 4859 12937
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 5592 12940 6469 12968
rect 5592 12928 5598 12940
rect 6457 12937 6469 12940
rect 6503 12968 6515 12971
rect 9398 12968 9404 12980
rect 6503 12940 9404 12968
rect 6503 12937 6515 12940
rect 6457 12931 6515 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10597 12971 10655 12977
rect 10597 12937 10609 12971
rect 10643 12968 10655 12971
rect 10870 12968 10876 12980
rect 10643 12940 10876 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 3786 12900 3792 12912
rect 2700 12872 3792 12900
rect 2038 12832 2044 12844
rect 1999 12804 2044 12832
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2700 12841 2728 12872
rect 3786 12860 3792 12872
rect 3844 12900 3850 12912
rect 9674 12900 9680 12912
rect 3844 12872 8340 12900
rect 3844 12860 3850 12872
rect 8312 12844 8340 12872
rect 9508 12872 9680 12900
rect 2685 12835 2743 12841
rect 2685 12801 2697 12835
rect 2731 12801 2743 12835
rect 2941 12835 2999 12841
rect 2941 12832 2953 12835
rect 2685 12795 2743 12801
rect 2792 12804 2953 12832
rect 2792 12764 2820 12804
rect 2941 12801 2953 12804
rect 2987 12801 2999 12835
rect 2941 12795 2999 12801
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 5169 12835 5227 12841
rect 5169 12832 5181 12835
rect 4672 12804 5181 12832
rect 4672 12792 4678 12804
rect 5169 12801 5181 12804
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 6730 12832 6736 12844
rect 5307 12804 6736 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 2240 12736 2820 12764
rect 2240 12705 2268 12736
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 5408 12736 5453 12764
rect 5408 12724 5414 12736
rect 2225 12699 2283 12705
rect 2225 12665 2237 12699
rect 2271 12665 2283 12699
rect 2225 12659 2283 12665
rect 4065 12699 4123 12705
rect 4065 12665 4077 12699
rect 4111 12696 4123 12699
rect 5552 12696 5580 12804
rect 6730 12792 6736 12804
rect 6788 12792 6794 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 8122 12835 8180 12841
rect 8122 12832 8134 12835
rect 7616 12804 8134 12832
rect 7616 12792 7622 12804
rect 8122 12801 8134 12804
rect 8168 12801 8180 12835
rect 8122 12795 8180 12801
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 9508 12841 9536 12872
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 9766 12860 9772 12912
rect 9824 12860 9830 12912
rect 10612 12900 10640 12931
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 21818 12968 21824 12980
rect 14936 12940 15240 12968
rect 21779 12940 21824 12968
rect 13906 12900 13912 12912
rect 9968 12872 10640 12900
rect 13867 12872 13912 12900
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8352 12804 8401 12832
rect 8352 12792 8358 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9784 12832 9812 12860
rect 9493 12795 9551 12801
rect 9600 12804 9812 12832
rect 9861 12835 9919 12841
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 9600 12764 9628 12804
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 9968 12832 9996 12872
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 14090 12900 14096 12912
rect 14051 12872 14096 12900
rect 14090 12860 14096 12872
rect 14148 12860 14154 12912
rect 14277 12903 14335 12909
rect 14277 12869 14289 12903
rect 14323 12900 14335 12903
rect 14936 12900 14964 12940
rect 14323 12872 14964 12900
rect 14323 12869 14335 12872
rect 14277 12863 14335 12869
rect 9907 12804 9996 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 11698 12832 11704 12844
rect 10100 12804 10145 12832
rect 11659 12804 11704 12832
rect 10100 12792 10106 12804
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12066 12832 12072 12844
rect 12027 12804 12072 12832
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 15212 12841 15240 12940
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 23569 12971 23627 12977
rect 23569 12937 23581 12971
rect 23615 12968 23627 12971
rect 23842 12968 23848 12980
rect 23615 12940 23848 12968
rect 23615 12937 23627 12940
rect 23569 12931 23627 12937
rect 23842 12928 23848 12940
rect 23900 12928 23906 12980
rect 24026 12928 24032 12980
rect 24084 12968 24090 12980
rect 24121 12971 24179 12977
rect 24121 12968 24133 12971
rect 24084 12940 24133 12968
rect 24084 12928 24090 12940
rect 24121 12937 24133 12940
rect 24167 12968 24179 12971
rect 24210 12968 24216 12980
rect 24167 12940 24216 12968
rect 24167 12937 24179 12940
rect 24121 12931 24179 12937
rect 24210 12928 24216 12940
rect 24268 12928 24274 12980
rect 32674 12968 32680 12980
rect 32635 12940 32680 12968
rect 32674 12928 32680 12940
rect 32732 12928 32738 12980
rect 35069 12971 35127 12977
rect 35069 12937 35081 12971
rect 35115 12968 35127 12971
rect 35894 12968 35900 12980
rect 35115 12940 35900 12968
rect 35115 12937 35127 12940
rect 35069 12931 35127 12937
rect 35894 12928 35900 12940
rect 35952 12928 35958 12980
rect 36722 12968 36728 12980
rect 36004 12940 36728 12968
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 16816 12872 18184 12900
rect 16816 12860 16822 12872
rect 12253 12835 12311 12841
rect 15013 12835 15071 12841
rect 12253 12801 12265 12835
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 14853 12807 15025 12835
rect 9355 12736 9628 12764
rect 9677 12767 9735 12773
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 9677 12733 9689 12767
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 9769 12767 9827 12773
rect 9769 12733 9781 12767
rect 9815 12764 9827 12767
rect 11882 12764 11888 12776
rect 9815 12736 9904 12764
rect 9815 12733 9827 12736
rect 9769 12727 9827 12733
rect 4111 12668 5580 12696
rect 4111 12665 4123 12668
rect 4065 12659 4123 12665
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 9692 12696 9720 12727
rect 9876 12708 9904 12736
rect 9968 12736 11888 12764
rect 9640 12668 9812 12696
rect 9640 12656 9646 12668
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 9784 12628 9812 12668
rect 9858 12656 9864 12708
rect 9916 12656 9922 12708
rect 9968 12628 9996 12736
rect 11882 12724 11888 12736
rect 11940 12724 11946 12776
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12032 12736 12077 12764
rect 12032 12724 12038 12736
rect 10042 12656 10048 12708
rect 10100 12696 10106 12708
rect 12268 12696 12296 12795
rect 10100 12668 12296 12696
rect 14853 12696 14881 12807
rect 15013 12801 15025 12807
rect 15059 12801 15071 12835
rect 15013 12795 15071 12801
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12801 15255 12835
rect 15197 12795 15255 12801
rect 15120 12764 15148 12795
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 18156 12841 18184 12872
rect 23106 12860 23112 12912
rect 23164 12900 23170 12912
rect 23750 12900 23756 12912
rect 23164 12872 23756 12900
rect 23164 12860 23170 12872
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 23860 12900 23888 12928
rect 24673 12903 24731 12909
rect 24673 12900 24685 12903
rect 23860 12872 24685 12900
rect 24673 12869 24685 12872
rect 24719 12869 24731 12903
rect 24673 12863 24731 12869
rect 32493 12903 32551 12909
rect 32493 12869 32505 12903
rect 32539 12900 32551 12903
rect 33134 12900 33140 12912
rect 32539 12872 33140 12900
rect 32539 12869 32551 12872
rect 32493 12863 32551 12869
rect 33134 12860 33140 12872
rect 33192 12900 33198 12912
rect 33318 12900 33324 12912
rect 33192 12872 33324 12900
rect 33192 12860 33198 12872
rect 33318 12860 33324 12872
rect 33376 12860 33382 12912
rect 35621 12903 35679 12909
rect 35621 12869 35633 12903
rect 35667 12900 35679 12903
rect 36004 12900 36032 12940
rect 36722 12928 36728 12940
rect 36780 12928 36786 12980
rect 38010 12928 38016 12980
rect 38068 12968 38074 12980
rect 40037 12971 40095 12977
rect 40037 12968 40049 12971
rect 38068 12940 40049 12968
rect 38068 12928 38074 12940
rect 40037 12937 40049 12940
rect 40083 12937 40095 12971
rect 40037 12931 40095 12937
rect 35667 12872 36032 12900
rect 35667 12869 35679 12872
rect 35621 12863 35679 12869
rect 37366 12860 37372 12912
rect 37424 12900 37430 12912
rect 37461 12903 37519 12909
rect 37461 12900 37473 12903
rect 37424 12872 37473 12900
rect 37424 12860 37430 12872
rect 37461 12869 37473 12872
rect 37507 12869 37519 12903
rect 37461 12863 37519 12869
rect 37645 12903 37703 12909
rect 37645 12869 37657 12903
rect 37691 12900 37703 12903
rect 37734 12900 37740 12912
rect 37691 12872 37740 12900
rect 37691 12869 37703 12872
rect 37645 12863 37703 12869
rect 37734 12860 37740 12872
rect 37792 12860 37798 12912
rect 38924 12903 38982 12909
rect 38924 12869 38936 12903
rect 38970 12900 38982 12903
rect 39206 12900 39212 12912
rect 38970 12872 39212 12900
rect 38970 12869 38982 12872
rect 38924 12863 38982 12869
rect 39206 12860 39212 12872
rect 39264 12860 39270 12912
rect 17885 12835 17943 12841
rect 15436 12804 16804 12832
rect 15436 12792 15442 12804
rect 16776 12776 16804 12804
rect 17885 12801 17897 12835
rect 17931 12832 17943 12835
rect 18141 12835 18199 12841
rect 17931 12804 18092 12832
rect 17931 12801 17943 12804
rect 17885 12795 17943 12801
rect 15286 12764 15292 12776
rect 15120 12736 15292 12764
rect 15286 12724 15292 12736
rect 15344 12764 15350 12776
rect 16114 12764 16120 12776
rect 15344 12736 16120 12764
rect 15344 12724 15350 12736
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 16758 12724 16764 12776
rect 16816 12724 16822 12776
rect 18064 12764 18092 12804
rect 18141 12801 18153 12835
rect 18187 12801 18199 12835
rect 18141 12795 18199 12801
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 18966 12835 19024 12841
rect 18966 12801 18978 12835
rect 19012 12801 19024 12835
rect 18966 12795 19024 12801
rect 19061 12835 19119 12841
rect 19061 12801 19073 12835
rect 19107 12832 19119 12835
rect 19150 12832 19156 12844
rect 19107 12804 19156 12832
rect 19107 12801 19119 12804
rect 19061 12795 19119 12801
rect 18601 12767 18659 12773
rect 18601 12764 18613 12767
rect 18064 12736 18613 12764
rect 18601 12733 18613 12736
rect 18647 12733 18659 12767
rect 18601 12727 18659 12733
rect 15746 12696 15752 12708
rect 14853 12668 15752 12696
rect 10100 12656 10106 12668
rect 15746 12656 15752 12668
rect 15804 12696 15810 12708
rect 15841 12699 15899 12705
rect 15841 12696 15853 12699
rect 15804 12668 15853 12696
rect 15804 12656 15810 12668
rect 15841 12665 15853 12668
rect 15887 12665 15899 12699
rect 15841 12659 15899 12665
rect 9784 12600 9996 12628
rect 11517 12631 11575 12637
rect 11517 12597 11529 12631
rect 11563 12628 11575 12631
rect 11606 12628 11612 12640
rect 11563 12600 11612 12628
rect 11563 12597 11575 12600
rect 11517 12591 11575 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 14737 12631 14795 12637
rect 14737 12597 14749 12631
rect 14783 12628 14795 12631
rect 15194 12628 15200 12640
rect 14783 12600 15200 12628
rect 14783 12597 14795 12600
rect 14737 12591 14795 12597
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 16761 12631 16819 12637
rect 16761 12628 16773 12631
rect 15712 12600 16773 12628
rect 15712 12588 15718 12600
rect 16761 12597 16773 12600
rect 16807 12597 16819 12631
rect 18892 12628 18920 12795
rect 18981 12708 19009 12795
rect 19150 12792 19156 12804
rect 19208 12792 19214 12844
rect 19242 12792 19248 12844
rect 19300 12832 19306 12844
rect 20990 12832 20996 12844
rect 19300 12804 19345 12832
rect 20951 12804 20996 12832
rect 19300 12792 19306 12804
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 22922 12832 22928 12844
rect 22835 12804 22928 12832
rect 22922 12792 22928 12804
rect 22980 12832 22986 12844
rect 23477 12835 23535 12841
rect 23477 12832 23489 12835
rect 22980 12804 23489 12832
rect 22980 12792 22986 12804
rect 23477 12801 23489 12804
rect 23523 12801 23535 12835
rect 23477 12795 23535 12801
rect 20717 12767 20775 12773
rect 20717 12733 20729 12767
rect 20763 12733 20775 12767
rect 23492 12764 23520 12795
rect 31662 12792 31668 12844
rect 31720 12832 31726 12844
rect 32309 12835 32367 12841
rect 32309 12832 32321 12835
rect 31720 12804 32321 12832
rect 31720 12792 31726 12804
rect 32309 12801 32321 12804
rect 32355 12801 32367 12835
rect 33594 12832 33600 12844
rect 32309 12795 32367 12801
rect 33152 12804 33600 12832
rect 33152 12773 33180 12804
rect 33594 12792 33600 12804
rect 33652 12792 33658 12844
rect 35710 12792 35716 12844
rect 35768 12832 35774 12844
rect 36081 12835 36139 12841
rect 36081 12832 36093 12835
rect 35768 12804 36093 12832
rect 35768 12792 35774 12804
rect 36081 12801 36093 12804
rect 36127 12801 36139 12835
rect 36244 12835 36302 12841
rect 36244 12832 36256 12835
rect 36081 12795 36139 12801
rect 36188 12804 36256 12832
rect 33137 12767 33195 12773
rect 33137 12764 33149 12767
rect 23492 12736 33149 12764
rect 20717 12727 20775 12733
rect 33137 12733 33149 12736
rect 33183 12733 33195 12767
rect 33410 12764 33416 12776
rect 33371 12736 33416 12764
rect 33137 12727 33195 12733
rect 18966 12656 18972 12708
rect 19024 12696 19030 12708
rect 20732 12696 20760 12727
rect 33410 12724 33416 12736
rect 33468 12724 33474 12776
rect 19024 12668 20760 12696
rect 19024 12656 19030 12668
rect 25590 12656 25596 12708
rect 25648 12696 25654 12708
rect 29178 12696 29184 12708
rect 25648 12668 29184 12696
rect 25648 12656 25654 12668
rect 29178 12656 29184 12668
rect 29236 12656 29242 12708
rect 36188 12696 36216 12804
rect 36244 12801 36256 12804
rect 36290 12801 36302 12835
rect 36244 12795 36302 12801
rect 36354 12792 36360 12844
rect 36412 12832 36418 12844
rect 36538 12841 36544 12844
rect 36495 12835 36544 12841
rect 36412 12804 36457 12832
rect 36412 12792 36418 12804
rect 36495 12801 36507 12835
rect 36541 12801 36544 12835
rect 36495 12795 36544 12801
rect 36538 12792 36544 12795
rect 36596 12792 36602 12844
rect 38654 12832 38660 12844
rect 38615 12804 38660 12832
rect 38654 12792 38660 12804
rect 38712 12792 38718 12844
rect 37277 12699 37335 12705
rect 37277 12696 37289 12699
rect 36188 12668 37289 12696
rect 37277 12665 37289 12668
rect 37323 12665 37335 12699
rect 37277 12659 37335 12665
rect 19150 12628 19156 12640
rect 18892 12600 19156 12628
rect 16761 12591 16819 12597
rect 19150 12588 19156 12600
rect 19208 12588 19214 12640
rect 27065 12631 27123 12637
rect 27065 12597 27077 12631
rect 27111 12628 27123 12631
rect 27246 12628 27252 12640
rect 27111 12600 27252 12628
rect 27111 12597 27123 12600
rect 27065 12591 27123 12597
rect 27246 12588 27252 12600
rect 27304 12588 27310 12640
rect 36722 12628 36728 12640
rect 36683 12600 36728 12628
rect 36722 12588 36728 12600
rect 36780 12588 36786 12640
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 7558 12424 7564 12436
rect 7519 12396 7564 12424
rect 7558 12384 7564 12396
rect 7616 12384 7622 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8128 12396 9045 12424
rect 3786 12288 3792 12300
rect 3747 12260 3792 12288
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 5592 12260 6101 12288
rect 5592 12248 5598 12260
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6178 12248 6184 12300
rect 6236 12288 6242 12300
rect 8018 12288 8024 12300
rect 6236 12260 6281 12288
rect 7979 12260 8024 12288
rect 6236 12248 6242 12260
rect 8018 12248 8024 12260
rect 8076 12248 8082 12300
rect 2590 12220 2596 12232
rect 2551 12192 2596 12220
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 2731 12192 5672 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 3050 12112 3056 12164
rect 3108 12152 3114 12164
rect 4034 12155 4092 12161
rect 4034 12152 4046 12155
rect 3108 12124 4046 12152
rect 3108 12112 3114 12124
rect 4034 12121 4046 12124
rect 4080 12121 4092 12155
rect 4034 12115 4092 12121
rect 2866 12084 2872 12096
rect 2827 12056 2872 12084
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5534 12084 5540 12096
rect 5215 12056 5540 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 5644 12093 5672 12192
rect 7006 12180 7012 12232
rect 7064 12220 7070 12232
rect 8128 12229 8156 12396
rect 9033 12393 9045 12396
rect 9079 12424 9091 12427
rect 14090 12424 14096 12436
rect 9079 12396 12434 12424
rect 14051 12396 14096 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 8294 12316 8300 12368
rect 8352 12356 8358 12368
rect 9122 12356 9128 12368
rect 8352 12328 9128 12356
rect 8352 12316 8358 12328
rect 9122 12316 9128 12328
rect 9180 12356 9186 12368
rect 12406 12356 12434 12396
rect 14090 12384 14096 12396
rect 14148 12384 14154 12436
rect 18230 12424 18236 12436
rect 14200 12396 18236 12424
rect 14200 12356 14228 12396
rect 18230 12384 18236 12396
rect 18288 12384 18294 12436
rect 21174 12384 21180 12436
rect 21232 12424 21238 12436
rect 21913 12427 21971 12433
rect 21913 12424 21925 12427
rect 21232 12396 21925 12424
rect 21232 12384 21238 12396
rect 21913 12393 21925 12396
rect 21959 12424 21971 12427
rect 22186 12424 22192 12436
rect 21959 12396 22192 12424
rect 21959 12393 21971 12396
rect 21913 12387 21971 12393
rect 22186 12384 22192 12396
rect 22244 12384 22250 12436
rect 22370 12384 22376 12436
rect 22428 12424 22434 12436
rect 22557 12427 22615 12433
rect 22557 12424 22569 12427
rect 22428 12396 22569 12424
rect 22428 12384 22434 12396
rect 22557 12393 22569 12396
rect 22603 12424 22615 12427
rect 27154 12424 27160 12436
rect 22603 12396 27160 12424
rect 22603 12393 22615 12396
rect 22557 12387 22615 12393
rect 27154 12384 27160 12396
rect 27212 12384 27218 12436
rect 35618 12384 35624 12436
rect 35676 12424 35682 12436
rect 35897 12427 35955 12433
rect 35897 12424 35909 12427
rect 35676 12396 35909 12424
rect 35676 12384 35682 12396
rect 35897 12393 35909 12396
rect 35943 12424 35955 12427
rect 36538 12424 36544 12436
rect 35943 12396 36544 12424
rect 35943 12393 35955 12396
rect 35897 12387 35955 12393
rect 36538 12384 36544 12396
rect 36596 12384 36602 12436
rect 37458 12384 37464 12436
rect 37516 12424 37522 12436
rect 38197 12427 38255 12433
rect 38197 12424 38209 12427
rect 37516 12396 38209 12424
rect 37516 12384 37522 12396
rect 38197 12393 38209 12396
rect 38243 12393 38255 12427
rect 38197 12387 38255 12393
rect 17497 12359 17555 12365
rect 9180 12328 9536 12356
rect 12406 12328 14228 12356
rect 16316 12328 17356 12356
rect 9180 12316 9186 12328
rect 9508 12297 9536 12328
rect 9493 12291 9551 12297
rect 9493 12257 9505 12291
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 16114 12248 16120 12300
rect 16172 12288 16178 12300
rect 16316 12288 16344 12328
rect 16172 12260 16344 12288
rect 17328 12288 17356 12328
rect 17497 12325 17509 12359
rect 17543 12356 17555 12359
rect 18138 12356 18144 12368
rect 17543 12328 18144 12356
rect 17543 12325 17555 12328
rect 17497 12319 17555 12325
rect 18138 12316 18144 12328
rect 18196 12316 18202 12368
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 19337 12359 19395 12365
rect 19337 12356 19349 12359
rect 19300 12328 19349 12356
rect 19300 12316 19306 12328
rect 19337 12325 19349 12328
rect 19383 12356 19395 12359
rect 28445 12359 28503 12365
rect 28445 12356 28457 12359
rect 19383 12328 28457 12356
rect 19383 12325 19395 12328
rect 19337 12319 19395 12325
rect 28445 12325 28457 12328
rect 28491 12356 28503 12359
rect 29362 12356 29368 12368
rect 28491 12328 29368 12356
rect 28491 12325 28503 12328
rect 28445 12319 28503 12325
rect 29362 12316 29368 12328
rect 29420 12316 29426 12368
rect 30653 12359 30711 12365
rect 30653 12325 30665 12359
rect 30699 12356 30711 12359
rect 30834 12356 30840 12368
rect 30699 12328 30840 12356
rect 30699 12325 30711 12328
rect 30653 12319 30711 12325
rect 30834 12316 30840 12328
rect 30892 12356 30898 12368
rect 31478 12356 31484 12368
rect 30892 12328 31484 12356
rect 30892 12316 30898 12328
rect 31478 12316 31484 12328
rect 31536 12316 31542 12368
rect 18966 12288 18972 12300
rect 17328 12260 18972 12288
rect 16172 12248 16178 12260
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 7064 12192 7757 12220
rect 7064 12180 7070 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 8297 12223 8355 12229
rect 8297 12189 8309 12223
rect 8343 12220 8355 12223
rect 8386 12220 8392 12232
rect 8343 12192 8392 12220
rect 8343 12189 8355 12192
rect 8297 12183 8355 12189
rect 7944 12152 7972 12183
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 9766 12229 9772 12232
rect 9760 12183 9772 12229
rect 9824 12220 9830 12232
rect 11333 12223 11391 12229
rect 9824 12192 9860 12220
rect 9766 12180 9772 12183
rect 9824 12180 9830 12192
rect 11333 12189 11345 12223
rect 11379 12220 11391 12223
rect 11422 12220 11428 12232
rect 11379 12192 11428 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 11606 12229 11612 12232
rect 11600 12183 11612 12229
rect 11664 12220 11670 12232
rect 13541 12223 13599 12229
rect 11664 12192 11700 12220
rect 11606 12180 11612 12183
rect 11664 12180 11670 12192
rect 13541 12189 13553 12223
rect 13587 12220 13599 12223
rect 13906 12220 13912 12232
rect 13587 12192 13912 12220
rect 13587 12189 13599 12192
rect 13541 12183 13599 12189
rect 13906 12180 13912 12192
rect 13964 12180 13970 12232
rect 15194 12220 15200 12232
rect 15252 12229 15258 12232
rect 15164 12192 15200 12220
rect 15194 12180 15200 12192
rect 15252 12183 15264 12229
rect 15470 12220 15476 12232
rect 15431 12192 15476 12220
rect 15252 12180 15258 12183
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16316 12229 16344 12260
rect 16209 12223 16267 12229
rect 16209 12220 16221 12223
rect 16080 12192 16221 12220
rect 16080 12180 16086 12192
rect 16209 12189 16221 12192
rect 16255 12189 16267 12223
rect 16209 12183 16267 12189
rect 16301 12223 16359 12229
rect 16301 12189 16313 12223
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12220 16635 12223
rect 16758 12220 16764 12232
rect 16623 12192 16764 12220
rect 16623 12189 16635 12192
rect 16577 12183 16635 12189
rect 9582 12152 9588 12164
rect 7944 12124 9588 12152
rect 9582 12112 9588 12124
rect 9640 12112 9646 12164
rect 12342 12112 12348 12164
rect 12400 12152 12406 12164
rect 13357 12155 13415 12161
rect 13357 12152 13369 12155
rect 12400 12124 13369 12152
rect 12400 12112 12406 12124
rect 13357 12121 13369 12124
rect 13403 12152 13415 12155
rect 13722 12152 13728 12164
rect 13403 12124 13728 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 13722 12112 13728 12124
rect 13780 12112 13786 12164
rect 16408 12152 16436 12183
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12220 17187 12223
rect 17494 12220 17500 12232
rect 17175 12192 17500 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 18230 12220 18236 12232
rect 18191 12192 18236 12220
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 18340 12229 18368 12260
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 18325 12223 18383 12229
rect 18601 12223 18659 12229
rect 18325 12189 18337 12223
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 18422 12217 18480 12223
rect 18422 12183 18434 12217
rect 18468 12214 18480 12217
rect 18468 12186 18552 12214
rect 18468 12183 18480 12186
rect 18422 12177 18480 12183
rect 14752 12124 16436 12152
rect 5629 12087 5687 12093
rect 5629 12053 5641 12087
rect 5675 12053 5687 12087
rect 5629 12047 5687 12053
rect 5997 12087 6055 12093
rect 5997 12053 6009 12087
rect 6043 12084 6055 12087
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6043 12056 6929 12084
rect 6043 12053 6055 12056
rect 5997 12047 6055 12053
rect 6917 12053 6929 12056
rect 6963 12084 6975 12087
rect 7098 12084 7104 12096
rect 6963 12056 7104 12084
rect 6963 12053 6975 12056
rect 6917 12047 6975 12053
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 9674 12044 9680 12096
rect 9732 12084 9738 12096
rect 10873 12087 10931 12093
rect 10873 12084 10885 12087
rect 9732 12056 10885 12084
rect 9732 12044 9738 12056
rect 10873 12053 10885 12056
rect 10919 12053 10931 12087
rect 10873 12047 10931 12053
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 12710 12084 12716 12096
rect 11756 12056 12716 12084
rect 11756 12044 11762 12056
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 13173 12087 13231 12093
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 14752 12084 14780 12124
rect 16666 12112 16672 12164
rect 16724 12152 16730 12164
rect 17313 12155 17371 12161
rect 17313 12152 17325 12155
rect 16724 12124 17325 12152
rect 16724 12112 16730 12124
rect 17313 12121 17325 12124
rect 17359 12121 17371 12155
rect 17313 12115 17371 12121
rect 13219 12056 14780 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 14826 12044 14832 12096
rect 14884 12084 14890 12096
rect 15933 12087 15991 12093
rect 15933 12084 15945 12087
rect 14884 12056 15945 12084
rect 14884 12044 14890 12056
rect 15933 12053 15945 12056
rect 15979 12053 15991 12087
rect 15933 12047 15991 12053
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 18138 12084 18144 12096
rect 18003 12056 18144 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 18322 12044 18328 12096
rect 18380 12084 18386 12096
rect 18524 12084 18552 12186
rect 18601 12189 18613 12223
rect 18647 12220 18659 12223
rect 18690 12220 18696 12232
rect 18647 12192 18696 12220
rect 18647 12189 18659 12192
rect 18601 12183 18659 12189
rect 18690 12180 18696 12192
rect 18748 12220 18754 12232
rect 19260 12220 19288 12316
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12288 19855 12291
rect 24489 12291 24547 12297
rect 19843 12260 21128 12288
rect 19843 12257 19855 12260
rect 19797 12251 19855 12257
rect 20162 12220 20168 12232
rect 18748 12192 19288 12220
rect 20123 12192 20168 12220
rect 18748 12180 18754 12192
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 20622 12180 20628 12232
rect 20680 12180 20686 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 20855 12223 20913 12229
rect 20855 12220 20867 12223
rect 20772 12192 20867 12220
rect 20772 12180 20778 12192
rect 20855 12189 20867 12192
rect 20901 12189 20913 12223
rect 20990 12220 20996 12232
rect 20951 12192 20996 12220
rect 20855 12183 20913 12189
rect 20990 12180 20996 12192
rect 21048 12180 21054 12232
rect 21100 12229 21128 12260
rect 24489 12257 24501 12291
rect 24535 12288 24547 12291
rect 24578 12288 24584 12300
rect 24535 12260 24584 12288
rect 24535 12257 24547 12260
rect 24489 12251 24547 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 25774 12288 25780 12300
rect 25424 12260 25780 12288
rect 21085 12223 21143 12229
rect 21085 12189 21097 12223
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12189 21327 12223
rect 24596 12220 24624 12248
rect 25179 12223 25237 12229
rect 25179 12220 25191 12223
rect 24596 12192 25191 12220
rect 21269 12183 21327 12189
rect 25179 12189 25191 12192
rect 25225 12189 25237 12223
rect 25314 12220 25320 12232
rect 25275 12192 25320 12220
rect 25179 12183 25237 12189
rect 19978 12152 19984 12164
rect 19891 12124 19984 12152
rect 19978 12112 19984 12124
rect 20036 12152 20042 12164
rect 20640 12152 20668 12180
rect 20036 12124 20668 12152
rect 20036 12112 20042 12124
rect 20622 12084 20628 12096
rect 18380 12056 18552 12084
rect 20583 12056 20628 12084
rect 18380 12044 18386 12056
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 21284 12084 21312 12183
rect 25314 12180 25320 12192
rect 25372 12180 25378 12232
rect 25424 12229 25452 12260
rect 25774 12248 25780 12260
rect 25832 12248 25838 12300
rect 31754 12288 31760 12300
rect 31128 12260 31760 12288
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12189 25467 12223
rect 25409 12183 25467 12189
rect 25498 12180 25504 12232
rect 25556 12220 25562 12232
rect 31128 12229 31156 12260
rect 31754 12248 31760 12260
rect 31812 12288 31818 12300
rect 32490 12288 32496 12300
rect 31812 12260 32496 12288
rect 31812 12248 31818 12260
rect 32490 12248 32496 12260
rect 32548 12248 32554 12300
rect 25593 12223 25651 12229
rect 25593 12220 25605 12223
rect 25556 12192 25605 12220
rect 25556 12180 25562 12192
rect 25593 12189 25605 12192
rect 25639 12220 25651 12223
rect 27433 12223 27491 12229
rect 27433 12220 27445 12223
rect 25639 12192 27445 12220
rect 25639 12189 25651 12192
rect 25593 12183 25651 12189
rect 27433 12189 27445 12192
rect 27479 12189 27491 12223
rect 27433 12183 27491 12189
rect 31113 12223 31171 12229
rect 31113 12189 31125 12223
rect 31159 12189 31171 12223
rect 31294 12220 31300 12232
rect 31255 12192 31300 12220
rect 31113 12183 31171 12189
rect 31294 12180 31300 12192
rect 31352 12180 31358 12232
rect 31389 12223 31447 12229
rect 31389 12189 31401 12223
rect 31435 12189 31447 12223
rect 31389 12183 31447 12189
rect 21726 12112 21732 12164
rect 21784 12152 21790 12164
rect 21821 12155 21879 12161
rect 21821 12152 21833 12155
rect 21784 12124 21833 12152
rect 21784 12112 21790 12124
rect 21821 12121 21833 12124
rect 21867 12121 21879 12155
rect 21821 12115 21879 12121
rect 27617 12155 27675 12161
rect 27617 12121 27629 12155
rect 27663 12152 27675 12155
rect 28258 12152 28264 12164
rect 27663 12124 28264 12152
rect 27663 12121 27675 12124
rect 27617 12115 27675 12121
rect 28258 12112 28264 12124
rect 28316 12112 28322 12164
rect 31018 12112 31024 12164
rect 31076 12152 31082 12164
rect 31404 12152 31432 12183
rect 31478 12180 31484 12232
rect 31536 12220 31542 12232
rect 33597 12223 33655 12229
rect 31536 12192 31581 12220
rect 31536 12180 31542 12192
rect 33597 12189 33609 12223
rect 33643 12220 33655 12223
rect 34514 12220 34520 12232
rect 33643 12192 34520 12220
rect 33643 12189 33655 12192
rect 33597 12183 33655 12189
rect 34514 12180 34520 12192
rect 34572 12180 34578 12232
rect 36817 12223 36875 12229
rect 36817 12189 36829 12223
rect 36863 12220 36875 12223
rect 38378 12220 38384 12232
rect 36863 12192 38384 12220
rect 36863 12189 36875 12192
rect 36817 12183 36875 12189
rect 38378 12180 38384 12192
rect 38436 12180 38442 12232
rect 31076 12124 31432 12152
rect 31757 12155 31815 12161
rect 31076 12112 31082 12124
rect 31757 12121 31769 12155
rect 31803 12152 31815 12155
rect 33330 12155 33388 12161
rect 33330 12152 33342 12155
rect 31803 12124 33342 12152
rect 31803 12121 31815 12124
rect 31757 12115 31815 12121
rect 33330 12121 33342 12124
rect 33376 12121 33388 12155
rect 33330 12115 33388 12121
rect 36722 12112 36728 12164
rect 36780 12152 36786 12164
rect 37062 12155 37120 12161
rect 37062 12152 37074 12155
rect 36780 12124 37074 12152
rect 36780 12112 36786 12124
rect 37062 12121 37074 12124
rect 37108 12121 37120 12155
rect 37062 12115 37120 12121
rect 22462 12084 22468 12096
rect 21284 12056 22468 12084
rect 22462 12044 22468 12056
rect 22520 12084 22526 12096
rect 23109 12087 23167 12093
rect 23109 12084 23121 12087
rect 22520 12056 23121 12084
rect 22520 12044 22526 12056
rect 23109 12053 23121 12056
rect 23155 12084 23167 12087
rect 23474 12084 23480 12096
rect 23155 12056 23480 12084
rect 23155 12053 23167 12056
rect 23109 12047 23167 12053
rect 23474 12044 23480 12056
rect 23532 12044 23538 12096
rect 24946 12084 24952 12096
rect 24907 12056 24952 12084
rect 24946 12044 24952 12056
rect 25004 12044 25010 12096
rect 32217 12087 32275 12093
rect 32217 12053 32229 12087
rect 32263 12084 32275 12087
rect 32398 12084 32404 12096
rect 32263 12056 32404 12084
rect 32263 12053 32275 12056
rect 32217 12047 32275 12053
rect 32398 12044 32404 12056
rect 32456 12044 32462 12096
rect 34606 12044 34612 12096
rect 34664 12084 34670 12096
rect 35802 12084 35808 12096
rect 34664 12056 35808 12084
rect 34664 12044 34670 12056
rect 35802 12044 35808 12056
rect 35860 12044 35866 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 3050 11880 3056 11892
rect 3011 11852 3056 11880
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 9858 11880 9864 11892
rect 5859 11852 9864 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 13722 11880 13728 11892
rect 13683 11852 13728 11880
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 15010 11880 15016 11892
rect 14792 11852 15016 11880
rect 14792 11840 14798 11852
rect 15010 11840 15016 11852
rect 15068 11880 15074 11892
rect 15562 11880 15568 11892
rect 15068 11852 15568 11880
rect 15068 11840 15074 11852
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 16666 11840 16672 11892
rect 16724 11880 16730 11892
rect 17037 11883 17095 11889
rect 17037 11880 17049 11883
rect 16724 11852 17049 11880
rect 16724 11840 16730 11852
rect 17037 11849 17049 11852
rect 17083 11849 17095 11883
rect 19889 11883 19947 11889
rect 17037 11843 17095 11849
rect 17144 11852 19288 11880
rect 6822 11772 6828 11824
rect 6880 11772 6886 11824
rect 14826 11772 14832 11824
rect 14884 11821 14890 11824
rect 14884 11812 14896 11821
rect 17144 11812 17172 11852
rect 19260 11812 19288 11852
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 19978 11880 19984 11892
rect 19935 11852 19984 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 23293 11883 23351 11889
rect 23293 11849 23305 11883
rect 23339 11880 23351 11883
rect 25314 11880 25320 11892
rect 23339 11852 25320 11880
rect 23339 11849 23351 11852
rect 23293 11843 23351 11849
rect 20438 11812 20444 11824
rect 14884 11784 14929 11812
rect 15028 11784 17172 11812
rect 17328 11784 18368 11812
rect 19260 11784 20444 11812
rect 14884 11775 14896 11784
rect 14884 11772 14890 11775
rect 2866 11744 2872 11756
rect 2827 11716 2872 11744
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 4706 11744 4712 11756
rect 4667 11716 4712 11744
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 5534 11744 5540 11756
rect 5495 11716 5540 11744
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6840 11744 6868 11772
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6696 11716 6929 11744
rect 6696 11704 6702 11716
rect 6917 11713 6929 11716
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 8018 11704 8024 11756
rect 8076 11744 8082 11756
rect 8858 11747 8916 11753
rect 8858 11744 8870 11747
rect 8076 11716 8870 11744
rect 8076 11704 8082 11716
rect 8858 11713 8870 11716
rect 8904 11713 8916 11747
rect 9122 11744 9128 11756
rect 9083 11716 9128 11744
rect 8858 11707 8916 11713
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 11790 11744 11796 11756
rect 11751 11716 11796 11744
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 15028 11744 15056 11784
rect 14108 11716 15056 11744
rect 15105 11747 15163 11753
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 4433 11679 4491 11685
rect 4433 11676 4445 11679
rect 2648 11648 4445 11676
rect 2648 11636 2654 11648
rect 4433 11645 4445 11648
rect 4479 11645 4491 11679
rect 4433 11639 4491 11645
rect 5169 11679 5227 11685
rect 5169 11645 5181 11679
rect 5215 11645 5227 11679
rect 5169 11639 5227 11645
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 6457 11679 6515 11685
rect 5675 11648 6408 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 5184 11608 5212 11639
rect 5534 11608 5540 11620
rect 5184 11580 5540 11608
rect 5534 11568 5540 11580
rect 5592 11608 5598 11620
rect 5718 11608 5724 11620
rect 5592 11580 5724 11608
rect 5592 11568 5598 11580
rect 5718 11568 5724 11580
rect 5776 11568 5782 11620
rect 6380 11540 6408 11648
rect 6457 11645 6469 11679
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 6472 11608 6500 11639
rect 6730 11636 6736 11688
rect 6788 11676 6794 11688
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6788 11648 6837 11676
rect 6788 11636 6794 11648
rect 6825 11645 6837 11648
rect 6871 11645 6883 11679
rect 6825 11639 6883 11645
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11517 11679 11575 11685
rect 11517 11676 11529 11679
rect 11388 11648 11529 11676
rect 11388 11636 11394 11648
rect 11517 11645 11529 11648
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 6472 11580 8248 11608
rect 8220 11552 8248 11580
rect 6914 11540 6920 11552
rect 6380 11512 6920 11540
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7558 11540 7564 11552
rect 7147 11512 7564 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 7745 11543 7803 11549
rect 7745 11509 7757 11543
rect 7791 11540 7803 11543
rect 7834 11540 7840 11552
rect 7791 11512 7840 11540
rect 7791 11509 7803 11512
rect 7745 11503 7803 11509
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 8202 11500 8208 11552
rect 8260 11500 8266 11552
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 14108 11540 14136 11716
rect 15105 11713 15117 11747
rect 15151 11744 15163 11747
rect 15470 11744 15476 11756
rect 15151 11716 15476 11744
rect 15151 11713 15163 11716
rect 15105 11707 15163 11713
rect 15470 11704 15476 11716
rect 15528 11744 15534 11756
rect 17328 11744 17356 11784
rect 18340 11756 18368 11784
rect 20438 11772 20444 11784
rect 20496 11772 20502 11824
rect 20622 11772 20628 11824
rect 20680 11812 20686 11824
rect 21002 11815 21060 11821
rect 21002 11812 21014 11815
rect 20680 11784 21014 11812
rect 20680 11772 20686 11784
rect 21002 11781 21014 11784
rect 21048 11781 21060 11815
rect 23308 11812 23336 11843
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 29638 11880 29644 11892
rect 29599 11852 29644 11880
rect 29638 11840 29644 11852
rect 29696 11840 29702 11892
rect 31294 11840 31300 11892
rect 31352 11880 31358 11892
rect 32125 11883 32183 11889
rect 32125 11880 32137 11883
rect 31352 11852 32137 11880
rect 31352 11840 31358 11852
rect 32125 11849 32137 11852
rect 32171 11849 32183 11883
rect 32125 11843 32183 11849
rect 34698 11840 34704 11892
rect 34756 11880 34762 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 34756 11852 35173 11880
rect 34756 11840 34762 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 35161 11843 35219 11849
rect 21002 11775 21060 11781
rect 22480 11784 23336 11812
rect 15528 11716 17356 11744
rect 15528 11704 15534 11716
rect 18138 11704 18144 11756
rect 18196 11753 18202 11756
rect 18196 11744 18208 11753
rect 18196 11716 18241 11744
rect 18196 11707 18208 11716
rect 18196 11704 18202 11707
rect 18322 11704 18328 11756
rect 18380 11744 18386 11756
rect 18417 11747 18475 11753
rect 18417 11744 18429 11747
rect 18380 11716 18429 11744
rect 18380 11704 18386 11716
rect 18417 11713 18429 11716
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11744 19027 11747
rect 19334 11744 19340 11756
rect 19015 11716 19340 11744
rect 19015 11713 19027 11716
rect 18969 11707 19027 11713
rect 19334 11704 19340 11716
rect 19392 11704 19398 11756
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 20714 11744 20720 11756
rect 20588 11716 20720 11744
rect 20588 11704 20594 11716
rect 20714 11704 20720 11716
rect 20772 11744 20778 11756
rect 22370 11744 22376 11756
rect 20772 11716 22376 11744
rect 20772 11704 20778 11716
rect 22370 11704 22376 11716
rect 22428 11704 22434 11756
rect 22480 11753 22508 11784
rect 24946 11772 24952 11824
rect 25004 11812 25010 11824
rect 25102 11815 25160 11821
rect 25102 11812 25114 11815
rect 25004 11784 25114 11812
rect 25004 11772 25010 11784
rect 25102 11781 25114 11784
rect 25148 11781 25160 11815
rect 25102 11775 25160 11781
rect 22465 11747 22523 11753
rect 22465 11713 22477 11747
rect 22511 11713 22523 11747
rect 22465 11707 22523 11713
rect 22554 11704 22560 11756
rect 22612 11744 22618 11756
rect 22612 11716 22657 11744
rect 22612 11704 22618 11716
rect 22738 11704 22744 11756
rect 22796 11744 22802 11756
rect 22796 11716 22841 11744
rect 22796 11704 22802 11716
rect 23106 11704 23112 11756
rect 23164 11744 23170 11756
rect 23201 11747 23259 11753
rect 23201 11744 23213 11747
rect 23164 11716 23213 11744
rect 23164 11704 23170 11716
rect 23201 11713 23213 11716
rect 23247 11713 23259 11747
rect 23382 11744 23388 11756
rect 23343 11716 23388 11744
rect 23201 11707 23259 11713
rect 23382 11704 23388 11716
rect 23440 11704 23446 11756
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 23532 11716 25912 11744
rect 23532 11704 23538 11716
rect 21269 11679 21327 11685
rect 21269 11645 21281 11679
rect 21315 11676 21327 11679
rect 21542 11676 21548 11688
rect 21315 11648 21548 11676
rect 21315 11645 21327 11648
rect 21269 11639 21327 11645
rect 21542 11636 21548 11648
rect 21600 11676 21606 11688
rect 24854 11676 24860 11688
rect 21600 11648 24860 11676
rect 21600 11636 21606 11648
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 19150 11608 19156 11620
rect 19111 11580 19156 11608
rect 19150 11568 19156 11580
rect 19208 11568 19214 11620
rect 22738 11608 22744 11620
rect 21744 11580 22744 11608
rect 12308 11512 14136 11540
rect 15841 11543 15899 11549
rect 12308 11500 12314 11512
rect 15841 11509 15853 11543
rect 15887 11540 15899 11543
rect 16022 11540 16028 11552
rect 15887 11512 16028 11540
rect 15887 11509 15899 11512
rect 15841 11503 15899 11509
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 21744 11540 21772 11580
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 25884 11608 25912 11716
rect 28258 11704 28264 11756
rect 28316 11744 28322 11756
rect 28353 11747 28411 11753
rect 28353 11744 28365 11747
rect 28316 11716 28365 11744
rect 28316 11704 28322 11716
rect 28353 11713 28365 11716
rect 28399 11713 28411 11747
rect 29656 11744 29684 11840
rect 30834 11812 30840 11824
rect 30484 11784 30840 11812
rect 30484 11753 30512 11784
rect 30834 11772 30840 11784
rect 30892 11772 30898 11824
rect 31662 11772 31668 11824
rect 31720 11812 31726 11824
rect 32493 11815 32551 11821
rect 32493 11812 32505 11815
rect 31720 11784 32505 11812
rect 31720 11772 31726 11784
rect 32493 11781 32505 11784
rect 32539 11781 32551 11815
rect 32493 11775 32551 11781
rect 35437 11815 35495 11821
rect 35437 11781 35449 11815
rect 35483 11812 35495 11815
rect 36262 11812 36268 11824
rect 35483 11784 36268 11812
rect 35483 11781 35495 11784
rect 35437 11775 35495 11781
rect 36262 11772 36268 11784
rect 36320 11772 36326 11824
rect 39482 11812 39488 11824
rect 39443 11784 39488 11812
rect 39482 11772 39488 11784
rect 39540 11772 39546 11824
rect 30377 11747 30435 11753
rect 30377 11744 30389 11747
rect 29656 11716 30389 11744
rect 28353 11707 28411 11713
rect 30377 11713 30389 11716
rect 30423 11713 30435 11747
rect 30377 11707 30435 11713
rect 30469 11747 30527 11753
rect 30469 11713 30481 11747
rect 30515 11713 30527 11747
rect 30469 11707 30527 11713
rect 28368 11676 28396 11707
rect 30558 11704 30564 11756
rect 30616 11744 30622 11756
rect 30745 11747 30803 11753
rect 30616 11716 30661 11744
rect 30616 11704 30622 11716
rect 30745 11713 30757 11747
rect 30791 11744 30803 11747
rect 31754 11744 31760 11756
rect 30791 11716 31760 11744
rect 30791 11713 30803 11716
rect 30745 11707 30803 11713
rect 31754 11704 31760 11716
rect 31812 11704 31818 11756
rect 32309 11747 32367 11753
rect 32309 11713 32321 11747
rect 32355 11744 32367 11747
rect 32398 11744 32404 11756
rect 32355 11716 32404 11744
rect 32355 11713 32367 11716
rect 32309 11707 32367 11713
rect 32398 11704 32404 11716
rect 32456 11704 32462 11756
rect 33226 11704 33232 11756
rect 33284 11744 33290 11756
rect 33410 11744 33416 11756
rect 33284 11716 33416 11744
rect 33284 11704 33290 11716
rect 33410 11704 33416 11716
rect 33468 11744 33474 11756
rect 34517 11747 34575 11753
rect 34517 11744 34529 11747
rect 33468 11716 34529 11744
rect 33468 11704 33474 11716
rect 34517 11713 34529 11716
rect 34563 11713 34575 11747
rect 35342 11744 35348 11756
rect 35255 11716 35348 11744
rect 34517 11707 34575 11713
rect 35342 11704 35348 11716
rect 35400 11704 35406 11756
rect 35526 11744 35532 11756
rect 35487 11716 35532 11744
rect 35526 11704 35532 11716
rect 35584 11704 35590 11756
rect 35618 11704 35624 11756
rect 35676 11744 35682 11756
rect 35713 11747 35771 11753
rect 35713 11744 35725 11747
rect 35676 11716 35725 11744
rect 35676 11704 35682 11716
rect 35713 11713 35725 11716
rect 35759 11713 35771 11747
rect 35713 11707 35771 11713
rect 37734 11704 37740 11756
rect 37792 11744 37798 11756
rect 38565 11747 38623 11753
rect 38565 11744 38577 11747
rect 37792 11716 38577 11744
rect 37792 11704 37798 11716
rect 38565 11713 38577 11716
rect 38611 11713 38623 11747
rect 38565 11707 38623 11713
rect 33244 11676 33272 11704
rect 28368 11648 33272 11676
rect 35360 11676 35388 11704
rect 38286 11676 38292 11688
rect 35360 11648 35756 11676
rect 38247 11648 38292 11676
rect 35728 11620 35756 11648
rect 38286 11636 38292 11648
rect 38344 11636 38350 11688
rect 28537 11611 28595 11617
rect 28537 11608 28549 11611
rect 25884 11580 28549 11608
rect 28537 11577 28549 11580
rect 28583 11608 28595 11611
rect 33962 11608 33968 11620
rect 28583 11580 33968 11608
rect 28583 11577 28595 11580
rect 28537 11571 28595 11577
rect 33962 11568 33968 11580
rect 34020 11568 34026 11620
rect 35710 11568 35716 11620
rect 35768 11568 35774 11620
rect 39114 11568 39120 11620
rect 39172 11608 39178 11620
rect 39301 11611 39359 11617
rect 39301 11608 39313 11611
rect 39172 11580 39313 11608
rect 39172 11568 39178 11580
rect 39301 11577 39313 11580
rect 39347 11577 39359 11611
rect 58158 11608 58164 11620
rect 58119 11580 58164 11608
rect 39301 11571 39359 11577
rect 58158 11568 58164 11580
rect 58216 11568 58222 11620
rect 16816 11512 21772 11540
rect 16816 11500 16822 11512
rect 21818 11500 21824 11552
rect 21876 11540 21882 11552
rect 22097 11543 22155 11549
rect 22097 11540 22109 11543
rect 21876 11512 22109 11540
rect 21876 11500 21882 11512
rect 22097 11509 22109 11512
rect 22143 11509 22155 11543
rect 22097 11503 22155 11509
rect 22186 11500 22192 11552
rect 22244 11540 22250 11552
rect 23106 11540 23112 11552
rect 22244 11512 23112 11540
rect 22244 11500 22250 11512
rect 23106 11500 23112 11512
rect 23164 11540 23170 11552
rect 23845 11543 23903 11549
rect 23845 11540 23857 11543
rect 23164 11512 23857 11540
rect 23164 11500 23170 11512
rect 23845 11509 23857 11512
rect 23891 11509 23903 11543
rect 23845 11503 23903 11509
rect 25038 11500 25044 11552
rect 25096 11540 25102 11552
rect 26237 11543 26295 11549
rect 26237 11540 26249 11543
rect 25096 11512 26249 11540
rect 25096 11500 25102 11512
rect 26237 11509 26249 11512
rect 26283 11509 26295 11543
rect 26237 11503 26295 11509
rect 30101 11543 30159 11549
rect 30101 11509 30113 11543
rect 30147 11540 30159 11543
rect 30282 11540 30288 11552
rect 30147 11512 30288 11540
rect 30147 11509 30159 11512
rect 30101 11503 30159 11509
rect 30282 11500 30288 11512
rect 30340 11500 30346 11552
rect 34609 11543 34667 11549
rect 34609 11509 34621 11543
rect 34655 11540 34667 11543
rect 38102 11540 38108 11552
rect 34655 11512 38108 11540
rect 34655 11509 34667 11512
rect 34609 11503 34667 11509
rect 38102 11500 38108 11512
rect 38160 11500 38166 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 8018 11336 8024 11348
rect 7979 11308 8024 11336
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 18690 11336 18696 11348
rect 18651 11308 18696 11336
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 20530 11336 20536 11348
rect 20491 11308 20536 11336
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 26234 11336 26240 11348
rect 25976 11308 26240 11336
rect 7190 11228 7196 11280
rect 7248 11268 7254 11280
rect 11517 11271 11575 11277
rect 7248 11240 7696 11268
rect 7248 11228 7254 11240
rect 7558 11200 7564 11212
rect 7519 11172 7564 11200
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 7668 11209 7696 11240
rect 11517 11237 11529 11271
rect 11563 11268 11575 11271
rect 11606 11268 11612 11280
rect 11563 11240 11612 11268
rect 11563 11237 11575 11240
rect 11517 11231 11575 11237
rect 11606 11228 11612 11240
rect 11664 11228 11670 11280
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11169 7711 11203
rect 21542 11200 21548 11212
rect 21503 11172 21548 11200
rect 7653 11163 7711 11169
rect 21542 11160 21548 11172
rect 21600 11160 21606 11212
rect 24854 11160 24860 11212
rect 24912 11200 24918 11212
rect 25976 11209 26004 11308
rect 26234 11296 26240 11308
rect 26292 11296 26298 11348
rect 36262 11336 36268 11348
rect 36223 11308 36268 11336
rect 36262 11296 36268 11308
rect 36320 11296 36326 11348
rect 38102 11336 38108 11348
rect 38063 11308 38108 11336
rect 38102 11296 38108 11308
rect 38160 11336 38166 11348
rect 39298 11336 39304 11348
rect 38160 11308 39304 11336
rect 38160 11296 38166 11308
rect 39298 11296 39304 11308
rect 39356 11296 39362 11348
rect 29914 11228 29920 11280
rect 29972 11268 29978 11280
rect 30190 11268 30196 11280
rect 29972 11240 30196 11268
rect 29972 11228 29978 11240
rect 30190 11228 30196 11240
rect 30248 11228 30254 11280
rect 39114 11268 39120 11280
rect 38948 11240 39120 11268
rect 25961 11203 26019 11209
rect 25961 11200 25973 11203
rect 24912 11172 25973 11200
rect 24912 11160 24918 11172
rect 25961 11169 25973 11172
rect 26007 11169 26019 11203
rect 25961 11163 26019 11169
rect 32490 11160 32496 11212
rect 32548 11200 32554 11212
rect 32585 11203 32643 11209
rect 32585 11200 32597 11203
rect 32548 11172 32597 11200
rect 32548 11160 32554 11172
rect 32585 11169 32597 11172
rect 32631 11169 32643 11203
rect 32585 11163 32643 11169
rect 32861 11203 32919 11209
rect 32861 11169 32873 11203
rect 32907 11200 32919 11203
rect 33226 11200 33232 11212
rect 32907 11172 33232 11200
rect 32907 11169 32919 11172
rect 32861 11163 32919 11169
rect 33226 11160 33232 11172
rect 33284 11160 33290 11212
rect 34514 11160 34520 11212
rect 34572 11200 34578 11212
rect 34885 11203 34943 11209
rect 34885 11200 34897 11203
rect 34572 11172 34897 11200
rect 34572 11160 34578 11172
rect 34885 11169 34897 11172
rect 34931 11169 34943 11203
rect 38948 11200 38976 11240
rect 39114 11228 39120 11240
rect 39172 11228 39178 11280
rect 40221 11203 40279 11209
rect 40221 11200 40233 11203
rect 38948 11172 39068 11200
rect 34885 11163 34943 11169
rect 7282 11132 7288 11144
rect 7195 11104 7288 11132
rect 7282 11092 7288 11104
rect 7340 11092 7346 11144
rect 7466 11132 7472 11144
rect 7427 11104 7472 11132
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 7834 11132 7840 11144
rect 7795 11104 7840 11132
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 11330 11132 11336 11144
rect 11291 11104 11336 11132
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 21818 11141 21824 11144
rect 21812 11095 21824 11141
rect 21876 11132 21882 11144
rect 21876 11104 21912 11132
rect 21818 11092 21824 11095
rect 21876 11092 21882 11104
rect 23106 11092 23112 11144
rect 23164 11132 23170 11144
rect 23382 11132 23388 11144
rect 23164 11104 23388 11132
rect 23164 11092 23170 11104
rect 23382 11092 23388 11104
rect 23440 11132 23446 11144
rect 23569 11135 23627 11141
rect 23569 11132 23581 11135
rect 23440 11104 23581 11132
rect 23440 11092 23446 11104
rect 23569 11101 23581 11104
rect 23615 11101 23627 11135
rect 23750 11132 23756 11144
rect 23711 11104 23756 11132
rect 23569 11095 23627 11101
rect 23750 11092 23756 11104
rect 23808 11092 23814 11144
rect 24946 11092 24952 11144
rect 25004 11132 25010 11144
rect 25041 11135 25099 11141
rect 25041 11132 25053 11135
rect 25004 11104 25053 11132
rect 25004 11092 25010 11104
rect 25041 11101 25053 11104
rect 25087 11101 25099 11135
rect 25314 11132 25320 11144
rect 25275 11104 25320 11132
rect 25041 11095 25099 11101
rect 25314 11092 25320 11104
rect 25372 11092 25378 11144
rect 30190 11132 30196 11144
rect 30151 11104 30196 11132
rect 30190 11092 30196 11104
rect 30248 11092 30254 11144
rect 30282 11092 30288 11144
rect 30340 11132 30346 11144
rect 30449 11135 30507 11141
rect 30449 11132 30461 11135
rect 30340 11104 30461 11132
rect 30340 11092 30346 11104
rect 30449 11101 30461 11104
rect 30495 11101 30507 11135
rect 30449 11095 30507 11101
rect 37645 11135 37703 11141
rect 37645 11101 37657 11135
rect 37691 11132 37703 11135
rect 38930 11132 38936 11144
rect 37691 11104 38936 11132
rect 37691 11101 37703 11104
rect 37645 11095 37703 11101
rect 38930 11092 38936 11104
rect 38988 11092 38994 11144
rect 39040 11141 39068 11172
rect 39132 11172 40233 11200
rect 39132 11141 39160 11172
rect 40221 11169 40233 11172
rect 40267 11169 40279 11203
rect 40221 11163 40279 11169
rect 39025 11135 39083 11141
rect 39025 11101 39037 11135
rect 39071 11101 39083 11135
rect 39025 11095 39083 11101
rect 39117 11135 39175 11141
rect 39117 11101 39129 11135
rect 39163 11101 39175 11135
rect 39298 11132 39304 11144
rect 39259 11104 39304 11132
rect 39117 11095 39175 11101
rect 39298 11092 39304 11104
rect 39356 11092 39362 11144
rect 40037 11135 40095 11141
rect 40037 11101 40049 11135
rect 40083 11132 40095 11135
rect 40402 11132 40408 11144
rect 40083 11104 40408 11132
rect 40083 11101 40095 11104
rect 40037 11095 40095 11101
rect 40402 11092 40408 11104
rect 40460 11092 40466 11144
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 7006 11064 7012 11076
rect 4856 11036 7012 11064
rect 4856 11024 4862 11036
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7300 11064 7328 11092
rect 8110 11064 8116 11076
rect 7300 11036 8116 11064
rect 8110 11024 8116 11036
rect 8168 11064 8174 11076
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8168 11036 8953 11064
rect 8168 11024 8174 11036
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 14918 11064 14924 11076
rect 9916 11036 14924 11064
rect 9916 11024 9922 11036
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 18141 11067 18199 11073
rect 18141 11033 18153 11067
rect 18187 11064 18199 11067
rect 18230 11064 18236 11076
rect 18187 11036 18236 11064
rect 18187 11033 18199 11036
rect 18141 11027 18199 11033
rect 18230 11024 18236 11036
rect 18288 11064 18294 11076
rect 18782 11064 18788 11076
rect 18288 11036 18788 11064
rect 18288 11024 18294 11036
rect 18782 11024 18788 11036
rect 18840 11024 18846 11076
rect 19150 11024 19156 11076
rect 19208 11064 19214 11076
rect 19429 11067 19487 11073
rect 19429 11064 19441 11067
rect 19208 11036 19441 11064
rect 19208 11024 19214 11036
rect 19429 11033 19441 11036
rect 19475 11064 19487 11067
rect 25590 11064 25596 11076
rect 19475 11036 25596 11064
rect 19475 11033 19487 11036
rect 19429 11027 19487 11033
rect 25590 11024 25596 11036
rect 25648 11024 25654 11076
rect 26234 11073 26240 11076
rect 26228 11027 26240 11073
rect 26292 11064 26298 11076
rect 26292 11036 26328 11064
rect 26234 11024 26240 11027
rect 26292 11024 26298 11036
rect 27706 11024 27712 11076
rect 27764 11064 27770 11076
rect 30006 11064 30012 11076
rect 27764 11036 30012 11064
rect 27764 11024 27770 11036
rect 30006 11024 30012 11036
rect 30064 11024 30070 11076
rect 35158 11073 35164 11076
rect 35152 11027 35164 11073
rect 35216 11064 35222 11076
rect 35216 11036 35252 11064
rect 35158 11024 35164 11027
rect 35216 11024 35222 11036
rect 38286 11024 38292 11076
rect 38344 11064 38350 11076
rect 39853 11067 39911 11073
rect 39853 11064 39865 11067
rect 38344 11036 39865 11064
rect 38344 11024 38350 11036
rect 39853 11033 39865 11036
rect 39899 11033 39911 11067
rect 39853 11027 39911 11033
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 7834 10996 7840 11008
rect 5500 10968 7840 10996
rect 5500 10956 5506 10968
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 22462 10956 22468 11008
rect 22520 10996 22526 11008
rect 22922 10996 22928 11008
rect 22520 10968 22928 10996
rect 22520 10956 22526 10968
rect 22922 10956 22928 10968
rect 22980 10956 22986 11008
rect 23382 10996 23388 11008
rect 23343 10968 23388 10996
rect 23382 10956 23388 10968
rect 23440 10956 23446 11008
rect 27338 10996 27344 11008
rect 27299 10968 27344 10996
rect 27338 10956 27344 10968
rect 27396 10956 27402 11008
rect 28442 10996 28448 11008
rect 28403 10968 28448 10996
rect 28442 10956 28448 10968
rect 28500 10956 28506 11008
rect 31018 10956 31024 11008
rect 31076 10996 31082 11008
rect 31573 10999 31631 11005
rect 31573 10996 31585 10999
rect 31076 10968 31585 10996
rect 31076 10956 31082 10968
rect 31573 10965 31585 10968
rect 31619 10965 31631 10999
rect 38654 10996 38660 11008
rect 38615 10968 38660 10996
rect 31573 10959 31631 10965
rect 38654 10956 38660 10968
rect 38712 10956 38718 11008
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 15654 10752 15660 10804
rect 15712 10792 15718 10804
rect 15930 10792 15936 10804
rect 15712 10764 15936 10792
rect 15712 10752 15718 10764
rect 15930 10752 15936 10764
rect 15988 10752 15994 10804
rect 23293 10795 23351 10801
rect 23293 10792 23305 10795
rect 22066 10764 23305 10792
rect 17034 10724 17040 10736
rect 16995 10696 17040 10724
rect 17034 10684 17040 10696
rect 17092 10684 17098 10736
rect 6638 10656 6644 10668
rect 6599 10628 6644 10656
rect 6638 10616 6644 10628
rect 6696 10616 6702 10668
rect 10594 10656 10600 10668
rect 10555 10628 10600 10656
rect 10594 10616 10600 10628
rect 10652 10656 10658 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 10652 10628 11529 10656
rect 10652 10616 10658 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 15930 10656 15936 10668
rect 15891 10628 15936 10656
rect 11517 10619 11575 10625
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 6365 10591 6423 10597
rect 6365 10557 6377 10591
rect 6411 10588 6423 10591
rect 6730 10588 6736 10600
rect 6411 10560 6736 10588
rect 6411 10557 6423 10560
rect 6365 10551 6423 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 10686 10588 10692 10600
rect 10647 10560 10692 10588
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 13262 10588 13268 10600
rect 10827 10560 13268 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 10796 10520 10824 10551
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 16117 10591 16175 10597
rect 16117 10557 16129 10591
rect 16163 10588 16175 10591
rect 16206 10588 16212 10600
rect 16163 10560 16212 10588
rect 16163 10557 16175 10560
rect 16117 10551 16175 10557
rect 16206 10548 16212 10560
rect 16264 10588 16270 10600
rect 22066 10588 22094 10764
rect 23293 10761 23305 10764
rect 23339 10792 23351 10795
rect 23750 10792 23756 10804
rect 23339 10764 23756 10792
rect 23339 10761 23351 10764
rect 23293 10755 23351 10761
rect 23750 10752 23756 10764
rect 23808 10752 23814 10804
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 25774 10792 25780 10804
rect 24811 10764 25780 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 25869 10795 25927 10801
rect 25869 10761 25881 10795
rect 25915 10792 25927 10795
rect 26234 10792 26240 10804
rect 25915 10764 26240 10792
rect 25915 10761 25927 10764
rect 25869 10755 25927 10761
rect 26234 10752 26240 10764
rect 26292 10752 26298 10804
rect 26418 10752 26424 10804
rect 26476 10792 26482 10804
rect 26476 10764 30374 10792
rect 26476 10752 26482 10764
rect 22278 10684 22284 10736
rect 22336 10724 22342 10736
rect 28442 10724 28448 10736
rect 22336 10696 28448 10724
rect 22336 10684 22342 10696
rect 28442 10684 28448 10696
rect 28500 10724 28506 10736
rect 28629 10727 28687 10733
rect 28629 10724 28641 10727
rect 28500 10696 28641 10724
rect 28500 10684 28506 10696
rect 28629 10693 28641 10696
rect 28675 10693 28687 10727
rect 28629 10687 28687 10693
rect 22462 10656 22468 10668
rect 22423 10628 22468 10656
rect 22462 10616 22468 10628
rect 22520 10616 22526 10668
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10656 22707 10659
rect 23382 10656 23388 10668
rect 22695 10628 23388 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 23382 10616 23388 10628
rect 23440 10656 23446 10668
rect 24397 10659 24455 10665
rect 24397 10656 24409 10659
rect 23440 10628 24409 10656
rect 23440 10616 23446 10628
rect 24397 10625 24409 10628
rect 24443 10625 24455 10659
rect 24397 10619 24455 10625
rect 24581 10659 24639 10665
rect 24581 10625 24593 10659
rect 24627 10656 24639 10659
rect 25038 10656 25044 10668
rect 24627 10628 25044 10656
rect 24627 10625 24639 10628
rect 24581 10619 24639 10625
rect 16264 10560 22094 10588
rect 22281 10591 22339 10597
rect 16264 10548 16270 10560
rect 22281 10557 22293 10591
rect 22327 10588 22339 10591
rect 22554 10588 22560 10600
rect 22327 10560 22560 10588
rect 22327 10557 22339 10560
rect 22281 10551 22339 10557
rect 22554 10548 22560 10560
rect 22612 10548 22618 10600
rect 6236 10492 10824 10520
rect 6236 10480 6242 10492
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 23566 10520 23572 10532
rect 17184 10492 23572 10520
rect 17184 10480 17190 10492
rect 23566 10480 23572 10492
rect 23624 10480 23630 10532
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9824 10424 10241 10452
rect 9824 10412 9830 10424
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 10229 10415 10287 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 19334 10452 19340 10464
rect 19295 10424 19340 10452
rect 19334 10412 19340 10424
rect 19392 10412 19398 10464
rect 24412 10452 24440 10619
rect 25038 10616 25044 10628
rect 25096 10616 25102 10668
rect 25222 10656 25228 10668
rect 25183 10628 25228 10656
rect 25222 10616 25228 10628
rect 25280 10616 25286 10668
rect 25406 10656 25412 10668
rect 25367 10628 25412 10656
rect 25406 10616 25412 10628
rect 25464 10616 25470 10668
rect 25501 10659 25559 10665
rect 25501 10625 25513 10659
rect 25547 10625 25559 10659
rect 25501 10619 25559 10625
rect 24946 10480 24952 10532
rect 25004 10520 25010 10532
rect 25516 10520 25544 10619
rect 25590 10616 25596 10668
rect 25648 10656 25654 10668
rect 27157 10659 27215 10665
rect 25648 10628 25693 10656
rect 25648 10616 25654 10628
rect 27157 10625 27169 10659
rect 27203 10656 27215 10659
rect 27430 10656 27436 10668
rect 27203 10628 27436 10656
rect 27203 10625 27215 10628
rect 27157 10619 27215 10625
rect 27172 10520 27200 10619
rect 27430 10616 27436 10628
rect 27488 10616 27494 10668
rect 27614 10656 27620 10668
rect 27575 10628 27620 10656
rect 27614 10616 27620 10628
rect 27672 10616 27678 10668
rect 27798 10656 27804 10668
rect 27759 10628 27804 10656
rect 27798 10616 27804 10628
rect 27856 10616 27862 10668
rect 27893 10659 27951 10665
rect 27893 10625 27905 10659
rect 27939 10625 27951 10659
rect 27893 10619 27951 10625
rect 27985 10659 28043 10665
rect 27985 10625 27997 10659
rect 28031 10656 28043 10659
rect 28074 10656 28080 10668
rect 28031 10628 28080 10656
rect 28031 10625 28043 10628
rect 27985 10619 28043 10625
rect 27338 10548 27344 10600
rect 27396 10588 27402 10600
rect 27908 10588 27936 10619
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 30346 10656 30374 10764
rect 30558 10752 30564 10804
rect 30616 10792 30622 10804
rect 30837 10795 30895 10801
rect 30837 10792 30849 10795
rect 30616 10764 30849 10792
rect 30616 10752 30622 10764
rect 30837 10761 30849 10764
rect 30883 10761 30895 10795
rect 30837 10755 30895 10761
rect 33962 10752 33968 10804
rect 34020 10792 34026 10804
rect 34517 10795 34575 10801
rect 34517 10792 34529 10795
rect 34020 10764 34529 10792
rect 34020 10752 34026 10764
rect 34517 10761 34529 10764
rect 34563 10761 34575 10795
rect 34517 10755 34575 10761
rect 35069 10795 35127 10801
rect 35069 10761 35081 10795
rect 35115 10792 35127 10795
rect 35158 10792 35164 10804
rect 35115 10764 35164 10792
rect 35115 10761 35127 10764
rect 35069 10755 35127 10761
rect 31018 10724 31024 10736
rect 30979 10696 31024 10724
rect 31018 10684 31024 10696
rect 31076 10684 31082 10736
rect 31205 10727 31263 10733
rect 31205 10693 31217 10727
rect 31251 10724 31263 10727
rect 31294 10724 31300 10736
rect 31251 10696 31300 10724
rect 31251 10693 31263 10696
rect 31205 10687 31263 10693
rect 31294 10684 31300 10696
rect 31352 10724 31358 10736
rect 31662 10724 31668 10736
rect 31352 10696 31668 10724
rect 31352 10684 31358 10696
rect 31662 10684 31668 10696
rect 31720 10684 31726 10736
rect 34532 10724 34560 10755
rect 35158 10752 35164 10764
rect 35216 10752 35222 10804
rect 40129 10795 40187 10801
rect 35452 10764 35756 10792
rect 35452 10724 35480 10764
rect 34532 10696 35480 10724
rect 33965 10659 34023 10665
rect 33965 10656 33977 10659
rect 30346 10628 33977 10656
rect 33965 10625 33977 10628
rect 34011 10656 34023 10659
rect 34790 10656 34796 10668
rect 34011 10628 34796 10656
rect 34011 10625 34023 10628
rect 33965 10619 34023 10625
rect 34790 10616 34796 10628
rect 34848 10656 34854 10668
rect 35728 10665 35756 10764
rect 40129 10761 40141 10795
rect 40175 10792 40187 10795
rect 40402 10792 40408 10804
rect 40175 10764 40408 10792
rect 40175 10761 40187 10764
rect 40129 10755 40187 10761
rect 40402 10752 40408 10764
rect 40460 10752 40466 10804
rect 36262 10684 36268 10736
rect 36320 10724 36326 10736
rect 36357 10727 36415 10733
rect 36357 10724 36369 10727
rect 36320 10696 36369 10724
rect 36320 10684 36326 10696
rect 36357 10693 36369 10696
rect 36403 10693 36415 10727
rect 36357 10687 36415 10693
rect 38654 10684 38660 10736
rect 38712 10724 38718 10736
rect 38994 10727 39052 10733
rect 38994 10724 39006 10727
rect 38712 10696 39006 10724
rect 38712 10684 38718 10696
rect 38994 10693 39006 10696
rect 39040 10693 39052 10727
rect 38994 10687 39052 10693
rect 35345 10659 35403 10665
rect 35345 10656 35357 10659
rect 34848 10628 35357 10656
rect 34848 10616 34854 10628
rect 35345 10625 35357 10628
rect 35391 10625 35403 10659
rect 35345 10619 35403 10625
rect 35434 10659 35492 10665
rect 35434 10625 35446 10659
rect 35480 10625 35492 10659
rect 35434 10619 35492 10625
rect 35529 10659 35587 10665
rect 35529 10625 35541 10659
rect 35575 10656 35587 10659
rect 35713 10659 35771 10665
rect 35575 10628 35664 10656
rect 35575 10625 35587 10628
rect 35529 10619 35587 10625
rect 27396 10560 27936 10588
rect 30285 10591 30343 10597
rect 27396 10548 27402 10560
rect 30285 10557 30297 10591
rect 30331 10588 30343 10591
rect 30466 10588 30472 10600
rect 30331 10560 30472 10588
rect 30331 10557 30343 10560
rect 30285 10551 30343 10557
rect 30466 10548 30472 10560
rect 30524 10548 30530 10600
rect 25004 10492 25544 10520
rect 25608 10492 27200 10520
rect 28169 10523 28227 10529
rect 25004 10480 25010 10492
rect 25608 10452 25636 10492
rect 28169 10489 28181 10523
rect 28215 10520 28227 10523
rect 31202 10520 31208 10532
rect 28215 10492 31208 10520
rect 28215 10489 28227 10492
rect 28169 10483 28227 10489
rect 31202 10480 31208 10492
rect 31260 10480 31266 10532
rect 26970 10452 26976 10464
rect 24412 10424 25636 10452
rect 26931 10424 26976 10452
rect 26970 10412 26976 10424
rect 27028 10412 27034 10464
rect 35452 10452 35480 10619
rect 35636 10588 35664 10628
rect 35713 10625 35725 10659
rect 35759 10625 35771 10659
rect 35713 10619 35771 10625
rect 36541 10659 36599 10665
rect 36541 10625 36553 10659
rect 36587 10656 36599 10659
rect 38286 10656 38292 10668
rect 36587 10628 38292 10656
rect 36587 10625 36599 10628
rect 36541 10619 36599 10625
rect 38286 10616 38292 10628
rect 38344 10616 38350 10668
rect 36173 10591 36231 10597
rect 36173 10588 36185 10591
rect 35636 10560 36185 10588
rect 36173 10557 36185 10560
rect 36219 10557 36231 10591
rect 36173 10551 36231 10557
rect 38378 10548 38384 10600
rect 38436 10588 38442 10600
rect 38749 10591 38807 10597
rect 38749 10588 38761 10591
rect 38436 10560 38761 10588
rect 38436 10548 38442 10560
rect 38749 10557 38761 10560
rect 38795 10557 38807 10591
rect 38749 10551 38807 10557
rect 39114 10452 39120 10464
rect 35452 10424 39120 10452
rect 39114 10412 39120 10424
rect 39172 10412 39178 10464
rect 58158 10452 58164 10464
rect 58119 10424 58164 10452
rect 58158 10412 58164 10424
rect 58216 10412 58222 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 5350 10248 5356 10260
rect 4571 10220 5356 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11054 10248 11060 10260
rect 10919 10220 11060 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11054 10208 11060 10220
rect 11112 10248 11118 10260
rect 13538 10248 13544 10260
rect 11112 10220 13544 10248
rect 11112 10208 11118 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 15838 10208 15844 10260
rect 15896 10248 15902 10260
rect 16301 10251 16359 10257
rect 16301 10248 16313 10251
rect 15896 10220 16313 10248
rect 15896 10208 15902 10220
rect 16301 10217 16313 10220
rect 16347 10217 16359 10251
rect 16301 10211 16359 10217
rect 16945 10251 17003 10257
rect 16945 10217 16957 10251
rect 16991 10248 17003 10251
rect 17034 10248 17040 10260
rect 16991 10220 17040 10248
rect 16991 10217 17003 10220
rect 16945 10211 17003 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 25406 10208 25412 10260
rect 25464 10248 25470 10260
rect 25685 10251 25743 10257
rect 25685 10248 25697 10251
rect 25464 10220 25697 10248
rect 25464 10208 25470 10220
rect 25685 10217 25697 10220
rect 25731 10217 25743 10251
rect 25685 10211 25743 10217
rect 32769 10251 32827 10257
rect 32769 10217 32781 10251
rect 32815 10248 32827 10251
rect 33778 10248 33784 10260
rect 32815 10220 33784 10248
rect 32815 10217 32827 10220
rect 32769 10211 32827 10217
rect 33778 10208 33784 10220
rect 33836 10208 33842 10260
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 12621 10183 12679 10189
rect 12621 10180 12633 10183
rect 12032 10152 12633 10180
rect 12032 10140 12038 10152
rect 12621 10149 12633 10152
rect 12667 10149 12679 10183
rect 12621 10143 12679 10149
rect 12802 10140 12808 10192
rect 12860 10180 12866 10192
rect 14277 10183 14335 10189
rect 14277 10180 14289 10183
rect 12860 10152 14289 10180
rect 12860 10140 12866 10152
rect 14277 10149 14289 10152
rect 14323 10180 14335 10183
rect 14734 10180 14740 10192
rect 14323 10152 14740 10180
rect 14323 10149 14335 10152
rect 14277 10143 14335 10149
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 25133 10183 25191 10189
rect 25133 10149 25145 10183
rect 25179 10180 25191 10183
rect 25590 10180 25596 10192
rect 25179 10152 25596 10180
rect 25179 10149 25191 10152
rect 25133 10143 25191 10149
rect 25590 10140 25596 10152
rect 25648 10140 25654 10192
rect 4062 10072 4068 10124
rect 4120 10112 4126 10124
rect 4522 10112 4528 10124
rect 4120 10084 4528 10112
rect 4120 10072 4126 10084
rect 4522 10072 4528 10084
rect 4580 10112 4586 10124
rect 4580 10084 10640 10112
rect 4580 10072 4586 10084
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 2501 10047 2559 10053
rect 2501 10013 2513 10047
rect 2547 10044 2559 10047
rect 2590 10044 2596 10056
rect 2547 10016 2596 10044
rect 2547 10013 2559 10016
rect 2501 10007 2559 10013
rect 2590 10004 2596 10016
rect 2648 10044 2654 10056
rect 9585 10047 9643 10053
rect 9585 10044 9597 10047
rect 2648 10016 9597 10044
rect 2648 10004 2654 10016
rect 9585 10013 9597 10016
rect 9631 10013 9643 10047
rect 9766 10044 9772 10056
rect 9727 10016 9772 10044
rect 9585 10007 9643 10013
rect 4338 9936 4344 9988
rect 4396 9976 4402 9988
rect 4617 9979 4675 9985
rect 4617 9976 4629 9979
rect 4396 9948 4629 9976
rect 4396 9936 4402 9948
rect 4617 9945 4629 9948
rect 4663 9945 4675 9979
rect 9600 9976 9628 10007
rect 9766 10004 9772 10016
rect 9824 10004 9830 10056
rect 10612 10044 10640 10084
rect 10686 10072 10692 10124
rect 10744 10112 10750 10124
rect 12897 10115 12955 10121
rect 12897 10112 12909 10115
rect 10744 10084 12909 10112
rect 10744 10072 10750 10084
rect 12897 10081 12909 10084
rect 12943 10081 12955 10115
rect 12897 10075 12955 10081
rect 25314 10072 25320 10124
rect 25372 10112 25378 10124
rect 29549 10115 29607 10121
rect 29549 10112 29561 10115
rect 25372 10084 29561 10112
rect 25372 10072 25378 10084
rect 29549 10081 29561 10084
rect 29595 10081 29607 10115
rect 31754 10112 31760 10124
rect 29549 10075 29607 10081
rect 30852 10084 31760 10112
rect 10612 10016 12020 10044
rect 11790 9976 11796 9988
rect 9600 9948 11796 9976
rect 4617 9939 4675 9945
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 1394 9868 1400 9920
rect 1452 9908 1458 9920
rect 2133 9911 2191 9917
rect 2133 9908 2145 9911
rect 1452 9880 2145 9908
rect 1452 9868 1458 9880
rect 2133 9877 2145 9880
rect 2179 9877 2191 9911
rect 6822 9908 6828 9920
rect 6783 9880 6828 9908
rect 2133 9871 2191 9877
rect 6822 9868 6828 9880
rect 6880 9868 6886 9920
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9214 9908 9220 9920
rect 9171 9880 9220 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9214 9868 9220 9880
rect 9272 9908 9278 9920
rect 9398 9908 9404 9920
rect 9272 9880 9404 9908
rect 9272 9868 9278 9880
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9953 9911 10011 9917
rect 9953 9877 9965 9911
rect 9999 9908 10011 9911
rect 11698 9908 11704 9920
rect 9999 9880 11704 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 11992 9908 12020 10016
rect 12526 10004 12532 10056
rect 12584 10044 12590 10056
rect 12805 10047 12863 10053
rect 12805 10044 12817 10047
rect 12584 10016 12817 10044
rect 12584 10004 12590 10016
rect 12805 10013 12817 10016
rect 12851 10013 12863 10047
rect 12805 10007 12863 10013
rect 14921 10047 14979 10053
rect 14921 10013 14933 10047
rect 14967 10044 14979 10047
rect 15838 10044 15844 10056
rect 14967 10016 15844 10044
rect 14967 10013 14979 10016
rect 14921 10007 14979 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 22278 10044 22284 10056
rect 16132 10016 22284 10044
rect 12158 9976 12164 9988
rect 12119 9948 12164 9976
rect 12158 9936 12164 9948
rect 12216 9976 12222 9988
rect 16132 9976 16160 10016
rect 22278 10004 22284 10016
rect 22336 10004 22342 10056
rect 25869 10047 25927 10053
rect 25869 10013 25881 10047
rect 25915 10044 25927 10047
rect 27338 10044 27344 10056
rect 25915 10016 27344 10044
rect 25915 10013 25927 10016
rect 25869 10007 25927 10013
rect 27338 10004 27344 10016
rect 27396 10004 27402 10056
rect 27430 10004 27436 10056
rect 27488 10044 27494 10056
rect 30852 10053 30880 10084
rect 31754 10072 31760 10084
rect 31812 10072 31818 10124
rect 28537 10047 28595 10053
rect 28537 10044 28549 10047
rect 27488 10016 28549 10044
rect 27488 10004 27494 10016
rect 28537 10013 28549 10016
rect 28583 10013 28595 10047
rect 28537 10007 28595 10013
rect 29825 10047 29883 10053
rect 29825 10013 29837 10047
rect 29871 10013 29883 10047
rect 29825 10007 29883 10013
rect 30837 10047 30895 10053
rect 30837 10013 30849 10047
rect 30883 10013 30895 10047
rect 30837 10007 30895 10013
rect 12216 9948 16160 9976
rect 16209 9979 16267 9985
rect 12216 9936 12222 9948
rect 16209 9945 16221 9979
rect 16255 9945 16267 9979
rect 16209 9939 16267 9945
rect 26053 9979 26111 9985
rect 26053 9945 26065 9979
rect 26099 9976 26111 9979
rect 26234 9976 26240 9988
rect 26099 9948 26240 9976
rect 26099 9945 26111 9948
rect 26053 9939 26111 9945
rect 12802 9908 12808 9920
rect 11992 9880 12808 9908
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 13044 9880 13277 9908
rect 13044 9868 13050 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 15378 9908 15384 9920
rect 15339 9880 15384 9908
rect 13265 9871 13323 9877
rect 15378 9868 15384 9880
rect 15436 9868 15442 9920
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 15930 9908 15936 9920
rect 15528 9880 15936 9908
rect 15528 9868 15534 9880
rect 15930 9868 15936 9880
rect 15988 9908 15994 9920
rect 16224 9908 16252 9939
rect 26234 9936 26240 9948
rect 26292 9976 26298 9988
rect 26970 9976 26976 9988
rect 26292 9948 26976 9976
rect 26292 9936 26298 9948
rect 26970 9936 26976 9948
rect 27028 9936 27034 9988
rect 29840 9976 29868 10007
rect 30926 10004 30932 10056
rect 30984 10044 30990 10056
rect 31021 10047 31079 10053
rect 31021 10044 31033 10047
rect 30984 10016 31033 10044
rect 30984 10004 30990 10016
rect 31021 10013 31033 10016
rect 31067 10013 31079 10047
rect 31021 10007 31079 10013
rect 31113 10047 31171 10053
rect 31113 10013 31125 10047
rect 31159 10013 31171 10047
rect 31113 10007 31171 10013
rect 31128 9976 31156 10007
rect 31202 10004 31208 10056
rect 31260 10044 31266 10056
rect 31846 10044 31852 10056
rect 31260 10016 31852 10044
rect 31260 10004 31266 10016
rect 31846 10004 31852 10016
rect 31904 10004 31910 10056
rect 32030 10004 32036 10056
rect 32088 10044 32094 10056
rect 32217 10047 32275 10053
rect 32217 10044 32229 10047
rect 32088 10016 32229 10044
rect 32088 10004 32094 10016
rect 32217 10013 32229 10016
rect 32263 10013 32275 10047
rect 32582 10044 32588 10056
rect 32543 10016 32588 10044
rect 32217 10007 32275 10013
rect 32582 10004 32588 10016
rect 32640 10004 32646 10056
rect 35529 10047 35587 10053
rect 35529 10013 35541 10047
rect 35575 10044 35587 10047
rect 35618 10044 35624 10056
rect 35575 10016 35624 10044
rect 35575 10013 35587 10016
rect 35529 10007 35587 10013
rect 35618 10004 35624 10016
rect 35676 10004 35682 10056
rect 35713 10047 35771 10053
rect 35713 10013 35725 10047
rect 35759 10044 35771 10047
rect 37274 10044 37280 10056
rect 35759 10016 37280 10044
rect 35759 10013 35771 10016
rect 35713 10007 35771 10013
rect 37274 10004 37280 10016
rect 37332 10004 37338 10056
rect 38565 10047 38623 10053
rect 38565 10013 38577 10047
rect 38611 10044 38623 10047
rect 39390 10044 39396 10056
rect 38611 10016 39396 10044
rect 38611 10013 38623 10016
rect 38565 10007 38623 10013
rect 39390 10004 39396 10016
rect 39448 10004 39454 10056
rect 31662 9976 31668 9988
rect 29840 9948 31668 9976
rect 30852 9920 30880 9948
rect 31662 9936 31668 9948
rect 31720 9936 31726 9988
rect 32401 9979 32459 9985
rect 32401 9945 32413 9979
rect 32447 9945 32459 9979
rect 32401 9939 32459 9945
rect 32493 9979 32551 9985
rect 32493 9945 32505 9979
rect 32539 9976 32551 9979
rect 33134 9976 33140 9988
rect 32539 9948 33140 9976
rect 32539 9945 32551 9948
rect 32493 9939 32551 9945
rect 15988 9880 16252 9908
rect 28721 9911 28779 9917
rect 15988 9868 15994 9880
rect 28721 9877 28733 9911
rect 28767 9908 28779 9911
rect 30374 9908 30380 9920
rect 28767 9880 30380 9908
rect 28767 9877 28779 9880
rect 28721 9871 28779 9877
rect 30374 9868 30380 9880
rect 30432 9868 30438 9920
rect 30834 9868 30840 9920
rect 30892 9868 30898 9920
rect 31478 9908 31484 9920
rect 31439 9880 31484 9908
rect 31478 9868 31484 9880
rect 31536 9868 31542 9920
rect 32214 9868 32220 9920
rect 32272 9908 32278 9920
rect 32416 9908 32444 9939
rect 33134 9936 33140 9948
rect 33192 9936 33198 9988
rect 38286 9936 38292 9988
rect 38344 9976 38350 9988
rect 38381 9979 38439 9985
rect 38381 9976 38393 9979
rect 38344 9948 38393 9976
rect 38344 9936 38350 9948
rect 38381 9945 38393 9948
rect 38427 9945 38439 9979
rect 38381 9939 38439 9945
rect 32272 9880 32444 9908
rect 35345 9911 35403 9917
rect 32272 9868 32278 9880
rect 35345 9877 35357 9911
rect 35391 9908 35403 9911
rect 35434 9908 35440 9920
rect 35391 9880 35440 9908
rect 35391 9877 35403 9880
rect 35345 9871 35403 9877
rect 35434 9868 35440 9880
rect 35492 9868 35498 9920
rect 38746 9908 38752 9920
rect 38707 9880 38752 9908
rect 38746 9868 38752 9880
rect 38804 9868 38810 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 9766 9704 9772 9716
rect 9508 9676 9772 9704
rect 8202 9636 8208 9648
rect 4356 9608 8208 9636
rect 4356 9580 4384 9608
rect 8202 9596 8208 9608
rect 8260 9636 8266 9648
rect 8363 9639 8421 9645
rect 8363 9636 8375 9639
rect 8260 9608 8375 9636
rect 8260 9596 8266 9608
rect 8363 9605 8375 9608
rect 8409 9605 8421 9639
rect 8363 9599 8421 9605
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9528 1458 9580
rect 2297 9571 2355 9577
rect 2297 9568 2309 9571
rect 1596 9540 2309 9568
rect 1596 9441 1624 9540
rect 2297 9537 2309 9540
rect 2343 9537 2355 9571
rect 2297 9531 2355 9537
rect 3510 9528 3516 9580
rect 3568 9568 3574 9580
rect 4338 9568 4344 9580
rect 3568 9540 4344 9568
rect 3568 9528 3574 9540
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 5534 9568 5540 9580
rect 5495 9540 5540 9568
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 6730 9528 6736 9580
rect 6788 9568 6794 9580
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6788 9540 6837 9568
rect 6788 9528 6794 9540
rect 6825 9537 6837 9540
rect 6871 9537 6883 9571
rect 6825 9531 6883 9537
rect 8573 9571 8631 9577
rect 8573 9537 8585 9571
rect 8619 9568 8631 9571
rect 9508 9568 9536 9676
rect 9766 9664 9772 9676
rect 9824 9704 9830 9716
rect 10226 9704 10232 9716
rect 9824 9676 10232 9704
rect 9824 9664 9830 9676
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 10965 9707 11023 9713
rect 10965 9704 10977 9707
rect 10744 9676 10977 9704
rect 10744 9664 10750 9676
rect 10965 9673 10977 9676
rect 11011 9673 11023 9707
rect 10965 9667 11023 9673
rect 12158 9664 12164 9716
rect 12216 9704 12222 9716
rect 12253 9707 12311 9713
rect 12253 9704 12265 9707
rect 12216 9676 12265 9704
rect 12216 9664 12222 9676
rect 12253 9673 12265 9676
rect 12299 9673 12311 9707
rect 12253 9667 12311 9673
rect 13538 9664 13544 9716
rect 13596 9704 13602 9716
rect 17034 9704 17040 9716
rect 13596 9676 17040 9704
rect 13596 9664 13602 9676
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 19426 9664 19432 9716
rect 19484 9664 19490 9716
rect 22848 9676 23520 9704
rect 11422 9636 11428 9648
rect 9600 9608 11428 9636
rect 9600 9577 9628 9608
rect 11422 9596 11428 9608
rect 11480 9596 11486 9648
rect 15746 9636 15752 9648
rect 15659 9608 15752 9636
rect 15746 9596 15752 9608
rect 15804 9636 15810 9648
rect 15804 9608 18736 9636
rect 15804 9596 15810 9608
rect 8619 9540 9536 9568
rect 9585 9571 9643 9577
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9852 9571 9910 9577
rect 9852 9537 9864 9571
rect 9898 9568 9910 9571
rect 11698 9568 11704 9580
rect 9898 9540 11560 9568
rect 11659 9540 11704 9568
rect 9898 9537 9910 9540
rect 9852 9531 9910 9537
rect 2038 9500 2044 9512
rect 1999 9472 2044 9500
rect 2038 9460 2044 9472
rect 2096 9460 2102 9512
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 5813 9503 5871 9509
rect 5813 9500 5825 9503
rect 5776 9472 5825 9500
rect 5776 9460 5782 9472
rect 5813 9469 5825 9472
rect 5859 9469 5871 9503
rect 5813 9463 5871 9469
rect 7006 9460 7012 9512
rect 7064 9500 7070 9512
rect 8205 9503 8263 9509
rect 8205 9500 8217 9503
rect 7064 9472 8217 9500
rect 7064 9460 7070 9472
rect 8205 9469 8217 9472
rect 8251 9469 8263 9503
rect 8205 9463 8263 9469
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9401 1639 9435
rect 1581 9395 1639 9401
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 7561 9435 7619 9441
rect 7561 9432 7573 9435
rect 7340 9404 7573 9432
rect 7340 9392 7346 9404
rect 7561 9401 7573 9404
rect 7607 9432 7619 9435
rect 8110 9432 8116 9444
rect 7607 9404 8116 9432
rect 7607 9401 7619 9404
rect 7561 9395 7619 9401
rect 8110 9392 8116 9404
rect 8168 9432 8174 9444
rect 11532 9441 11560 9540
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 11790 9528 11796 9580
rect 11848 9568 11854 9580
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 11848 9540 13185 9568
rect 11848 9528 11854 9540
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13354 9568 13360 9580
rect 13315 9540 13360 9568
rect 13173 9531 13231 9537
rect 13354 9528 13360 9540
rect 13412 9528 13418 9580
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14734 9568 14740 9580
rect 14507 9540 14740 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 11974 9460 11980 9512
rect 12032 9500 12038 9512
rect 15194 9500 15200 9512
rect 12032 9472 15200 9500
rect 12032 9460 12038 9472
rect 15194 9460 15200 9472
rect 15252 9500 15258 9512
rect 15378 9500 15384 9512
rect 15252 9472 15384 9500
rect 15252 9460 15258 9472
rect 15378 9460 15384 9472
rect 15436 9500 15442 9512
rect 15580 9500 15608 9531
rect 15436 9472 15608 9500
rect 15436 9460 15442 9472
rect 15764 9441 15792 9596
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 18472 9540 18613 9568
rect 18472 9528 18478 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 18708 9568 18736 9608
rect 18966 9596 18972 9648
rect 19024 9636 19030 9648
rect 19444 9636 19472 9664
rect 19024 9608 19472 9636
rect 19024 9596 19030 9608
rect 20070 9596 20076 9648
rect 20128 9636 20134 9648
rect 20530 9636 20536 9648
rect 20128 9608 20536 9636
rect 20128 9596 20134 9608
rect 20530 9596 20536 9608
rect 20588 9636 20594 9648
rect 20717 9639 20775 9645
rect 20717 9636 20729 9639
rect 20588 9608 20729 9636
rect 20588 9596 20594 9608
rect 20717 9605 20729 9608
rect 20763 9605 20775 9639
rect 22848 9636 22876 9676
rect 20717 9599 20775 9605
rect 20824 9608 22876 9636
rect 20254 9568 20260 9580
rect 18708 9540 20260 9568
rect 18601 9531 18659 9537
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20824 9500 20852 9608
rect 22922 9596 22928 9648
rect 22980 9636 22986 9648
rect 23385 9639 23443 9645
rect 23385 9636 23397 9639
rect 22980 9608 23397 9636
rect 22980 9596 22986 9608
rect 23385 9605 23397 9608
rect 23431 9605 23443 9639
rect 23492 9636 23520 9676
rect 28534 9664 28540 9716
rect 28592 9704 28598 9716
rect 29178 9704 29184 9716
rect 28592 9676 29184 9704
rect 28592 9664 28598 9676
rect 29178 9664 29184 9676
rect 29236 9664 29242 9716
rect 31018 9664 31024 9716
rect 31076 9704 31082 9716
rect 31076 9676 31340 9704
rect 31076 9664 31082 9676
rect 23566 9636 23572 9648
rect 23492 9608 23572 9636
rect 23385 9599 23443 9605
rect 23566 9596 23572 9608
rect 23624 9636 23630 9648
rect 24762 9636 24768 9648
rect 23624 9608 24768 9636
rect 23624 9596 23630 9608
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 25038 9596 25044 9648
rect 25096 9636 25102 9648
rect 25501 9639 25559 9645
rect 25501 9636 25513 9639
rect 25096 9608 25513 9636
rect 25096 9596 25102 9608
rect 25501 9605 25513 9608
rect 25547 9605 25559 9639
rect 25501 9599 25559 9605
rect 28994 9596 29000 9648
rect 29052 9636 29058 9648
rect 29733 9639 29791 9645
rect 29733 9636 29745 9639
rect 29052 9608 29745 9636
rect 29052 9596 29058 9608
rect 29733 9605 29745 9608
rect 29779 9605 29791 9639
rect 29733 9599 29791 9605
rect 29917 9639 29975 9645
rect 29917 9605 29929 9639
rect 29963 9636 29975 9639
rect 30926 9636 30932 9648
rect 29963 9608 30932 9636
rect 29963 9605 29975 9608
rect 29917 9599 29975 9605
rect 30926 9596 30932 9608
rect 30984 9596 30990 9648
rect 31312 9645 31340 9676
rect 39390 9664 39396 9716
rect 39448 9704 39454 9716
rect 39761 9707 39819 9713
rect 39761 9704 39773 9707
rect 39448 9676 39773 9704
rect 39448 9664 39454 9676
rect 39761 9673 39773 9676
rect 39807 9673 39819 9707
rect 39761 9667 39819 9673
rect 31297 9639 31355 9645
rect 31297 9605 31309 9639
rect 31343 9605 31355 9639
rect 31297 9599 31355 9605
rect 31662 9596 31668 9648
rect 31720 9636 31726 9648
rect 31720 9608 32444 9636
rect 31720 9596 31726 9608
rect 23109 9571 23167 9577
rect 23109 9568 23121 9571
rect 17144 9472 20852 9500
rect 20916 9540 23121 9568
rect 11517 9435 11575 9441
rect 8168 9404 9536 9432
rect 8168 9392 8174 9404
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4433 9367 4491 9373
rect 4433 9364 4445 9367
rect 4028 9336 4445 9364
rect 4028 9324 4034 9336
rect 4433 9333 4445 9336
rect 4479 9364 4491 9367
rect 6178 9364 6184 9376
rect 4479 9336 6184 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6914 9364 6920 9376
rect 6827 9336 6920 9364
rect 6914 9324 6920 9336
rect 6972 9364 6978 9376
rect 7650 9364 7656 9376
rect 6972 9336 7656 9364
rect 6972 9324 6978 9336
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 8757 9367 8815 9373
rect 8757 9333 8769 9367
rect 8803 9364 8815 9367
rect 9398 9364 9404 9376
rect 8803 9336 9404 9364
rect 8803 9333 8815 9336
rect 8757 9327 8815 9333
rect 9398 9324 9404 9336
rect 9456 9324 9462 9376
rect 9508 9364 9536 9404
rect 11517 9401 11529 9435
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 15749 9435 15807 9441
rect 15749 9401 15761 9435
rect 15795 9401 15807 9435
rect 15749 9395 15807 9401
rect 13078 9364 13084 9376
rect 9508 9336 13084 9364
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 13541 9367 13599 9373
rect 13541 9333 13553 9367
rect 13587 9364 13599 9367
rect 14458 9364 14464 9376
rect 13587 9336 14464 9364
rect 13587 9333 13599 9336
rect 13541 9327 13599 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14645 9367 14703 9373
rect 14645 9333 14657 9367
rect 14691 9364 14703 9367
rect 15010 9364 15016 9376
rect 14691 9336 15016 9364
rect 14691 9333 14703 9336
rect 14645 9327 14703 9333
rect 15010 9324 15016 9336
rect 15068 9364 15074 9376
rect 17144 9364 17172 9472
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 20916 9432 20944 9540
rect 23109 9537 23121 9540
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9537 23351 9571
rect 23474 9568 23480 9580
rect 23435 9540 23480 9568
rect 23293 9531 23351 9537
rect 21818 9500 21824 9512
rect 21779 9472 21824 9500
rect 21818 9460 21824 9472
rect 21876 9460 21882 9512
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 20404 9404 20944 9432
rect 22112 9432 22140 9463
rect 22186 9460 22192 9512
rect 22244 9500 22250 9512
rect 23308 9500 23336 9531
rect 23474 9528 23480 9540
rect 23532 9528 23538 9580
rect 25222 9568 25228 9580
rect 25183 9540 25228 9568
rect 25222 9528 25228 9540
rect 25280 9528 25286 9580
rect 25406 9568 25412 9580
rect 25367 9540 25412 9568
rect 25406 9528 25412 9540
rect 25464 9528 25470 9580
rect 25593 9571 25651 9577
rect 25593 9537 25605 9571
rect 25639 9537 25651 9571
rect 25593 9531 25651 9537
rect 22244 9472 23336 9500
rect 23492 9500 23520 9528
rect 25608 9500 25636 9531
rect 28074 9528 28080 9580
rect 28132 9568 28138 9580
rect 28537 9571 28595 9577
rect 28537 9568 28549 9571
rect 28132 9540 28549 9568
rect 28132 9528 28138 9540
rect 28537 9537 28549 9540
rect 28583 9537 28595 9571
rect 28537 9531 28595 9537
rect 29549 9571 29607 9577
rect 29549 9537 29561 9571
rect 29595 9568 29607 9571
rect 30374 9568 30380 9580
rect 29595 9540 30380 9568
rect 29595 9537 29607 9540
rect 29549 9531 29607 9537
rect 28261 9503 28319 9509
rect 28261 9500 28273 9503
rect 23492 9472 28273 9500
rect 22244 9460 22250 9472
rect 23106 9432 23112 9444
rect 22112 9404 23112 9432
rect 20404 9392 20410 9404
rect 23106 9392 23112 9404
rect 23164 9392 23170 9444
rect 15068 9336 17172 9364
rect 18141 9367 18199 9373
rect 15068 9324 15074 9336
rect 18141 9333 18153 9367
rect 18187 9364 18199 9367
rect 18414 9364 18420 9376
rect 18187 9336 18420 9364
rect 18187 9333 18199 9336
rect 18141 9327 18199 9333
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 18782 9364 18788 9376
rect 18743 9336 18788 9364
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 23308 9364 23336 9472
rect 28261 9469 28273 9472
rect 28307 9469 28319 9503
rect 28552 9500 28580 9531
rect 30374 9528 30380 9540
rect 30432 9528 30438 9580
rect 31018 9568 31024 9580
rect 30979 9540 31024 9568
rect 31018 9528 31024 9540
rect 31076 9528 31082 9580
rect 31202 9568 31208 9580
rect 31163 9540 31208 9568
rect 31202 9528 31208 9540
rect 31260 9528 31266 9580
rect 31389 9571 31447 9577
rect 31389 9537 31401 9571
rect 31435 9537 31447 9571
rect 31389 9531 31447 9537
rect 30561 9503 30619 9509
rect 28552 9472 30512 9500
rect 28261 9463 28319 9469
rect 23661 9435 23719 9441
rect 23661 9401 23673 9435
rect 23707 9432 23719 9435
rect 25682 9432 25688 9444
rect 23707 9404 25688 9432
rect 23707 9401 23719 9404
rect 23661 9395 23719 9401
rect 25682 9392 25688 9404
rect 25740 9392 25746 9444
rect 25777 9435 25835 9441
rect 25777 9401 25789 9435
rect 25823 9432 25835 9435
rect 26050 9432 26056 9444
rect 25823 9404 26056 9432
rect 25823 9401 25835 9404
rect 25777 9395 25835 9401
rect 26050 9392 26056 9404
rect 26108 9392 26114 9444
rect 28276 9432 28304 9463
rect 28718 9432 28724 9444
rect 28276 9404 28724 9432
rect 28718 9392 28724 9404
rect 28776 9392 28782 9444
rect 30484 9432 30512 9472
rect 30561 9469 30573 9503
rect 30607 9500 30619 9503
rect 31110 9500 31116 9512
rect 30607 9472 31116 9500
rect 30607 9469 30619 9472
rect 30561 9463 30619 9469
rect 31110 9460 31116 9472
rect 31168 9460 31174 9512
rect 31404 9500 31432 9531
rect 31754 9528 31760 9580
rect 31812 9568 31818 9580
rect 32125 9571 32183 9577
rect 32125 9568 32137 9571
rect 31812 9540 32137 9568
rect 31812 9528 31818 9540
rect 32125 9537 32137 9540
rect 32171 9537 32183 9571
rect 32306 9568 32312 9580
rect 32267 9540 32312 9568
rect 32125 9531 32183 9537
rect 32306 9528 32312 9540
rect 32364 9528 32370 9580
rect 32416 9577 32444 9608
rect 32950 9596 32956 9648
rect 33008 9636 33014 9648
rect 33229 9639 33287 9645
rect 33229 9636 33241 9639
rect 33008 9608 33241 9636
rect 33008 9596 33014 9608
rect 33229 9605 33241 9608
rect 33275 9605 33287 9639
rect 33229 9599 33287 9605
rect 35244 9639 35302 9645
rect 35244 9605 35256 9639
rect 35290 9636 35302 9639
rect 35342 9636 35348 9648
rect 35290 9608 35348 9636
rect 35290 9605 35302 9608
rect 35244 9599 35302 9605
rect 35342 9596 35348 9608
rect 35400 9596 35406 9648
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9537 32459 9571
rect 32401 9531 32459 9537
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9568 32551 9571
rect 32968 9568 32996 9596
rect 38654 9577 38660 9580
rect 32539 9540 32996 9568
rect 32539 9537 32551 9540
rect 32493 9531 32551 9537
rect 38648 9531 38660 9577
rect 38712 9568 38718 9580
rect 38712 9540 38748 9568
rect 38654 9528 38660 9531
rect 38712 9528 38718 9540
rect 32582 9500 32588 9512
rect 31404 9472 32588 9500
rect 31404 9432 31432 9472
rect 32582 9460 32588 9472
rect 32640 9460 32646 9512
rect 34698 9460 34704 9512
rect 34756 9500 34762 9512
rect 34977 9503 35035 9509
rect 34977 9500 34989 9503
rect 34756 9472 34989 9500
rect 34756 9460 34762 9472
rect 34977 9469 34989 9472
rect 35023 9469 35035 9503
rect 34977 9463 35035 9469
rect 37918 9460 37924 9512
rect 37976 9500 37982 9512
rect 38378 9500 38384 9512
rect 37976 9472 38384 9500
rect 37976 9460 37982 9472
rect 38378 9460 38384 9472
rect 38436 9460 38442 9512
rect 31570 9432 31576 9444
rect 30484 9404 31432 9432
rect 31531 9404 31576 9432
rect 31570 9392 31576 9404
rect 31628 9392 31634 9444
rect 25406 9364 25412 9376
rect 23308 9336 25412 9364
rect 25406 9324 25412 9336
rect 25464 9324 25470 9376
rect 30374 9324 30380 9376
rect 30432 9364 30438 9376
rect 31294 9364 31300 9376
rect 30432 9336 31300 9364
rect 30432 9324 30438 9336
rect 31294 9324 31300 9336
rect 31352 9324 31358 9376
rect 32769 9367 32827 9373
rect 32769 9333 32781 9367
rect 32815 9364 32827 9367
rect 33134 9364 33140 9376
rect 32815 9336 33140 9364
rect 32815 9333 32827 9336
rect 32769 9327 32827 9333
rect 33134 9324 33140 9336
rect 33192 9324 33198 9376
rect 35618 9324 35624 9376
rect 35676 9364 35682 9376
rect 36357 9367 36415 9373
rect 36357 9364 36369 9367
rect 35676 9336 36369 9364
rect 35676 9324 35682 9336
rect 36357 9333 36369 9336
rect 36403 9333 36415 9367
rect 36357 9327 36415 9333
rect 37461 9367 37519 9373
rect 37461 9333 37473 9367
rect 37507 9364 37519 9367
rect 37550 9364 37556 9376
rect 37507 9336 37556 9364
rect 37507 9333 37519 9336
rect 37461 9327 37519 9333
rect 37550 9324 37556 9336
rect 37608 9324 37614 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 2409 9163 2467 9169
rect 2409 9160 2421 9163
rect 2372 9132 2421 9160
rect 2372 9120 2378 9132
rect 2409 9129 2421 9132
rect 2455 9129 2467 9163
rect 2409 9123 2467 9129
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 13538 9160 13544 9172
rect 3016 9132 6776 9160
rect 3016 9120 3022 9132
rect 5166 9052 5172 9104
rect 5224 9092 5230 9104
rect 6549 9095 6607 9101
rect 6549 9092 6561 9095
rect 5224 9064 6561 9092
rect 5224 9052 5230 9064
rect 6549 9061 6561 9064
rect 6595 9061 6607 9095
rect 6549 9055 6607 9061
rect 3053 9027 3111 9033
rect 3053 8993 3065 9027
rect 3099 9024 3111 9027
rect 3970 9024 3976 9036
rect 3099 8996 3976 9024
rect 3099 8993 3111 8996
rect 3053 8987 3111 8993
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 5350 9024 5356 9036
rect 5311 8996 5356 9024
rect 5350 8984 5356 8996
rect 5408 8984 5414 9036
rect 5994 9024 6000 9036
rect 5736 8996 6000 9024
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 5534 8956 5540 8968
rect 4295 8928 5540 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 2869 8891 2927 8897
rect 2869 8857 2881 8891
rect 2915 8888 2927 8891
rect 3418 8888 3424 8900
rect 2915 8860 3424 8888
rect 2915 8857 2927 8860
rect 2869 8851 2927 8857
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 4080 8888 4108 8919
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5077 8891 5135 8897
rect 4080 8860 4752 8888
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 2774 8820 2780 8832
rect 1995 8792 2780 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 2774 8780 2780 8792
rect 2832 8820 2838 8832
rect 3881 8823 3939 8829
rect 2832 8792 2877 8820
rect 2832 8780 2838 8792
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 3970 8820 3976 8832
rect 3927 8792 3976 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4724 8829 4752 8860
rect 5077 8857 5089 8891
rect 5123 8888 5135 8891
rect 5626 8888 5632 8900
rect 5123 8860 5632 8888
rect 5123 8857 5135 8860
rect 5077 8851 5135 8857
rect 5626 8848 5632 8860
rect 5684 8888 5690 8900
rect 5736 8888 5764 8996
rect 5994 8984 6000 8996
rect 6052 9024 6058 9036
rect 6178 9024 6184 9036
rect 6052 8996 6184 9024
rect 6052 8984 6058 8996
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 5902 8956 5908 8968
rect 5863 8928 5908 8956
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 6748 8965 6776 9132
rect 10152 9132 13544 9160
rect 8478 9092 8484 9104
rect 6840 9064 8484 9092
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8925 6791 8959
rect 6840 8956 6868 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7190 9024 7196 9036
rect 6963 8996 7196 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7190 8984 7196 8996
rect 7248 9024 7254 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7248 8996 8033 9024
rect 7248 8984 7254 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6840 8928 7021 8956
rect 6733 8919 6791 8925
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7282 8956 7288 8968
rect 7243 8928 7288 8956
rect 7101 8919 7159 8925
rect 5684 8860 5764 8888
rect 5684 8848 5690 8860
rect 5810 8848 5816 8900
rect 5868 8888 5874 8900
rect 7116 8888 7144 8919
rect 7282 8916 7288 8928
rect 7340 8916 7346 8968
rect 10152 8965 10180 9132
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 16022 9160 16028 9172
rect 15528 9132 16028 9160
rect 15528 9120 15534 9132
rect 16022 9120 16028 9132
rect 16080 9160 16086 9172
rect 18693 9163 18751 9169
rect 16080 9132 18644 9160
rect 16080 9120 16086 9132
rect 11422 9092 11428 9104
rect 11383 9064 11428 9092
rect 11422 9052 11428 9064
rect 11480 9052 11486 9104
rect 14093 9095 14151 9101
rect 14093 9061 14105 9095
rect 14139 9061 14151 9095
rect 14093 9055 14151 9061
rect 12526 9024 12532 9036
rect 12487 8996 12532 9024
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 12621 9027 12679 9033
rect 12621 8993 12633 9027
rect 12667 9024 12679 9027
rect 13998 9024 14004 9036
rect 12667 8996 14004 9024
rect 12667 8993 12679 8996
rect 12621 8987 12679 8993
rect 13998 8984 14004 8996
rect 14056 9024 14062 9036
rect 14108 9024 14136 9055
rect 14056 8996 14136 9024
rect 15473 9027 15531 9033
rect 14056 8984 14062 8996
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 18616 9024 18644 9132
rect 18693 9129 18705 9163
rect 18739 9160 18751 9163
rect 19426 9160 19432 9172
rect 18739 9132 19432 9160
rect 18739 9129 18751 9132
rect 18693 9123 18751 9129
rect 19426 9120 19432 9132
rect 19484 9160 19490 9172
rect 20346 9160 20352 9172
rect 19484 9132 20352 9160
rect 19484 9120 19490 9132
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 20622 9160 20628 9172
rect 20535 9132 20628 9160
rect 20622 9120 20628 9132
rect 20680 9160 20686 9172
rect 25222 9160 25228 9172
rect 20680 9132 25228 9160
rect 20680 9120 20686 9132
rect 25222 9120 25228 9132
rect 25280 9120 25286 9172
rect 27706 9160 27712 9172
rect 27667 9132 27712 9160
rect 27706 9120 27712 9132
rect 27764 9120 27770 9172
rect 30098 9160 30104 9172
rect 30059 9132 30104 9160
rect 30098 9120 30104 9132
rect 30156 9120 30162 9172
rect 31665 9163 31723 9169
rect 31665 9129 31677 9163
rect 31711 9160 31723 9163
rect 32306 9160 32312 9172
rect 31711 9132 32312 9160
rect 31711 9129 31723 9132
rect 31665 9123 31723 9129
rect 32306 9120 32312 9132
rect 32364 9120 32370 9172
rect 32677 9163 32735 9169
rect 32677 9129 32689 9163
rect 32723 9160 32735 9163
rect 34238 9160 34244 9172
rect 32723 9132 34244 9160
rect 32723 9129 32735 9132
rect 32677 9123 32735 9129
rect 34238 9120 34244 9132
rect 34296 9120 34302 9172
rect 34977 9163 35035 9169
rect 34977 9129 34989 9163
rect 35023 9160 35035 9163
rect 35342 9160 35348 9172
rect 35023 9132 35348 9160
rect 35023 9129 35035 9132
rect 34977 9123 35035 9129
rect 35342 9120 35348 9132
rect 35400 9120 35406 9172
rect 20254 9052 20260 9104
rect 20312 9092 20318 9104
rect 24486 9092 24492 9104
rect 20312 9064 24492 9092
rect 20312 9052 20318 9064
rect 24486 9052 24492 9064
rect 24544 9052 24550 9104
rect 27798 9092 27804 9104
rect 27448 9064 27804 9092
rect 21177 9027 21235 9033
rect 15519 8996 17356 9024
rect 18616 8996 19380 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 12986 8956 12992 8968
rect 12947 8928 12992 8956
rect 10137 8919 10195 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 17328 8965 17356 8996
rect 16117 8959 16175 8965
rect 16117 8956 16129 8959
rect 14516 8928 16129 8956
rect 14516 8916 14522 8928
rect 16117 8925 16129 8928
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8956 17371 8959
rect 18322 8956 18328 8968
rect 17359 8928 18328 8956
rect 17359 8925 17371 8928
rect 17313 8919 17371 8925
rect 18322 8916 18328 8928
rect 18380 8956 18386 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 18380 8928 19257 8956
rect 18380 8916 18386 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19352 8956 19380 8996
rect 21177 8993 21189 9027
rect 21223 9024 21235 9027
rect 21818 9024 21824 9036
rect 21223 8996 21824 9024
rect 21223 8993 21235 8996
rect 21177 8987 21235 8993
rect 21818 8984 21824 8996
rect 21876 9024 21882 9036
rect 21913 9027 21971 9033
rect 21913 9024 21925 9027
rect 21876 8996 21925 9024
rect 21876 8984 21882 8996
rect 21913 8993 21925 8996
rect 21959 8993 21971 9027
rect 21913 8987 21971 8993
rect 22066 8996 27200 9024
rect 19352 8928 19656 8956
rect 19245 8919 19303 8925
rect 5868 8860 7144 8888
rect 8205 8891 8263 8897
rect 5868 8848 5874 8860
rect 8205 8857 8217 8891
rect 8251 8888 8263 8891
rect 8294 8888 8300 8900
rect 8251 8860 8300 8888
rect 8251 8857 8263 8860
rect 8205 8851 8263 8857
rect 8294 8848 8300 8860
rect 8352 8888 8358 8900
rect 9401 8891 9459 8897
rect 9401 8888 9413 8891
rect 8352 8860 9413 8888
rect 8352 8848 8358 8860
rect 9401 8857 9413 8860
rect 9447 8857 9459 8891
rect 9401 8851 9459 8857
rect 9585 8891 9643 8897
rect 9585 8857 9597 8891
rect 9631 8888 9643 8891
rect 11882 8888 11888 8900
rect 9631 8860 11888 8888
rect 9631 8857 9643 8860
rect 9585 8851 9643 8857
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 15228 8891 15286 8897
rect 15228 8857 15240 8891
rect 15274 8888 15286 8891
rect 15274 8860 15976 8888
rect 15274 8857 15286 8860
rect 15228 8851 15286 8857
rect 4709 8823 4767 8829
rect 4709 8789 4721 8823
rect 4755 8789 4767 8823
rect 4709 8783 4767 8789
rect 5169 8823 5227 8829
rect 5169 8789 5181 8823
rect 5215 8820 5227 8823
rect 5258 8820 5264 8832
rect 5215 8792 5264 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 6086 8820 6092 8832
rect 6047 8792 6092 8820
rect 6086 8780 6092 8792
rect 6144 8780 6150 8832
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 11974 8820 11980 8832
rect 6236 8792 11980 8820
rect 6236 8780 6242 8792
rect 11974 8780 11980 8792
rect 12032 8780 12038 8832
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 15948 8829 15976 8860
rect 17402 8848 17408 8900
rect 17460 8888 17466 8900
rect 17558 8891 17616 8897
rect 17558 8888 17570 8891
rect 17460 8860 17570 8888
rect 17460 8848 17466 8860
rect 17558 8857 17570 8860
rect 17604 8857 17616 8891
rect 17558 8851 17616 8857
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 19490 8891 19548 8897
rect 19490 8888 19502 8891
rect 19116 8860 19502 8888
rect 19116 8848 19122 8860
rect 19490 8857 19502 8860
rect 19536 8857 19548 8891
rect 19628 8888 19656 8928
rect 20530 8916 20536 8968
rect 20588 8956 20594 8968
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 20588 8928 21097 8956
rect 20588 8916 20594 8928
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21266 8956 21272 8968
rect 21227 8928 21272 8956
rect 21085 8919 21143 8925
rect 21266 8916 21272 8928
rect 21324 8916 21330 8968
rect 21358 8916 21364 8968
rect 21416 8956 21422 8968
rect 22066 8956 22094 8996
rect 21416 8928 22094 8956
rect 22189 8959 22247 8965
rect 21416 8916 21422 8928
rect 22189 8925 22201 8959
rect 22235 8956 22247 8959
rect 23474 8956 23480 8968
rect 22235 8928 23480 8956
rect 22235 8925 22247 8928
rect 22189 8919 22247 8925
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 27172 8965 27200 8996
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 27341 8959 27399 8965
rect 27341 8925 27353 8959
rect 27387 8956 27399 8959
rect 27448 8956 27476 9064
rect 27798 9052 27804 9064
rect 27856 9092 27862 9104
rect 27856 9064 31248 9092
rect 27856 9052 27862 9064
rect 28460 9033 28488 9064
rect 31220 9036 31248 9064
rect 35434 9052 35440 9104
rect 35492 9092 35498 9104
rect 35492 9064 35664 9092
rect 35492 9052 35498 9064
rect 28445 9027 28503 9033
rect 28445 8993 28457 9027
rect 28491 8993 28503 9027
rect 28445 8987 28503 8993
rect 28718 8984 28724 9036
rect 28776 9024 28782 9036
rect 28776 8996 29960 9024
rect 28776 8984 28782 8996
rect 27387 8928 27476 8956
rect 27525 8959 27583 8965
rect 27387 8925 27399 8928
rect 27341 8919 27399 8925
rect 27525 8925 27537 8959
rect 27571 8956 27583 8959
rect 28074 8956 28080 8968
rect 27571 8928 28080 8956
rect 27571 8925 27583 8928
rect 27525 8919 27583 8925
rect 28074 8916 28080 8928
rect 28132 8916 28138 8968
rect 28169 8959 28227 8965
rect 28169 8925 28181 8959
rect 28215 8925 28227 8959
rect 28169 8919 28227 8925
rect 24026 8888 24032 8900
rect 19628 8860 24032 8888
rect 19490 8851 19548 8857
rect 24026 8848 24032 8860
rect 24084 8848 24090 8900
rect 25958 8888 25964 8900
rect 24320 8860 25964 8888
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 12216 8792 12357 8820
rect 12216 8780 12222 8792
rect 12345 8789 12357 8792
rect 12391 8789 12403 8823
rect 12345 8783 12403 8789
rect 15933 8823 15991 8829
rect 15933 8789 15945 8823
rect 15979 8789 15991 8823
rect 16574 8820 16580 8832
rect 16535 8792 16580 8820
rect 15933 8783 15991 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 18782 8780 18788 8832
rect 18840 8820 18846 8832
rect 24320 8820 24348 8860
rect 25958 8848 25964 8860
rect 26016 8848 26022 8900
rect 27430 8848 27436 8900
rect 27488 8888 27494 8900
rect 28184 8888 28212 8919
rect 28534 8916 28540 8968
rect 28592 8956 28598 8968
rect 29932 8965 29960 8996
rect 31202 8984 31208 9036
rect 31260 9024 31266 9036
rect 32214 9024 32220 9036
rect 31260 8996 32220 9024
rect 31260 8984 31266 8996
rect 32214 8984 32220 8996
rect 32272 8984 32278 9036
rect 35636 9024 35664 9064
rect 37642 9024 37648 9036
rect 35544 8996 35664 9024
rect 35912 8996 37648 9024
rect 29549 8959 29607 8965
rect 29549 8956 29561 8959
rect 28592 8928 29561 8956
rect 28592 8916 28598 8928
rect 29549 8925 29561 8928
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 29917 8959 29975 8965
rect 29917 8925 29929 8959
rect 29963 8925 29975 8959
rect 31294 8956 31300 8968
rect 31255 8928 31300 8956
rect 29917 8919 29975 8925
rect 31294 8916 31300 8928
rect 31352 8916 31358 8968
rect 32122 8956 32128 8968
rect 32083 8928 32128 8956
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 32398 8956 32404 8968
rect 32359 8928 32404 8956
rect 32398 8916 32404 8928
rect 32456 8916 32462 8968
rect 32493 8959 32551 8965
rect 32493 8925 32505 8959
rect 32539 8956 32551 8959
rect 32582 8956 32588 8968
rect 32539 8928 32588 8956
rect 32539 8925 32551 8928
rect 32493 8919 32551 8925
rect 32582 8916 32588 8928
rect 32640 8916 32646 8968
rect 34790 8916 34796 8968
rect 34848 8956 34854 8968
rect 35207 8959 35265 8965
rect 35207 8956 35219 8959
rect 34848 8928 35219 8956
rect 34848 8916 34854 8928
rect 35207 8925 35219 8928
rect 35253 8925 35265 8959
rect 35207 8919 35265 8925
rect 35358 8956 35416 8962
rect 35358 8922 35370 8956
rect 35404 8922 35416 8956
rect 35358 8916 35416 8922
rect 35458 8956 35516 8962
rect 35458 8922 35470 8956
rect 35504 8953 35516 8956
rect 35544 8953 35572 8996
rect 35504 8925 35572 8953
rect 35504 8922 35516 8925
rect 35458 8916 35516 8922
rect 35618 8916 35624 8968
rect 35676 8956 35682 8968
rect 35802 8956 35808 8968
rect 35676 8928 35808 8956
rect 35676 8916 35682 8928
rect 35802 8916 35808 8928
rect 35860 8916 35866 8968
rect 29733 8891 29791 8897
rect 29733 8888 29745 8891
rect 27488 8860 27533 8888
rect 28092 8860 29745 8888
rect 27488 8848 27494 8860
rect 28092 8832 28120 8860
rect 29733 8857 29745 8860
rect 29779 8857 29791 8891
rect 29733 8851 29791 8857
rect 29825 8891 29883 8897
rect 29825 8857 29837 8891
rect 29871 8857 29883 8891
rect 29825 8851 29883 8857
rect 31481 8891 31539 8897
rect 31481 8857 31493 8891
rect 31527 8888 31539 8891
rect 31570 8888 31576 8900
rect 31527 8860 31576 8888
rect 31527 8857 31539 8860
rect 31481 8851 31539 8857
rect 24486 8820 24492 8832
rect 18840 8792 24348 8820
rect 24447 8792 24492 8820
rect 18840 8780 18846 8792
rect 24486 8780 24492 8792
rect 24544 8780 24550 8832
rect 25406 8780 25412 8832
rect 25464 8820 25470 8832
rect 28074 8820 28080 8832
rect 25464 8792 28080 8820
rect 25464 8780 25470 8792
rect 28074 8780 28080 8792
rect 28132 8780 28138 8832
rect 29840 8820 29868 8851
rect 31496 8820 31524 8851
rect 31570 8848 31576 8860
rect 31628 8848 31634 8900
rect 32214 8848 32220 8900
rect 32272 8888 32278 8900
rect 32309 8891 32367 8897
rect 32309 8888 32321 8891
rect 32272 8860 32321 8888
rect 32272 8848 32278 8860
rect 32309 8857 32321 8860
rect 32355 8857 32367 8891
rect 32309 8851 32367 8857
rect 35373 8888 35401 8916
rect 35912 8888 35940 8996
rect 37642 8984 37648 8996
rect 37700 8984 37706 9036
rect 36906 8956 36912 8968
rect 36867 8928 36912 8956
rect 36906 8916 36912 8928
rect 36964 8916 36970 8968
rect 37550 8956 37556 8968
rect 37511 8928 37556 8956
rect 37550 8916 37556 8928
rect 37608 8916 37614 8968
rect 58158 8956 58164 8968
rect 58119 8928 58164 8956
rect 58158 8916 58164 8928
rect 58216 8916 58222 8968
rect 35373 8860 35940 8888
rect 36725 8891 36783 8897
rect 35373 8832 35401 8860
rect 36725 8857 36737 8891
rect 36771 8888 36783 8891
rect 37274 8888 37280 8900
rect 36771 8860 37280 8888
rect 36771 8857 36783 8860
rect 36725 8851 36783 8857
rect 37274 8848 37280 8860
rect 37332 8848 37338 8900
rect 29840 8792 31524 8820
rect 35342 8780 35348 8832
rect 35400 8780 35406 8832
rect 37090 8820 37096 8832
rect 37051 8792 37096 8820
rect 37090 8780 37096 8792
rect 37148 8780 37154 8832
rect 37918 8780 37924 8832
rect 37976 8820 37982 8832
rect 38841 8823 38899 8829
rect 38841 8820 38853 8823
rect 37976 8792 38853 8820
rect 37976 8780 37982 8792
rect 38841 8789 38853 8792
rect 38887 8789 38899 8823
rect 38841 8783 38899 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 2004 8588 4629 8616
rect 2004 8576 2010 8588
rect 4617 8585 4629 8588
rect 4663 8616 4675 8619
rect 5626 8616 5632 8628
rect 4663 8588 5632 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5810 8616 5816 8628
rect 5771 8588 5816 8616
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 5960 8588 6745 8616
rect 5960 8576 5966 8588
rect 6733 8585 6745 8588
rect 6779 8585 6791 8619
rect 6733 8579 6791 8585
rect 7929 8619 7987 8625
rect 7929 8585 7941 8619
rect 7975 8616 7987 8619
rect 8662 8616 8668 8628
rect 7975 8588 8668 8616
rect 7975 8585 7987 8588
rect 7929 8579 7987 8585
rect 8662 8576 8668 8588
rect 8720 8616 8726 8628
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 8720 8588 9413 8616
rect 8720 8576 8726 8588
rect 9401 8585 9413 8588
rect 9447 8616 9459 8619
rect 9582 8616 9588 8628
rect 9447 8588 9588 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 10321 8619 10379 8625
rect 10321 8616 10333 8619
rect 9732 8588 10333 8616
rect 9732 8576 9738 8588
rect 10321 8585 10333 8588
rect 10367 8616 10379 8619
rect 12986 8616 12992 8628
rect 10367 8588 12992 8616
rect 10367 8585 10379 8588
rect 10321 8579 10379 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13354 8576 13360 8628
rect 13412 8616 13418 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13412 8588 13553 8616
rect 13412 8576 13418 8588
rect 13541 8585 13553 8588
rect 13587 8585 13599 8619
rect 13998 8616 14004 8628
rect 13959 8588 14004 8616
rect 13541 8579 13599 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 15105 8619 15163 8625
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15470 8616 15476 8628
rect 15151 8588 15476 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 17313 8619 17371 8625
rect 17313 8585 17325 8619
rect 17359 8616 17371 8619
rect 17402 8616 17408 8628
rect 17359 8588 17408 8616
rect 17359 8585 17371 8588
rect 17313 8579 17371 8585
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17954 8616 17960 8628
rect 17512 8588 17960 8616
rect 3418 8508 3424 8560
rect 3476 8548 3482 8560
rect 12342 8548 12348 8560
rect 3476 8520 10732 8548
rect 3476 8508 3482 8520
rect 2038 8440 2044 8492
rect 2096 8480 2102 8492
rect 2498 8480 2504 8492
rect 2096 8452 2504 8480
rect 2096 8440 2102 8452
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 2768 8483 2826 8489
rect 2768 8449 2780 8483
rect 2814 8480 2826 8483
rect 3786 8480 3792 8492
rect 2814 8452 3792 8480
rect 2814 8449 2826 8452
rect 2768 8443 2826 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5810 8480 5816 8492
rect 5215 8452 5816 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 8386 8480 8392 8492
rect 7147 8452 8392 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 2038 8344 2044 8356
rect 1999 8316 2044 8344
rect 2038 8304 2044 8316
rect 2096 8304 2102 8356
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 5258 8344 5264 8356
rect 3927 8316 5264 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 5258 8304 5264 8316
rect 5316 8344 5322 8356
rect 5552 8344 5580 8375
rect 5316 8316 5580 8344
rect 5316 8304 5322 8316
rect 5644 8276 5672 8375
rect 6932 8344 6960 8443
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8480 8999 8483
rect 9766 8480 9772 8492
rect 8987 8452 9772 8480
rect 8987 8449 8999 8452
rect 8941 8443 8999 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 10704 8489 10732 8520
rect 10796 8520 12348 8548
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 8018 8412 8024 8424
rect 7979 8384 8024 8412
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8202 8412 8208 8424
rect 8163 8384 8208 8412
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 10796 8421 10824 8520
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 13078 8508 13084 8560
rect 13136 8548 13142 8560
rect 16758 8548 16764 8560
rect 13136 8520 16764 8548
rect 13136 8508 13142 8520
rect 16758 8508 16764 8520
rect 16816 8508 16822 8560
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8480 11759 8483
rect 11790 8480 11796 8492
rect 11747 8452 11796 8480
rect 11747 8449 11759 8452
rect 11701 8443 11759 8449
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 11882 8440 11888 8492
rect 11940 8480 11946 8492
rect 12069 8483 12127 8489
rect 11940 8452 11985 8480
rect 11940 8440 11946 8452
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12618 8480 12624 8492
rect 12299 8452 12624 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 11977 8415 12035 8421
rect 11977 8381 11989 8415
rect 12023 8381 12035 8415
rect 12084 8412 12112 8443
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 13906 8480 13912 8492
rect 13867 8452 13912 8480
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 12084 8384 12296 8412
rect 11977 8375 12035 8381
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 6932 8316 7573 8344
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 7561 8307 7619 8313
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 10796 8344 10824 8375
rect 7708 8316 10824 8344
rect 10965 8347 11023 8353
rect 7708 8304 7714 8316
rect 10965 8313 10977 8347
rect 11011 8344 11023 8347
rect 11992 8344 12020 8375
rect 12268 8356 12296 8384
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 14093 8415 14151 8421
rect 14093 8412 14105 8415
rect 13320 8384 14105 8412
rect 13320 8372 13326 8384
rect 14093 8381 14105 8384
rect 14139 8381 14151 8415
rect 14093 8375 14151 8381
rect 11011 8316 12020 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 12250 8304 12256 8356
rect 12308 8344 12314 8356
rect 12434 8344 12440 8356
rect 12308 8316 12440 8344
rect 12308 8304 12314 8316
rect 12434 8304 12440 8316
rect 12492 8304 12498 8356
rect 12986 8344 12992 8356
rect 12947 8316 12992 8344
rect 12986 8304 12992 8316
rect 13044 8344 13050 8356
rect 14936 8344 14964 8443
rect 16022 8440 16028 8492
rect 16080 8480 16086 8492
rect 17512 8480 17540 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 19058 8616 19064 8628
rect 19019 8588 19064 8616
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 20993 8619 21051 8625
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 21266 8616 21272 8628
rect 21039 8588 21272 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 21266 8576 21272 8588
rect 21324 8576 21330 8628
rect 24486 8576 24492 8628
rect 24544 8616 24550 8628
rect 28902 8616 28908 8628
rect 24544 8588 25912 8616
rect 28863 8588 28908 8616
rect 24544 8576 24550 8588
rect 19521 8551 19579 8557
rect 19521 8548 19533 8551
rect 18616 8520 19533 8548
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 16080 8452 17601 8480
rect 16080 8440 16086 8452
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 17954 8480 17960 8492
rect 17915 8452 17960 8480
rect 17773 8443 17831 8449
rect 13044 8316 14964 8344
rect 17696 8344 17724 8443
rect 17788 8412 17816 8443
rect 17954 8440 17960 8452
rect 18012 8480 18018 8492
rect 18616 8489 18644 8520
rect 19521 8517 19533 8520
rect 19567 8517 19579 8551
rect 19521 8511 19579 8517
rect 19705 8551 19763 8557
rect 19705 8517 19717 8551
rect 19751 8548 19763 8551
rect 20622 8548 20628 8560
rect 19751 8520 20628 8548
rect 19751 8517 19763 8520
rect 19705 8511 19763 8517
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 23692 8551 23750 8557
rect 23692 8517 23704 8551
rect 23738 8548 23750 8551
rect 24397 8551 24455 8557
rect 24397 8548 24409 8551
rect 23738 8520 24409 8548
rect 23738 8517 23750 8520
rect 23692 8511 23750 8517
rect 24397 8517 24409 8520
rect 24443 8517 24455 8551
rect 24397 8511 24455 8517
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 18012 8452 18429 8480
rect 18012 8440 18018 8452
rect 18417 8449 18429 8452
rect 18463 8449 18475 8483
rect 18417 8443 18475 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 18690 8440 18696 8492
rect 18748 8480 18754 8492
rect 18831 8483 18889 8489
rect 18748 8452 18793 8480
rect 18748 8440 18754 8452
rect 18831 8449 18843 8483
rect 18877 8480 18889 8483
rect 18966 8480 18972 8492
rect 18877 8452 18972 8480
rect 18877 8449 18889 8452
rect 18831 8443 18889 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8480 19947 8483
rect 19978 8480 19984 8492
rect 19935 8452 19984 8480
rect 19935 8449 19947 8452
rect 19889 8443 19947 8449
rect 19978 8440 19984 8452
rect 20036 8440 20042 8492
rect 24688 8489 24716 8588
rect 24946 8548 24952 8560
rect 24780 8520 24952 8548
rect 24780 8489 24808 8520
rect 24946 8508 24952 8520
rect 25004 8548 25010 8560
rect 25498 8548 25504 8560
rect 25004 8520 25504 8548
rect 25004 8508 25010 8520
rect 25498 8508 25504 8520
rect 25556 8508 25562 8560
rect 24673 8483 24731 8489
rect 24673 8449 24685 8483
rect 24719 8449 24731 8483
rect 24673 8443 24731 8449
rect 24765 8483 24823 8489
rect 24765 8449 24777 8483
rect 24811 8449 24823 8483
rect 24765 8443 24823 8449
rect 24854 8440 24860 8492
rect 24912 8480 24918 8492
rect 25041 8483 25099 8489
rect 24912 8452 24957 8480
rect 24912 8440 24918 8452
rect 25041 8449 25053 8483
rect 25087 8480 25099 8483
rect 25130 8480 25136 8492
rect 25087 8452 25136 8480
rect 25087 8449 25099 8452
rect 25041 8443 25099 8449
rect 25130 8440 25136 8452
rect 25188 8440 25194 8492
rect 19242 8412 19248 8424
rect 17788 8384 19248 8412
rect 19242 8372 19248 8384
rect 19300 8372 19306 8424
rect 23937 8415 23995 8421
rect 23937 8381 23949 8415
rect 23983 8412 23995 8415
rect 25682 8412 25688 8424
rect 23983 8384 25688 8412
rect 23983 8381 23995 8384
rect 23937 8375 23995 8381
rect 25682 8372 25688 8384
rect 25740 8372 25746 8424
rect 25884 8412 25912 8588
rect 28902 8576 28908 8588
rect 28960 8576 28966 8628
rect 29825 8619 29883 8625
rect 29825 8585 29837 8619
rect 29871 8616 29883 8619
rect 30006 8616 30012 8628
rect 29871 8588 30012 8616
rect 29871 8585 29883 8588
rect 29825 8579 29883 8585
rect 30006 8576 30012 8588
rect 30064 8616 30070 8628
rect 30190 8616 30196 8628
rect 30064 8588 30196 8616
rect 30064 8576 30070 8588
rect 30190 8576 30196 8588
rect 30248 8576 30254 8628
rect 30466 8576 30472 8628
rect 30524 8616 30530 8628
rect 32217 8619 32275 8625
rect 32217 8616 32229 8619
rect 30524 8588 32229 8616
rect 30524 8576 30530 8588
rect 26053 8551 26111 8557
rect 26053 8517 26065 8551
rect 26099 8548 26111 8551
rect 27430 8548 27436 8560
rect 26099 8520 27436 8548
rect 26099 8517 26111 8520
rect 26053 8511 26111 8517
rect 27430 8508 27436 8520
rect 27488 8508 27494 8560
rect 28074 8508 28080 8560
rect 28132 8548 28138 8560
rect 28537 8551 28595 8557
rect 28537 8548 28549 8551
rect 28132 8520 28549 8548
rect 28132 8508 28138 8520
rect 28537 8517 28549 8520
rect 28583 8517 28595 8551
rect 28537 8511 28595 8517
rect 28629 8551 28687 8557
rect 28629 8517 28641 8551
rect 28675 8548 28687 8551
rect 28994 8548 29000 8560
rect 28675 8520 29000 8548
rect 28675 8517 28687 8520
rect 28629 8511 28687 8517
rect 28994 8508 29000 8520
rect 29052 8508 29058 8560
rect 31128 8492 31156 8588
rect 32217 8585 32229 8588
rect 32263 8616 32275 8619
rect 37550 8616 37556 8628
rect 32263 8588 37556 8616
rect 32263 8585 32275 8588
rect 32217 8579 32275 8585
rect 37550 8576 37556 8588
rect 37608 8576 37614 8628
rect 38565 8619 38623 8625
rect 38565 8585 38577 8619
rect 38611 8616 38623 8619
rect 38654 8616 38660 8628
rect 38611 8588 38660 8616
rect 38611 8585 38623 8588
rect 38565 8579 38623 8585
rect 38654 8576 38660 8588
rect 38712 8576 38718 8628
rect 34790 8548 34796 8560
rect 34751 8520 34796 8548
rect 34790 8508 34796 8520
rect 34848 8508 34854 8560
rect 37090 8508 37096 8560
rect 37148 8548 37154 8560
rect 37148 8520 37667 8548
rect 37148 8508 37154 8520
rect 37639 8492 37667 8520
rect 38746 8508 38752 8560
rect 38804 8548 38810 8560
rect 38804 8520 39068 8548
rect 38804 8508 38810 8520
rect 26234 8480 26240 8492
rect 26195 8452 26240 8480
rect 26234 8440 26240 8452
rect 26292 8440 26298 8492
rect 28350 8480 28356 8492
rect 28311 8452 28356 8480
rect 28350 8440 28356 8452
rect 28408 8440 28414 8492
rect 28718 8480 28724 8492
rect 28679 8452 28724 8480
rect 28718 8440 28724 8452
rect 28776 8440 28782 8492
rect 31110 8480 31116 8492
rect 31071 8452 31116 8480
rect 31110 8440 31116 8452
rect 31168 8440 31174 8492
rect 36633 8483 36691 8489
rect 36633 8480 36645 8483
rect 32232 8452 36645 8480
rect 26418 8412 26424 8424
rect 25884 8384 26424 8412
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 18690 8344 18696 8356
rect 17696 8316 18696 8344
rect 13044 8304 13050 8316
rect 18690 8304 18696 8316
rect 18748 8304 18754 8356
rect 25958 8304 25964 8356
rect 26016 8344 26022 8356
rect 29546 8344 29552 8356
rect 26016 8316 29552 8344
rect 26016 8304 26022 8316
rect 29546 8304 29552 8316
rect 29604 8344 29610 8356
rect 32232 8344 32260 8452
rect 36633 8449 36645 8452
rect 36679 8480 36691 8483
rect 37274 8480 37280 8492
rect 36679 8452 37280 8480
rect 36679 8449 36691 8452
rect 36633 8443 36691 8449
rect 37274 8440 37280 8452
rect 37332 8440 37338 8492
rect 37461 8483 37519 8489
rect 37461 8449 37473 8483
rect 37507 8449 37519 8483
rect 37461 8443 37519 8449
rect 37624 8486 37682 8492
rect 37624 8452 37636 8486
rect 37670 8452 37682 8486
rect 37624 8446 37682 8452
rect 35526 8372 35532 8424
rect 35584 8412 35590 8424
rect 37476 8412 37504 8443
rect 37734 8440 37740 8492
rect 37792 8480 37798 8492
rect 37875 8483 37933 8489
rect 37792 8452 37837 8480
rect 37792 8440 37798 8452
rect 37875 8449 37887 8483
rect 37921 8480 37933 8483
rect 38838 8480 38844 8492
rect 37921 8452 38844 8480
rect 37921 8449 37933 8452
rect 37875 8443 37933 8449
rect 38838 8440 38844 8452
rect 38896 8440 38902 8492
rect 39040 8489 39068 8520
rect 38933 8483 38991 8489
rect 38933 8449 38945 8483
rect 38979 8449 38991 8483
rect 38933 8443 38991 8449
rect 39025 8483 39083 8489
rect 39025 8449 39037 8483
rect 39071 8449 39083 8483
rect 39025 8443 39083 8449
rect 39209 8483 39267 8489
rect 39209 8449 39221 8483
rect 39255 8480 39267 8483
rect 39298 8480 39304 8492
rect 39255 8452 39304 8480
rect 39255 8449 39267 8452
rect 39209 8443 39267 8449
rect 35584 8384 37504 8412
rect 35584 8372 35590 8384
rect 38654 8372 38660 8424
rect 38712 8412 38718 8424
rect 38948 8412 38976 8443
rect 39114 8412 39120 8424
rect 38712 8384 39120 8412
rect 38712 8372 38718 8384
rect 39114 8372 39120 8384
rect 39172 8372 39178 8424
rect 29604 8316 32260 8344
rect 29604 8304 29610 8316
rect 34698 8304 34704 8356
rect 34756 8344 34762 8356
rect 37918 8344 37924 8356
rect 34756 8316 37924 8344
rect 34756 8304 34762 8316
rect 37918 8304 37924 8316
rect 37976 8304 37982 8356
rect 39224 8344 39252 8443
rect 39298 8440 39304 8452
rect 39356 8480 39362 8492
rect 39669 8483 39727 8489
rect 39669 8480 39681 8483
rect 39356 8452 39681 8480
rect 39356 8440 39362 8452
rect 39669 8449 39681 8452
rect 39715 8449 39727 8483
rect 39669 8443 39727 8449
rect 38028 8316 39252 8344
rect 6730 8276 6736 8288
rect 5644 8248 6736 8276
rect 6730 8236 6736 8248
rect 6788 8276 6794 8288
rect 6914 8276 6920 8288
rect 6788 8248 6920 8276
rect 6788 8236 6794 8248
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 11514 8276 11520 8288
rect 11475 8248 11520 8276
rect 11514 8236 11520 8248
rect 11572 8236 11578 8288
rect 16022 8276 16028 8288
rect 15983 8248 16028 8276
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 17678 8236 17684 8288
rect 17736 8276 17742 8288
rect 18966 8276 18972 8288
rect 17736 8248 18972 8276
rect 17736 8236 17742 8248
rect 18966 8236 18972 8248
rect 19024 8236 19030 8288
rect 22557 8279 22615 8285
rect 22557 8245 22569 8279
rect 22603 8276 22615 8279
rect 22922 8276 22928 8288
rect 22603 8248 22928 8276
rect 22603 8245 22615 8248
rect 22557 8239 22615 8245
rect 22922 8236 22928 8248
rect 22980 8236 22986 8288
rect 25590 8236 25596 8288
rect 25648 8276 25654 8288
rect 25869 8279 25927 8285
rect 25869 8276 25881 8279
rect 25648 8248 25881 8276
rect 25648 8236 25654 8248
rect 25869 8245 25881 8248
rect 25915 8245 25927 8279
rect 25869 8239 25927 8245
rect 36078 8236 36084 8288
rect 36136 8276 36142 8288
rect 38028 8276 38056 8316
rect 36136 8248 38056 8276
rect 38105 8279 38163 8285
rect 36136 8236 36142 8248
rect 38105 8245 38117 8279
rect 38151 8276 38163 8279
rect 38194 8276 38200 8288
rect 38151 8248 38200 8276
rect 38151 8245 38163 8248
rect 38105 8239 38163 8245
rect 38194 8236 38200 8248
rect 38252 8236 38258 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 7466 8072 7472 8084
rect 4939 8044 7472 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 7837 8075 7895 8081
rect 7837 8041 7849 8075
rect 7883 8072 7895 8075
rect 8018 8072 8024 8084
rect 7883 8044 8024 8072
rect 7883 8041 7895 8044
rect 7837 8035 7895 8041
rect 8018 8032 8024 8044
rect 8076 8032 8082 8084
rect 17678 8072 17684 8084
rect 9140 8044 12434 8072
rect 17639 8044 17684 8072
rect 2498 7896 2504 7948
rect 2556 7936 2562 7948
rect 6457 7939 6515 7945
rect 6457 7936 6469 7939
rect 2556 7908 6469 7936
rect 2556 7896 2562 7908
rect 6457 7905 6469 7908
rect 6503 7905 6515 7939
rect 6457 7899 6515 7905
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 6713 7871 6771 7877
rect 6713 7868 6725 7871
rect 6144 7840 6725 7868
rect 6144 7828 6150 7840
rect 6713 7837 6725 7840
rect 6759 7837 6771 7871
rect 6713 7831 6771 7837
rect 7006 7828 7012 7880
rect 7064 7868 7070 7880
rect 9140 7868 9168 8044
rect 12406 8004 12434 8044
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 18012 8044 18245 8072
rect 18012 8032 18018 8044
rect 18233 8041 18245 8044
rect 18279 8041 18291 8075
rect 19242 8072 19248 8084
rect 19203 8044 19248 8072
rect 18233 8035 18291 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 23198 8072 23204 8084
rect 23159 8044 23204 8072
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 24765 8075 24823 8081
rect 24765 8041 24777 8075
rect 24811 8072 24823 8075
rect 24854 8072 24860 8084
rect 24811 8044 24860 8072
rect 24811 8041 24823 8044
rect 24765 8035 24823 8041
rect 24854 8032 24860 8044
rect 24912 8032 24918 8084
rect 27065 8075 27123 8081
rect 24964 8044 26648 8072
rect 12406 7976 14596 8004
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12437 7939 12495 7945
rect 12437 7936 12449 7939
rect 11940 7908 12449 7936
rect 11940 7896 11946 7908
rect 12437 7905 12449 7908
rect 12483 7905 12495 7939
rect 13446 7936 13452 7948
rect 12437 7899 12495 7905
rect 12636 7908 13452 7936
rect 7064 7840 9168 7868
rect 10229 7871 10287 7877
rect 7064 7828 7070 7840
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 11422 7868 11428 7880
rect 10275 7840 11428 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 11698 7828 11704 7880
rect 11756 7868 11762 7880
rect 12636 7877 12664 7908
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 14568 7877 14596 7976
rect 16850 7964 16856 8016
rect 16908 8004 16914 8016
rect 16945 8007 17003 8013
rect 16945 8004 16957 8007
rect 16908 7976 16957 8004
rect 16908 7964 16914 7976
rect 16945 7973 16957 7976
rect 16991 8004 17003 8007
rect 16991 7976 22692 8004
rect 16991 7973 17003 7976
rect 16945 7967 17003 7973
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 18748 7908 21128 7936
rect 18748 7896 18754 7908
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 11756 7840 12265 7868
rect 11756 7828 11762 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 12520 7871 12578 7877
rect 12520 7868 12532 7871
rect 12253 7831 12311 7837
rect 12452 7840 12532 7868
rect 2133 7803 2191 7809
rect 2133 7769 2145 7803
rect 2179 7800 2191 7803
rect 3050 7800 3056 7812
rect 2179 7772 3056 7800
rect 2179 7769 2191 7772
rect 2133 7763 2191 7769
rect 3050 7760 3056 7772
rect 3108 7760 3114 7812
rect 5445 7803 5503 7809
rect 5445 7769 5457 7803
rect 5491 7800 5503 7803
rect 6362 7800 6368 7812
rect 5491 7772 6368 7800
rect 5491 7769 5503 7772
rect 5445 7763 5503 7769
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 7282 7760 7288 7812
rect 7340 7800 7346 7812
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 7340 7772 9505 7800
rect 7340 7760 7346 7772
rect 9493 7769 9505 7772
rect 9539 7769 9551 7803
rect 9493 7763 9551 7769
rect 10496 7803 10554 7809
rect 10496 7769 10508 7803
rect 10542 7800 10554 7803
rect 11514 7800 11520 7812
rect 10542 7772 11520 7800
rect 10542 7769 10554 7772
rect 10496 7763 10554 7769
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 12158 7760 12164 7812
rect 12216 7800 12222 7812
rect 12452 7800 12480 7840
rect 12520 7837 12532 7840
rect 12566 7837 12578 7871
rect 12520 7831 12578 7837
rect 12617 7871 12675 7877
rect 12617 7837 12629 7871
rect 12663 7837 12675 7871
rect 12617 7831 12675 7837
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15286 7868 15292 7880
rect 14599 7840 15292 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 12820 7800 12848 7831
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15562 7868 15568 7880
rect 15523 7840 15568 7868
rect 15562 7828 15568 7840
rect 15620 7828 15626 7880
rect 19426 7868 19432 7880
rect 19387 7840 19432 7868
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 19536 7840 21005 7868
rect 12216 7772 12480 7800
rect 12636 7772 12848 7800
rect 12216 7760 12222 7772
rect 12636 7744 12664 7772
rect 15378 7760 15384 7812
rect 15436 7800 15442 7812
rect 15810 7803 15868 7809
rect 15810 7800 15822 7803
rect 15436 7772 15822 7800
rect 15436 7760 15442 7772
rect 15810 7769 15822 7772
rect 15856 7769 15868 7803
rect 19536 7800 19564 7840
rect 20993 7837 21005 7840
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 15810 7763 15868 7769
rect 17604 7772 19564 7800
rect 19613 7803 19671 7809
rect 2682 7732 2688 7744
rect 2643 7704 2688 7732
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3694 7732 3700 7744
rect 3283 7704 3700 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3694 7692 3700 7704
rect 3752 7692 3758 7744
rect 5997 7735 6055 7741
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 7190 7732 7196 7744
rect 6043 7704 7196 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 7190 7692 7196 7704
rect 7248 7692 7254 7744
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8720 7704 8953 7732
rect 8720 7692 8726 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 11609 7735 11667 7741
rect 11609 7701 11621 7735
rect 11655 7732 11667 7735
rect 11790 7732 11796 7744
rect 11655 7704 11796 7732
rect 11655 7701 11667 7704
rect 11609 7695 11667 7701
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12069 7735 12127 7741
rect 12069 7701 12081 7735
rect 12115 7732 12127 7735
rect 12526 7732 12532 7744
rect 12115 7704 12532 7732
rect 12115 7701 12127 7704
rect 12069 7695 12127 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 12618 7692 12624 7744
rect 12676 7692 12682 7744
rect 13449 7735 13507 7741
rect 13449 7701 13461 7735
rect 13495 7732 13507 7735
rect 13538 7732 13544 7744
rect 13495 7704 13544 7732
rect 13495 7701 13507 7704
rect 13449 7695 13507 7701
rect 13538 7692 13544 7704
rect 13596 7732 13602 7744
rect 13906 7732 13912 7744
rect 13596 7704 13912 7732
rect 13596 7692 13602 7704
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 17604 7732 17632 7772
rect 19613 7769 19625 7803
rect 19659 7800 19671 7803
rect 19978 7800 19984 7812
rect 19659 7772 19984 7800
rect 19659 7769 19671 7772
rect 19613 7763 19671 7769
rect 19978 7760 19984 7772
rect 20036 7760 20042 7812
rect 14691 7704 17632 7732
rect 21008 7732 21036 7831
rect 21100 7809 21128 7908
rect 22664 7877 22692 7976
rect 24118 7964 24124 8016
rect 24176 8004 24182 8016
rect 24964 8004 24992 8044
rect 24176 7976 24992 8004
rect 26620 8004 26648 8044
rect 27065 8041 27077 8075
rect 27111 8072 27123 8075
rect 27430 8072 27436 8084
rect 27111 8044 27436 8072
rect 27111 8041 27123 8044
rect 27065 8035 27123 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 28994 8032 29000 8084
rect 29052 8072 29058 8084
rect 30193 8075 30251 8081
rect 30193 8072 30205 8075
rect 29052 8044 30205 8072
rect 29052 8032 29058 8044
rect 30193 8041 30205 8044
rect 30239 8041 30251 8075
rect 34977 8075 35035 8081
rect 34977 8072 34989 8075
rect 30193 8035 30251 8041
rect 30300 8044 34989 8072
rect 30300 8004 30328 8044
rect 34977 8041 34989 8044
rect 35023 8041 35035 8075
rect 36078 8072 36084 8084
rect 36039 8044 36084 8072
rect 34977 8035 35035 8041
rect 36078 8032 36084 8044
rect 36136 8032 36142 8084
rect 37274 8072 37280 8084
rect 37235 8044 37280 8072
rect 37274 8032 37280 8044
rect 37332 8032 37338 8084
rect 39301 8075 39359 8081
rect 39301 8072 39313 8075
rect 37752 8044 39313 8072
rect 26620 7976 30328 8004
rect 24176 7964 24182 7976
rect 36906 7964 36912 8016
rect 36964 8004 36970 8016
rect 37752 8004 37780 8044
rect 39301 8041 39313 8044
rect 39347 8041 39359 8075
rect 39301 8035 39359 8041
rect 36964 7976 37780 8004
rect 36964 7964 36970 7976
rect 25682 7936 25688 7948
rect 22940 7908 24624 7936
rect 25643 7908 25688 7936
rect 22940 7880 22968 7908
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 22649 7871 22707 7877
rect 21223 7840 22600 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 22572 7812 22600 7840
rect 22649 7837 22661 7871
rect 22695 7837 22707 7871
rect 22922 7868 22928 7880
rect 22883 7840 22928 7868
rect 22649 7831 22707 7837
rect 22922 7828 22928 7840
rect 22980 7828 22986 7880
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7868 23075 7871
rect 23198 7868 23204 7880
rect 23063 7840 23204 7868
rect 23063 7837 23075 7840
rect 23017 7831 23075 7837
rect 23198 7828 23204 7840
rect 23256 7828 23262 7880
rect 24596 7877 24624 7908
rect 25682 7896 25688 7908
rect 25740 7896 25746 7948
rect 37918 7936 37924 7948
rect 35268 7908 37780 7936
rect 37879 7908 37924 7936
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7837 24639 7871
rect 26234 7868 26240 7880
rect 24581 7831 24639 7837
rect 25424 7840 26240 7868
rect 21085 7803 21143 7809
rect 21085 7769 21097 7803
rect 21131 7800 21143 7803
rect 21131 7772 22094 7800
rect 21131 7769 21143 7772
rect 21085 7763 21143 7769
rect 21637 7735 21695 7741
rect 21637 7732 21649 7735
rect 21008 7704 21649 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 21637 7701 21649 7704
rect 21683 7732 21695 7735
rect 21726 7732 21732 7744
rect 21683 7704 21732 7732
rect 21683 7701 21695 7704
rect 21637 7695 21695 7701
rect 21726 7692 21732 7704
rect 21784 7692 21790 7744
rect 22066 7732 22094 7772
rect 22554 7760 22560 7812
rect 22612 7800 22618 7812
rect 22833 7803 22891 7809
rect 22833 7800 22845 7803
rect 22612 7772 22845 7800
rect 22612 7760 22618 7772
rect 22833 7769 22845 7772
rect 22879 7769 22891 7803
rect 22833 7763 22891 7769
rect 24302 7760 24308 7812
rect 24360 7800 24366 7812
rect 24397 7803 24455 7809
rect 24397 7800 24409 7803
rect 24360 7772 24409 7800
rect 24360 7760 24366 7772
rect 24397 7769 24409 7772
rect 24443 7800 24455 7803
rect 25424 7800 25452 7840
rect 26234 7828 26240 7840
rect 26292 7828 26298 7880
rect 31317 7871 31375 7877
rect 31317 7837 31329 7871
rect 31363 7868 31375 7871
rect 31478 7868 31484 7880
rect 31363 7840 31484 7868
rect 31363 7837 31375 7840
rect 31317 7831 31375 7837
rect 31478 7828 31484 7840
rect 31536 7828 31542 7880
rect 31573 7871 31631 7877
rect 31573 7837 31585 7871
rect 31619 7868 31631 7871
rect 33870 7868 33876 7880
rect 31619 7840 33876 7868
rect 31619 7837 31631 7840
rect 31573 7831 31631 7837
rect 33870 7828 33876 7840
rect 33928 7828 33934 7880
rect 35268 7877 35296 7908
rect 35161 7871 35219 7877
rect 35161 7837 35173 7871
rect 35207 7837 35219 7871
rect 35161 7831 35219 7837
rect 35253 7871 35311 7877
rect 35253 7837 35265 7871
rect 35299 7837 35311 7871
rect 35253 7831 35311 7837
rect 35529 7871 35587 7877
rect 35529 7837 35541 7871
rect 35575 7868 35587 7871
rect 35618 7868 35624 7880
rect 35575 7840 35624 7868
rect 35575 7837 35587 7840
rect 35529 7831 35587 7837
rect 24443 7772 25452 7800
rect 25952 7803 26010 7809
rect 24443 7769 24455 7772
rect 24397 7763 24455 7769
rect 25952 7769 25964 7803
rect 25998 7800 26010 7803
rect 26050 7800 26056 7812
rect 25998 7772 26056 7800
rect 25998 7769 26010 7772
rect 25952 7763 26010 7769
rect 26050 7760 26056 7772
rect 26108 7760 26114 7812
rect 25774 7732 25780 7744
rect 22066 7704 25780 7732
rect 25774 7692 25780 7704
rect 25832 7692 25838 7744
rect 35176 7732 35204 7831
rect 35618 7828 35624 7840
rect 35676 7828 35682 7880
rect 35345 7803 35403 7809
rect 35345 7769 35357 7803
rect 35391 7800 35403 7803
rect 35434 7800 35440 7812
rect 35391 7772 35440 7800
rect 35391 7769 35403 7772
rect 35345 7763 35403 7769
rect 35434 7760 35440 7772
rect 35492 7760 35498 7812
rect 37752 7800 37780 7908
rect 37918 7896 37924 7908
rect 37976 7896 37982 7948
rect 38194 7877 38200 7880
rect 38188 7868 38200 7877
rect 38155 7840 38200 7868
rect 38188 7831 38200 7840
rect 38194 7828 38200 7831
rect 38252 7828 38258 7880
rect 58158 7868 58164 7880
rect 58119 7840 58164 7868
rect 58158 7828 58164 7840
rect 58216 7828 58222 7880
rect 38838 7800 38844 7812
rect 37752 7772 38844 7800
rect 38838 7760 38844 7772
rect 38896 7760 38902 7812
rect 35710 7732 35716 7744
rect 35176 7704 35716 7732
rect 35710 7692 35716 7704
rect 35768 7692 35774 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 3878 7528 3884 7540
rect 3839 7500 3884 7528
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 6840 7500 7757 7528
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5718 7392 5724 7404
rect 5583 7364 5724 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5718 7352 5724 7364
rect 5776 7392 5782 7404
rect 6840 7392 6868 7500
rect 7745 7497 7757 7500
rect 7791 7528 7803 7531
rect 9674 7528 9680 7540
rect 7791 7500 9680 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 9858 7528 9864 7540
rect 9819 7500 9864 7528
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 11701 7531 11759 7537
rect 11701 7528 11713 7531
rect 10980 7500 11713 7528
rect 6914 7420 6920 7472
rect 6972 7460 6978 7472
rect 6972 7432 8248 7460
rect 6972 7420 6978 7432
rect 5776 7364 6868 7392
rect 5776 7352 5782 7364
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8220 7401 8248 7432
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 10873 7463 10931 7469
rect 10873 7460 10885 7463
rect 9824 7432 10885 7460
rect 9824 7420 9830 7432
rect 10873 7429 10885 7432
rect 10919 7429 10931 7463
rect 10873 7423 10931 7429
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 8076 7364 8125 7392
rect 8076 7352 8082 7364
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 10980 7392 11008 7500
rect 11701 7497 11713 7500
rect 11747 7528 11759 7531
rect 11882 7528 11888 7540
rect 11747 7500 11888 7528
rect 11747 7497 11759 7500
rect 11701 7491 11759 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 15197 7531 15255 7537
rect 12492 7500 12537 7528
rect 12492 7488 12498 7500
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15654 7528 15660 7540
rect 15243 7500 15660 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15654 7488 15660 7500
rect 15712 7528 15718 7540
rect 20349 7531 20407 7537
rect 20349 7528 20361 7531
rect 15712 7500 20361 7528
rect 15712 7488 15718 7500
rect 20349 7497 20361 7500
rect 20395 7528 20407 7531
rect 22925 7531 22983 7537
rect 20395 7500 20944 7528
rect 20395 7497 20407 7500
rect 20349 7491 20407 7497
rect 15105 7463 15163 7469
rect 15105 7429 15117 7463
rect 15151 7460 15163 7463
rect 15286 7460 15292 7472
rect 15151 7432 15292 7460
rect 15151 7429 15163 7432
rect 15105 7423 15163 7429
rect 15286 7420 15292 7432
rect 15344 7420 15350 7472
rect 16850 7460 16856 7472
rect 16811 7432 16856 7460
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 17310 7420 17316 7472
rect 17368 7460 17374 7472
rect 17368 7432 19656 7460
rect 17368 7420 17374 7432
rect 8444 7364 11008 7392
rect 11517 7395 11575 7401
rect 8444 7352 8450 7364
rect 11517 7361 11529 7395
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 5626 7324 5632 7336
rect 2363 7296 5632 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 5810 7324 5816 7336
rect 5771 7296 5816 7324
rect 5810 7284 5816 7296
rect 5868 7284 5874 7336
rect 6454 7324 6460 7336
rect 6415 7296 6460 7324
rect 6454 7284 6460 7296
rect 6512 7284 6518 7336
rect 6730 7324 6736 7336
rect 6691 7296 6736 7324
rect 6730 7284 6736 7296
rect 6788 7284 6794 7336
rect 11330 7324 11336 7336
rect 7760 7296 11336 7324
rect 6472 7256 6500 7284
rect 7760 7256 7788 7296
rect 11330 7284 11336 7296
rect 11388 7324 11394 7336
rect 11532 7324 11560 7355
rect 11606 7352 11612 7404
rect 11664 7392 11670 7404
rect 17037 7395 17095 7401
rect 11664 7364 16160 7392
rect 11664 7352 11670 7364
rect 11388 7296 11560 7324
rect 11388 7284 11394 7296
rect 6472 7228 7788 7256
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 8849 7259 8907 7265
rect 8849 7256 8861 7259
rect 7892 7228 8861 7256
rect 7892 7216 7898 7228
rect 8849 7225 8861 7228
rect 8895 7225 8907 7259
rect 8849 7219 8907 7225
rect 13265 7259 13323 7265
rect 13265 7225 13277 7259
rect 13311 7256 13323 7259
rect 15010 7256 15016 7268
rect 13311 7228 15016 7256
rect 13311 7225 13323 7228
rect 13265 7219 13323 7225
rect 15010 7216 15016 7228
rect 15068 7216 15074 7268
rect 16132 7265 16160 7364
rect 17037 7361 17049 7395
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 18049 7395 18107 7401
rect 18049 7361 18061 7395
rect 18095 7392 18107 7395
rect 18690 7392 18696 7404
rect 18095 7364 18696 7392
rect 18095 7361 18107 7364
rect 18049 7355 18107 7361
rect 16117 7259 16175 7265
rect 16117 7225 16129 7259
rect 16163 7256 16175 7259
rect 16758 7256 16764 7268
rect 16163 7228 16764 7256
rect 16163 7225 16175 7228
rect 16117 7219 16175 7225
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 17052 7256 17080 7355
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 19521 7395 19579 7401
rect 19521 7361 19533 7395
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 18322 7324 18328 7336
rect 18283 7296 18328 7324
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 19536 7256 19564 7355
rect 19628 7324 19656 7432
rect 20916 7401 20944 7500
rect 22925 7497 22937 7531
rect 22971 7528 22983 7531
rect 23290 7528 23296 7540
rect 22971 7500 23296 7528
rect 22971 7497 22983 7500
rect 22925 7491 22983 7497
rect 23290 7488 23296 7500
rect 23348 7488 23354 7540
rect 24210 7488 24216 7540
rect 24268 7528 24274 7540
rect 26050 7528 26056 7540
rect 24268 7500 24532 7528
rect 26011 7500 26056 7528
rect 24268 7488 24274 7500
rect 22649 7463 22707 7469
rect 21008 7432 22416 7460
rect 20901 7395 20959 7401
rect 20901 7361 20913 7395
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 21008 7324 21036 7432
rect 22388 7401 22416 7432
rect 22649 7429 22661 7463
rect 22695 7460 22707 7463
rect 23842 7460 23848 7472
rect 22695 7432 23848 7460
rect 22695 7429 22707 7432
rect 22649 7423 22707 7429
rect 23842 7420 23848 7432
rect 23900 7420 23906 7472
rect 24121 7463 24179 7469
rect 24121 7429 24133 7463
rect 24167 7460 24179 7463
rect 24394 7460 24400 7472
rect 24167 7432 24400 7460
rect 24167 7429 24179 7432
rect 24121 7423 24179 7429
rect 24394 7420 24400 7432
rect 24452 7420 24458 7472
rect 24504 7460 24532 7500
rect 26050 7488 26056 7500
rect 26108 7488 26114 7540
rect 27157 7531 27215 7537
rect 27157 7497 27169 7531
rect 27203 7528 27215 7531
rect 27706 7528 27712 7540
rect 27203 7500 27712 7528
rect 27203 7497 27215 7500
rect 27157 7491 27215 7497
rect 27706 7488 27712 7500
rect 27764 7528 27770 7540
rect 35989 7531 36047 7537
rect 35989 7528 36001 7531
rect 27764 7500 28488 7528
rect 27764 7488 27770 7500
rect 28460 7469 28488 7500
rect 31726 7500 36001 7528
rect 28445 7463 28503 7469
rect 24504 7432 27108 7460
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7392 21143 7395
rect 22373 7395 22431 7401
rect 21131 7364 22094 7392
rect 21131 7361 21143 7364
rect 21085 7355 21143 7361
rect 19628 7296 21036 7324
rect 22066 7324 22094 7364
rect 22373 7361 22385 7395
rect 22419 7361 22431 7395
rect 22554 7392 22560 7404
rect 22515 7364 22560 7392
rect 22373 7355 22431 7361
rect 22554 7352 22560 7364
rect 22612 7352 22618 7404
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7392 22799 7395
rect 23198 7392 23204 7404
rect 22787 7364 23204 7392
rect 22787 7361 22799 7364
rect 22741 7355 22799 7361
rect 23198 7352 23204 7364
rect 23256 7352 23262 7404
rect 24302 7392 24308 7404
rect 24263 7364 24308 7392
rect 24302 7352 24308 7364
rect 24360 7352 24366 7404
rect 25130 7352 25136 7404
rect 25188 7392 25194 7404
rect 25409 7395 25467 7401
rect 25409 7392 25421 7395
rect 25188 7364 25421 7392
rect 25188 7352 25194 7364
rect 25409 7361 25421 7364
rect 25455 7361 25467 7395
rect 25590 7392 25596 7404
rect 25551 7364 25596 7392
rect 25409 7355 25467 7361
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 25685 7395 25743 7401
rect 25685 7361 25697 7395
rect 25731 7361 25743 7395
rect 25685 7355 25743 7361
rect 25777 7395 25835 7401
rect 25777 7361 25789 7395
rect 25823 7392 25835 7395
rect 25958 7392 25964 7404
rect 25823 7364 25964 7392
rect 25823 7361 25835 7364
rect 25777 7355 25835 7361
rect 22572 7324 22600 7352
rect 22066 7296 22600 7324
rect 25498 7284 25504 7336
rect 25556 7324 25562 7336
rect 25700 7324 25728 7355
rect 25958 7352 25964 7364
rect 26016 7352 26022 7404
rect 26973 7395 27031 7401
rect 26973 7361 26985 7395
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 25556 7296 25728 7324
rect 25556 7284 25562 7296
rect 19978 7256 19984 7268
rect 17052 7228 19380 7256
rect 19536 7228 19984 7256
rect 19352 7200 19380 7228
rect 19978 7216 19984 7228
rect 20036 7256 20042 7268
rect 21269 7259 21327 7265
rect 21269 7256 21281 7259
rect 20036 7228 21281 7256
rect 20036 7216 20042 7228
rect 21269 7225 21281 7228
rect 21315 7256 21327 7259
rect 26988 7256 27016 7355
rect 27080 7324 27108 7432
rect 28445 7429 28457 7463
rect 28491 7429 28503 7463
rect 28445 7423 28503 7429
rect 30561 7463 30619 7469
rect 30561 7429 30573 7463
rect 30607 7460 30619 7463
rect 31018 7460 31024 7472
rect 30607 7432 31024 7460
rect 30607 7429 30619 7432
rect 30561 7423 30619 7429
rect 27614 7352 27620 7404
rect 27672 7392 27678 7404
rect 28261 7395 28319 7401
rect 28261 7392 28273 7395
rect 27672 7364 28273 7392
rect 27672 7352 27678 7364
rect 28261 7361 28273 7364
rect 28307 7392 28319 7395
rect 28350 7392 28356 7404
rect 28307 7364 28356 7392
rect 28307 7361 28319 7364
rect 28261 7355 28319 7361
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 28460 7392 28488 7423
rect 31018 7420 31024 7432
rect 31076 7420 31082 7472
rect 30745 7395 30803 7401
rect 30745 7392 30757 7395
rect 28460 7364 30757 7392
rect 30745 7361 30757 7364
rect 30791 7392 30803 7395
rect 31202 7392 31208 7404
rect 30791 7364 31208 7392
rect 30791 7361 30803 7364
rect 30745 7355 30803 7361
rect 31202 7352 31208 7364
rect 31260 7352 31266 7404
rect 31726 7324 31754 7500
rect 35989 7497 36001 7500
rect 36035 7497 36047 7531
rect 35989 7491 36047 7497
rect 33134 7420 33140 7472
rect 33192 7460 33198 7472
rect 33606 7463 33664 7469
rect 33606 7460 33618 7463
rect 33192 7432 33618 7460
rect 33192 7420 33198 7432
rect 33606 7429 33618 7432
rect 33652 7429 33664 7463
rect 33606 7423 33664 7429
rect 35434 7420 35440 7472
rect 35492 7460 35498 7472
rect 36357 7463 36415 7469
rect 36357 7460 36369 7463
rect 35492 7432 36369 7460
rect 35492 7420 35498 7432
rect 36357 7429 36369 7432
rect 36403 7429 36415 7463
rect 38838 7460 38844 7472
rect 38799 7432 38844 7460
rect 36357 7423 36415 7429
rect 38838 7420 38844 7432
rect 38896 7420 38902 7472
rect 33870 7392 33876 7404
rect 33831 7364 33876 7392
rect 33870 7352 33876 7364
rect 33928 7352 33934 7404
rect 35115 7395 35173 7401
rect 35115 7392 35127 7395
rect 34348 7364 35127 7392
rect 27080 7296 31754 7324
rect 21315 7228 27016 7256
rect 21315 7225 21327 7228
rect 21269 7219 21327 7225
rect 31570 7216 31576 7268
rect 31628 7256 31634 7268
rect 32493 7259 32551 7265
rect 32493 7256 32505 7259
rect 31628 7228 32505 7256
rect 31628 7216 31634 7228
rect 32493 7225 32505 7228
rect 32539 7225 32551 7259
rect 32493 7219 32551 7225
rect 1762 7188 1768 7200
rect 1723 7160 1768 7188
rect 1762 7148 1768 7160
rect 1820 7148 1826 7200
rect 2869 7191 2927 7197
rect 2869 7157 2881 7191
rect 2915 7188 2927 7191
rect 3142 7188 3148 7200
rect 2915 7160 3148 7188
rect 2915 7157 2927 7160
rect 2869 7151 2927 7157
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3421 7191 3479 7197
rect 3421 7157 3433 7191
rect 3467 7188 3479 7191
rect 3970 7188 3976 7200
rect 3467 7160 3976 7188
rect 3467 7157 3479 7160
rect 3421 7151 3479 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 7742 7188 7748 7200
rect 4571 7160 7748 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8389 7191 8447 7197
rect 8389 7157 8401 7191
rect 8435 7188 8447 7191
rect 9214 7188 9220 7200
rect 8435 7160 9220 7188
rect 8435 7157 8447 7160
rect 8389 7151 8447 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 10318 7188 10324 7200
rect 10279 7160 10324 7188
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 13817 7191 13875 7197
rect 13817 7157 13829 7191
rect 13863 7188 13875 7191
rect 14274 7188 14280 7200
rect 13863 7160 14280 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 14369 7191 14427 7197
rect 14369 7157 14381 7191
rect 14415 7188 14427 7191
rect 14734 7188 14740 7200
rect 14415 7160 14740 7188
rect 14415 7157 14427 7160
rect 14369 7151 14427 7157
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 16666 7188 16672 7200
rect 16627 7160 16672 7188
rect 16666 7148 16672 7160
rect 16724 7148 16730 7200
rect 17589 7191 17647 7197
rect 17589 7157 17601 7191
rect 17635 7188 17647 7191
rect 17954 7188 17960 7200
rect 17635 7160 17960 7188
rect 17635 7157 17647 7160
rect 17589 7151 17647 7157
rect 17954 7148 17960 7160
rect 18012 7148 18018 7200
rect 19334 7188 19340 7200
rect 19295 7160 19340 7188
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 23474 7188 23480 7200
rect 23435 7160 23480 7188
rect 23474 7148 23480 7160
rect 23532 7148 23538 7200
rect 23937 7191 23995 7197
rect 23937 7157 23949 7191
rect 23983 7188 23995 7191
rect 24578 7188 24584 7200
rect 23983 7160 24584 7188
rect 23983 7157 23995 7160
rect 23937 7151 23995 7157
rect 24578 7148 24584 7160
rect 24636 7148 24642 7200
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25958 7188 25964 7200
rect 24995 7160 25964 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 27982 7148 27988 7200
rect 28040 7188 28046 7200
rect 28077 7191 28135 7197
rect 28077 7188 28089 7191
rect 28040 7160 28089 7188
rect 28040 7148 28046 7160
rect 28077 7157 28089 7160
rect 28123 7157 28135 7191
rect 28077 7151 28135 7157
rect 29822 7148 29828 7200
rect 29880 7188 29886 7200
rect 30377 7191 30435 7197
rect 30377 7188 30389 7191
rect 29880 7160 30389 7188
rect 29880 7148 29886 7160
rect 30377 7157 30389 7160
rect 30423 7157 30435 7191
rect 30377 7151 30435 7157
rect 30926 7148 30932 7200
rect 30984 7188 30990 7200
rect 34348 7197 34376 7364
rect 35115 7361 35127 7364
rect 35161 7361 35173 7395
rect 35250 7392 35256 7404
rect 35211 7364 35256 7392
rect 35115 7355 35173 7361
rect 35130 7256 35158 7355
rect 35250 7352 35256 7364
rect 35308 7352 35314 7404
rect 35345 7395 35403 7401
rect 35345 7361 35357 7395
rect 35391 7361 35403 7395
rect 35526 7392 35532 7404
rect 35487 7364 35532 7392
rect 35345 7355 35403 7361
rect 35360 7324 35388 7355
rect 35526 7352 35532 7364
rect 35584 7352 35590 7404
rect 35710 7352 35716 7404
rect 35768 7392 35774 7404
rect 36173 7395 36231 7401
rect 36173 7392 36185 7395
rect 35768 7364 36185 7392
rect 35768 7352 35774 7364
rect 36173 7361 36185 7364
rect 36219 7361 36231 7395
rect 36173 7355 36231 7361
rect 36262 7352 36268 7404
rect 36320 7392 36326 7404
rect 36541 7395 36599 7401
rect 36320 7364 36365 7392
rect 36320 7352 36326 7364
rect 36541 7361 36553 7395
rect 36587 7392 36599 7395
rect 37090 7392 37096 7404
rect 36587 7364 37096 7392
rect 36587 7361 36599 7364
rect 36541 7355 36599 7361
rect 37090 7352 37096 7364
rect 37148 7352 37154 7404
rect 38286 7352 38292 7404
rect 38344 7392 38350 7404
rect 38657 7395 38715 7401
rect 38657 7392 38669 7395
rect 38344 7364 38669 7392
rect 38344 7352 38350 7364
rect 38657 7361 38669 7364
rect 38703 7361 38715 7395
rect 38657 7355 38715 7361
rect 36906 7324 36912 7336
rect 35360 7296 36912 7324
rect 36906 7284 36912 7296
rect 36964 7284 36970 7336
rect 36170 7256 36176 7268
rect 35130 7228 36176 7256
rect 36170 7216 36176 7228
rect 36228 7216 36234 7268
rect 34333 7191 34391 7197
rect 34333 7188 34345 7191
rect 30984 7160 34345 7188
rect 30984 7148 30990 7160
rect 34333 7157 34345 7160
rect 34379 7157 34391 7191
rect 34333 7151 34391 7157
rect 34790 7148 34796 7200
rect 34848 7188 34854 7200
rect 34885 7191 34943 7197
rect 34885 7188 34897 7191
rect 34848 7160 34897 7188
rect 34848 7148 34854 7160
rect 34885 7157 34897 7160
rect 34931 7157 34943 7191
rect 34885 7151 34943 7157
rect 38930 7148 38936 7200
rect 38988 7188 38994 7200
rect 39025 7191 39083 7197
rect 39025 7188 39037 7191
rect 38988 7160 39037 7188
rect 38988 7148 38994 7160
rect 39025 7157 39037 7160
rect 39071 7157 39083 7191
rect 39025 7151 39083 7157
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 3234 6984 3240 6996
rect 2556 6956 3240 6984
rect 2556 6944 2562 6956
rect 3234 6944 3240 6956
rect 3292 6944 3298 6996
rect 15378 6984 15384 6996
rect 15339 6956 15384 6984
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 27614 6984 27620 6996
rect 27575 6956 27620 6984
rect 27614 6944 27620 6956
rect 27672 6944 27678 6996
rect 30926 6984 30932 6996
rect 28092 6956 30932 6984
rect 3878 6876 3884 6928
rect 3936 6916 3942 6928
rect 9858 6916 9864 6928
rect 3936 6888 4384 6916
rect 3936 6876 3942 6888
rect 2501 6851 2559 6857
rect 2501 6817 2513 6851
rect 2547 6848 2559 6851
rect 2590 6848 2596 6860
rect 2547 6820 2596 6848
rect 2547 6817 2559 6820
rect 2501 6811 2559 6817
rect 2590 6808 2596 6820
rect 2648 6808 2654 6860
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 4120 6820 4292 6848
rect 4120 6808 4126 6820
rect 2314 6780 2320 6792
rect 2275 6752 2320 6780
rect 2314 6740 2320 6752
rect 2372 6740 2378 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4264 6789 4292 6820
rect 4356 6789 4384 6888
rect 9140 6888 9864 6916
rect 5534 6848 5540 6860
rect 4540 6820 5540 6848
rect 4540 6789 4568 6820
rect 5534 6808 5540 6820
rect 5592 6848 5598 6860
rect 6730 6848 6736 6860
rect 5592 6820 6736 6848
rect 5592 6808 5598 6820
rect 6730 6808 6736 6820
rect 6788 6848 6794 6860
rect 6788 6820 8248 6848
rect 6788 6808 6794 6820
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3936 6752 3985 6780
rect 3936 6740 3942 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6749 4215 6783
rect 4157 6743 4215 6749
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 3602 6712 3608 6724
rect 1719 6684 3608 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 3602 6672 3608 6684
rect 3660 6672 3666 6724
rect 2130 6644 2136 6656
rect 2091 6616 2136 6644
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3326 6644 3332 6656
rect 3283 6616 3332 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 3326 6604 3332 6616
rect 3384 6604 3390 6656
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 3476 6616 3801 6644
rect 3476 6604 3482 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 4172 6644 4200 6743
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 6420 6752 6469 6780
rect 6420 6740 6426 6752
rect 6457 6749 6469 6752
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 7190 6740 7196 6792
rect 7248 6780 7254 6792
rect 7285 6783 7343 6789
rect 7285 6780 7297 6783
rect 7248 6752 7297 6780
rect 7248 6740 7254 6752
rect 7285 6749 7297 6752
rect 7331 6749 7343 6783
rect 7285 6743 7343 6749
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 7892 6752 8125 6780
rect 7892 6740 7898 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 8220 6780 8248 6820
rect 9140 6789 9168 6888
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 23474 6916 23480 6928
rect 23387 6888 23480 6916
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 14921 6851 14979 6857
rect 9272 6820 9317 6848
rect 9416 6820 11192 6848
rect 9272 6808 9278 6820
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8220 6752 8953 6780
rect 8113 6743 8171 6749
rect 8941 6749 8953 6752
rect 8987 6780 8999 6783
rect 9125 6783 9183 6789
rect 8987 6752 9076 6780
rect 8987 6749 8999 6752
rect 8941 6743 8999 6749
rect 5074 6672 5080 6724
rect 5132 6712 5138 6724
rect 5445 6715 5503 6721
rect 5445 6712 5457 6715
rect 5132 6684 5457 6712
rect 5132 6672 5138 6684
rect 5445 6681 5457 6684
rect 5491 6712 5503 6715
rect 5810 6712 5816 6724
rect 5491 6684 5816 6712
rect 5491 6681 5503 6684
rect 5445 6675 5503 6681
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 8294 6712 8300 6724
rect 6472 6684 8300 6712
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 4172 6616 5549 6644
rect 3789 6607 3847 6613
rect 5537 6613 5549 6616
rect 5583 6644 5595 6647
rect 6472 6644 6500 6684
rect 8294 6672 8300 6684
rect 8352 6712 8358 6724
rect 9048 6712 9076 6752
rect 9125 6749 9137 6783
rect 9171 6749 9183 6783
rect 9306 6780 9312 6792
rect 9267 6752 9312 6780
rect 9125 6743 9183 6749
rect 9306 6740 9312 6752
rect 9364 6740 9370 6792
rect 9416 6712 9444 6820
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 11054 6780 11060 6792
rect 9539 6752 11060 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11164 6780 11192 6820
rect 14921 6817 14933 6851
rect 14967 6848 14979 6851
rect 15194 6848 15200 6860
rect 14967 6820 15200 6848
rect 14967 6817 14979 6820
rect 14921 6811 14979 6817
rect 15194 6808 15200 6820
rect 15252 6848 15258 6860
rect 16666 6848 16672 6860
rect 15252 6820 15700 6848
rect 15252 6808 15258 6820
rect 11164 6752 12434 6780
rect 8352 6684 8984 6712
rect 9048 6684 9444 6712
rect 10689 6715 10747 6721
rect 8352 6672 8358 6684
rect 8956 6656 8984 6684
rect 10689 6681 10701 6715
rect 10735 6712 10747 6715
rect 12250 6712 12256 6724
rect 10735 6684 12256 6712
rect 10735 6681 10747 6684
rect 10689 6675 10747 6681
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 12406 6712 12434 6752
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 12814 6783 12872 6789
rect 12814 6780 12826 6783
rect 12584 6752 12826 6780
rect 12584 6740 12590 6752
rect 12814 6749 12826 6752
rect 12860 6749 12872 6783
rect 13078 6780 13084 6792
rect 13039 6752 13084 6780
rect 12814 6743 12872 6749
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 15672 6789 15700 6820
rect 15856 6820 16672 6848
rect 15856 6789 15884 6820
rect 16666 6808 16672 6820
rect 16724 6808 16730 6860
rect 16945 6851 17003 6857
rect 16945 6817 16957 6851
rect 16991 6848 17003 6851
rect 17034 6848 17040 6860
rect 16991 6820 17040 6848
rect 16991 6817 17003 6820
rect 16945 6811 17003 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 19426 6808 19432 6860
rect 19484 6808 19490 6860
rect 22186 6848 22192 6860
rect 22147 6820 22192 6848
rect 22186 6808 22192 6820
rect 22244 6808 22250 6860
rect 15657 6783 15715 6789
rect 15657 6749 15669 6783
rect 15703 6749 15715 6783
rect 15657 6743 15715 6749
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 15749 6743 15807 6749
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 16022 6780 16028 6792
rect 15983 6752 16028 6780
rect 15841 6743 15899 6749
rect 12618 6712 12624 6724
rect 12406 6684 12624 6712
rect 12618 6672 12624 6684
rect 12676 6672 12682 6724
rect 15764 6712 15792 6743
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6780 18015 6783
rect 18782 6780 18788 6792
rect 18003 6752 18788 6780
rect 18003 6749 18015 6752
rect 17957 6743 18015 6749
rect 18782 6740 18788 6752
rect 18840 6780 18846 6792
rect 19444 6780 19472 6808
rect 18840 6752 19472 6780
rect 18840 6740 18846 6752
rect 21818 6740 21824 6792
rect 21876 6780 21882 6792
rect 21913 6783 21971 6789
rect 21913 6780 21925 6783
rect 21876 6752 21925 6780
rect 21876 6740 21882 6752
rect 21913 6749 21925 6752
rect 21959 6749 21971 6783
rect 23400 6780 23428 6888
rect 23474 6876 23480 6888
rect 23532 6916 23538 6928
rect 28092 6916 28120 6956
rect 30926 6944 30932 6956
rect 30984 6944 30990 6996
rect 31018 6944 31024 6996
rect 31076 6984 31082 6996
rect 31389 6987 31447 6993
rect 31389 6984 31401 6987
rect 31076 6956 31401 6984
rect 31076 6944 31082 6956
rect 31389 6953 31401 6956
rect 31435 6953 31447 6987
rect 36906 6984 36912 6996
rect 36867 6956 36912 6984
rect 31389 6947 31447 6953
rect 36906 6944 36912 6956
rect 36964 6944 36970 6996
rect 36998 6916 37004 6928
rect 23532 6888 28120 6916
rect 34961 6888 37004 6916
rect 23532 6876 23538 6888
rect 25130 6848 25136 6860
rect 24412 6820 25136 6848
rect 23457 6783 23515 6789
rect 23457 6780 23469 6783
rect 23400 6752 23469 6780
rect 21913 6743 21971 6749
rect 23457 6749 23469 6752
rect 23503 6749 23515 6783
rect 23457 6743 23515 6749
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6749 23627 6783
rect 23569 6743 23627 6749
rect 23661 6783 23719 6789
rect 23661 6749 23673 6783
rect 23707 6780 23719 6783
rect 23750 6780 23756 6792
rect 23707 6752 23756 6780
rect 23707 6749 23719 6752
rect 23661 6743 23719 6749
rect 15930 6712 15936 6724
rect 15764 6684 15936 6712
rect 15930 6672 15936 6684
rect 15988 6712 15994 6724
rect 18322 6712 18328 6724
rect 15988 6684 18328 6712
rect 15988 6672 15994 6684
rect 18322 6672 18328 6684
rect 18380 6672 18386 6724
rect 19429 6715 19487 6721
rect 19429 6681 19441 6715
rect 19475 6712 19487 6715
rect 20162 6712 20168 6724
rect 19475 6684 20168 6712
rect 19475 6681 19487 6684
rect 19429 6675 19487 6681
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 23584 6712 23612 6743
rect 23750 6740 23756 6752
rect 23808 6740 23814 6792
rect 24412 6789 24440 6820
rect 25130 6808 25136 6820
rect 25188 6808 25194 6860
rect 25774 6848 25780 6860
rect 25735 6820 25780 6848
rect 25774 6808 25780 6820
rect 25832 6808 25838 6860
rect 27246 6848 27252 6860
rect 25976 6820 27252 6848
rect 23845 6783 23903 6789
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 23891 6752 24409 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 24578 6780 24584 6792
rect 24539 6752 24584 6780
rect 24397 6743 24455 6749
rect 24578 6740 24584 6752
rect 24636 6740 24642 6792
rect 24673 6783 24731 6789
rect 24673 6749 24685 6783
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 24688 6712 24716 6743
rect 24762 6740 24768 6792
rect 24820 6780 24826 6792
rect 25976 6780 26004 6820
rect 27246 6808 27252 6820
rect 27304 6848 27310 6860
rect 28997 6851 29055 6857
rect 27304 6820 27614 6848
rect 27304 6808 27310 6820
rect 24820 6752 26004 6780
rect 26053 6783 26111 6789
rect 24820 6740 24826 6752
rect 26053 6749 26065 6783
rect 26099 6780 26111 6783
rect 27430 6780 27436 6792
rect 26099 6752 27436 6780
rect 26099 6749 26111 6752
rect 26053 6743 26111 6749
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 27586 6780 27614 6820
rect 28997 6817 29009 6851
rect 29043 6848 29055 6851
rect 30006 6848 30012 6860
rect 29043 6820 30012 6848
rect 29043 6817 29055 6820
rect 28997 6811 29055 6817
rect 30006 6808 30012 6820
rect 30064 6808 30070 6860
rect 34961 6789 34989 6888
rect 36998 6876 37004 6888
rect 37056 6876 37062 6928
rect 35434 6848 35440 6860
rect 35084 6820 35440 6848
rect 35084 6789 35112 6820
rect 35434 6808 35440 6820
rect 35492 6808 35498 6860
rect 36449 6851 36507 6857
rect 36449 6817 36461 6851
rect 36495 6848 36507 6851
rect 38378 6848 38384 6860
rect 36495 6820 38384 6848
rect 36495 6817 36507 6820
rect 36449 6811 36507 6817
rect 38378 6808 38384 6820
rect 38436 6808 38442 6860
rect 38654 6808 38660 6860
rect 38712 6848 38718 6860
rect 38712 6820 38884 6848
rect 38712 6808 38718 6820
rect 34057 6783 34115 6789
rect 34057 6780 34069 6783
rect 27586 6752 34069 6780
rect 34057 6749 34069 6752
rect 34103 6780 34115 6783
rect 34931 6783 34989 6789
rect 34931 6780 34943 6783
rect 34103 6752 34943 6780
rect 34103 6749 34115 6752
rect 34057 6743 34115 6749
rect 34931 6749 34943 6752
rect 34977 6749 34989 6783
rect 34931 6743 34989 6749
rect 35069 6783 35127 6789
rect 35069 6749 35081 6783
rect 35115 6749 35127 6783
rect 35069 6743 35127 6749
rect 35182 6783 35240 6789
rect 35182 6749 35194 6783
rect 35228 6780 35240 6783
rect 35345 6783 35403 6789
rect 35228 6752 35296 6780
rect 35228 6749 35240 6752
rect 35182 6743 35240 6749
rect 25498 6712 25504 6724
rect 23584 6684 25504 6712
rect 25498 6672 25504 6684
rect 25556 6672 25562 6724
rect 27522 6672 27528 6724
rect 27580 6712 27586 6724
rect 28730 6715 28788 6721
rect 28730 6712 28742 6715
rect 27580 6684 28742 6712
rect 27580 6672 27586 6684
rect 28730 6681 28742 6684
rect 28776 6681 28788 6715
rect 28730 6675 28788 6681
rect 30276 6715 30334 6721
rect 30276 6681 30288 6715
rect 30322 6712 30334 6715
rect 30374 6712 30380 6724
rect 30322 6684 30380 6712
rect 30322 6681 30334 6684
rect 30276 6675 30334 6681
rect 30374 6672 30380 6684
rect 30432 6672 30438 6724
rect 6638 6644 6644 6656
rect 5583 6616 6500 6644
rect 6599 6616 6644 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 7469 6647 7527 6653
rect 7469 6644 7481 6647
rect 6880 6616 7481 6644
rect 6880 6604 6886 6616
rect 7469 6613 7481 6616
rect 7515 6613 7527 6647
rect 7469 6607 7527 6613
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6644 7987 6647
rect 8018 6644 8024 6656
rect 7975 6616 8024 6644
rect 7975 6613 7987 6616
rect 7929 6607 7987 6613
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 8938 6604 8944 6656
rect 8996 6604 9002 6656
rect 9674 6644 9680 6656
rect 9635 6616 9680 6644
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 11238 6644 11244 6656
rect 11199 6616 11244 6644
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11698 6644 11704 6656
rect 11572 6616 11704 6644
rect 11572 6604 11578 6616
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 16850 6644 16856 6656
rect 14415 6616 16856 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 18414 6644 18420 6656
rect 18375 6616 18420 6644
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 20714 6644 20720 6656
rect 20675 6616 20720 6644
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 20990 6604 20996 6656
rect 21048 6644 21054 6656
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 21048 6616 21189 6644
rect 21048 6604 21054 6616
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 23201 6647 23259 6653
rect 23201 6613 23213 6647
rect 23247 6644 23259 6647
rect 23566 6644 23572 6656
rect 23247 6616 23572 6644
rect 23247 6613 23259 6616
rect 23201 6607 23259 6613
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 25038 6644 25044 6656
rect 24999 6616 25044 6644
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 27062 6644 27068 6656
rect 27023 6616 27068 6644
rect 27062 6604 27068 6616
rect 27120 6644 27126 6656
rect 30650 6644 30656 6656
rect 27120 6616 30656 6644
rect 27120 6604 27126 6616
rect 30650 6604 30656 6616
rect 30708 6644 30714 6656
rect 31110 6644 31116 6656
rect 30708 6616 31116 6644
rect 30708 6604 30714 6616
rect 31110 6604 31116 6616
rect 31168 6604 31174 6656
rect 34606 6604 34612 6656
rect 34664 6644 34670 6656
rect 34701 6647 34759 6653
rect 34701 6644 34713 6647
rect 34664 6616 34713 6644
rect 34664 6604 34670 6616
rect 34701 6613 34713 6616
rect 34747 6613 34759 6647
rect 35268 6644 35296 6752
rect 35345 6749 35357 6783
rect 35391 6780 35403 6783
rect 35526 6780 35532 6792
rect 35391 6752 35532 6780
rect 35391 6749 35403 6752
rect 35345 6743 35403 6749
rect 35526 6740 35532 6752
rect 35584 6740 35590 6792
rect 35805 6783 35863 6789
rect 35805 6749 35817 6783
rect 35851 6749 35863 6783
rect 35986 6780 35992 6792
rect 35947 6752 35992 6780
rect 35805 6743 35863 6749
rect 35820 6712 35848 6743
rect 35986 6740 35992 6752
rect 36044 6740 36050 6792
rect 36081 6783 36139 6789
rect 36081 6749 36093 6783
rect 36127 6749 36139 6783
rect 36081 6743 36139 6749
rect 35894 6712 35900 6724
rect 35820 6684 35900 6712
rect 35894 6672 35900 6684
rect 35952 6672 35958 6724
rect 36096 6656 36124 6743
rect 36170 6740 36176 6792
rect 36228 6780 36234 6792
rect 36228 6752 36273 6780
rect 36228 6740 36234 6752
rect 36998 6740 37004 6792
rect 37056 6780 37062 6792
rect 38856 6789 38884 6820
rect 38749 6783 38807 6789
rect 38749 6780 38761 6783
rect 37056 6752 38761 6780
rect 37056 6740 37062 6752
rect 38749 6749 38761 6752
rect 38795 6749 38807 6783
rect 38749 6743 38807 6749
rect 38841 6783 38899 6789
rect 38841 6749 38853 6783
rect 38887 6749 38899 6783
rect 38841 6743 38899 6749
rect 37090 6712 37096 6724
rect 37051 6684 37096 6712
rect 37090 6672 37096 6684
rect 37148 6672 37154 6724
rect 37277 6715 37335 6721
rect 37277 6681 37289 6715
rect 37323 6712 37335 6715
rect 37366 6712 37372 6724
rect 37323 6684 37372 6712
rect 37323 6681 37335 6684
rect 37277 6675 37335 6681
rect 37366 6672 37372 6684
rect 37424 6672 37430 6724
rect 38013 6715 38071 6721
rect 38013 6681 38025 6715
rect 38059 6712 38071 6715
rect 38764 6712 38792 6743
rect 38930 6740 38936 6792
rect 38988 6780 38994 6792
rect 39117 6783 39175 6789
rect 38988 6752 39033 6780
rect 38988 6740 38994 6752
rect 39117 6749 39129 6783
rect 39163 6780 39175 6783
rect 39298 6780 39304 6792
rect 39163 6752 39304 6780
rect 39163 6749 39175 6752
rect 39117 6743 39175 6749
rect 39298 6740 39304 6752
rect 39356 6740 39362 6792
rect 39853 6715 39911 6721
rect 39853 6712 39865 6715
rect 38059 6684 38700 6712
rect 38764 6684 39865 6712
rect 38059 6681 38071 6684
rect 38013 6675 38071 6681
rect 35342 6644 35348 6656
rect 35268 6616 35348 6644
rect 34701 6607 34759 6613
rect 35342 6604 35348 6616
rect 35400 6604 35406 6656
rect 36078 6604 36084 6656
rect 36136 6604 36142 6656
rect 38473 6647 38531 6653
rect 38473 6613 38485 6647
rect 38519 6644 38531 6647
rect 38562 6644 38568 6656
rect 38519 6616 38568 6644
rect 38519 6613 38531 6616
rect 38473 6607 38531 6613
rect 38562 6604 38568 6616
rect 38620 6604 38626 6656
rect 38672 6644 38700 6684
rect 39853 6681 39865 6684
rect 39899 6681 39911 6715
rect 39853 6675 39911 6681
rect 39298 6644 39304 6656
rect 38672 6616 39304 6644
rect 39298 6604 39304 6616
rect 39356 6604 39362 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 6454 6440 6460 6452
rect 6415 6412 6460 6440
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 11238 6400 11244 6452
rect 11296 6440 11302 6452
rect 14826 6440 14832 6452
rect 11296 6412 14832 6440
rect 11296 6400 11302 6412
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 15289 6443 15347 6449
rect 15289 6409 15301 6443
rect 15335 6440 15347 6443
rect 17310 6440 17316 6452
rect 15335 6412 17316 6440
rect 15335 6409 15347 6412
rect 15289 6403 15347 6409
rect 3234 6372 3240 6384
rect 3195 6344 3240 6372
rect 3234 6332 3240 6344
rect 3292 6332 3298 6384
rect 3326 6332 3332 6384
rect 3384 6372 3390 6384
rect 4985 6375 5043 6381
rect 4985 6372 4997 6375
rect 3384 6344 4997 6372
rect 3384 6332 3390 6344
rect 4985 6341 4997 6344
rect 5031 6372 5043 6375
rect 6546 6372 6552 6384
rect 5031 6344 6552 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 6546 6332 6552 6344
rect 6604 6332 6610 6384
rect 11422 6372 11428 6384
rect 9140 6344 11428 6372
rect 1489 6307 1547 6313
rect 1489 6273 1501 6307
rect 1535 6304 1547 6307
rect 2130 6304 2136 6316
rect 1535 6276 2136 6304
rect 1535 6273 1547 6276
rect 1489 6267 1547 6273
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6304 2835 6307
rect 5813 6307 5871 6313
rect 5813 6304 5825 6307
rect 2823 6276 5825 6304
rect 2823 6273 2835 6276
rect 2777 6267 2835 6273
rect 5813 6273 5825 6276
rect 5859 6304 5871 6307
rect 6270 6304 6276 6316
rect 5859 6276 6276 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6270 6264 6276 6276
rect 6328 6264 6334 6316
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6304 7159 6307
rect 7282 6304 7288 6316
rect 7147 6276 7288 6304
rect 7147 6273 7159 6276
rect 7101 6267 7159 6273
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 6380 6236 6408 6267
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8018 6304 8024 6316
rect 7975 6276 8024 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8386 6304 8392 6316
rect 8347 6276 8392 6304
rect 8386 6264 8392 6276
rect 8444 6264 8450 6316
rect 9140 6313 9168 6344
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 12345 6375 12403 6381
rect 12345 6341 12357 6375
rect 12391 6372 12403 6375
rect 12391 6344 13032 6372
rect 12391 6341 12403 6344
rect 12345 6335 12403 6341
rect 9125 6307 9183 6313
rect 9125 6273 9137 6307
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9392 6307 9450 6313
rect 9392 6273 9404 6307
rect 9438 6304 9450 6307
rect 9674 6304 9680 6316
rect 9438 6276 9680 6304
rect 9438 6273 9450 6276
rect 9392 6267 9450 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 12894 6236 12900 6248
rect 5408 6208 6408 6236
rect 7116 6208 9168 6236
rect 5408 6196 5414 6208
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 7116 6168 7144 6208
rect 4764 6140 7144 6168
rect 7285 6171 7343 6177
rect 4764 6128 4770 6140
rect 7285 6137 7297 6171
rect 7331 6168 7343 6171
rect 8386 6168 8392 6180
rect 7331 6140 8392 6168
rect 7331 6137 7343 6140
rect 7285 6131 7343 6137
rect 8386 6128 8392 6140
rect 8444 6128 8450 6180
rect 1670 6100 1676 6112
rect 1631 6072 1676 6100
rect 1670 6060 1676 6072
rect 1728 6060 1734 6112
rect 2222 6100 2228 6112
rect 2183 6072 2228 6100
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 4614 6100 4620 6112
rect 2740 6072 4620 6100
rect 2740 6060 2746 6072
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 5626 6100 5632 6112
rect 5587 6072 5632 6100
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 7616 6072 7757 6100
rect 7616 6060 7622 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 8573 6103 8631 6109
rect 8573 6069 8585 6103
rect 8619 6100 8631 6103
rect 9030 6100 9036 6112
rect 8619 6072 9036 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 9140 6100 9168 6208
rect 10152 6208 12900 6236
rect 10152 6100 10180 6208
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 13004 6236 13032 6344
rect 13078 6332 13084 6384
rect 13136 6372 13142 6384
rect 15562 6372 15568 6384
rect 13136 6344 15568 6372
rect 13136 6332 13142 6344
rect 13924 6313 13952 6344
rect 15562 6332 15568 6344
rect 15620 6332 15626 6384
rect 15948 6381 15976 6412
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 20530 6400 20536 6452
rect 20588 6440 20594 6452
rect 21910 6440 21916 6452
rect 20588 6412 21916 6440
rect 20588 6400 20594 6412
rect 21910 6400 21916 6412
rect 21968 6400 21974 6452
rect 23658 6440 23664 6452
rect 23619 6412 23664 6440
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 24026 6400 24032 6452
rect 24084 6440 24090 6452
rect 24213 6443 24271 6449
rect 24213 6440 24225 6443
rect 24084 6412 24225 6440
rect 24084 6400 24090 6412
rect 24213 6409 24225 6412
rect 24259 6440 24271 6443
rect 24762 6440 24768 6452
rect 24259 6412 24768 6440
rect 24259 6409 24271 6412
rect 24213 6403 24271 6409
rect 24762 6400 24768 6412
rect 24820 6400 24826 6452
rect 25130 6440 25136 6452
rect 25043 6412 25136 6440
rect 25130 6400 25136 6412
rect 25188 6440 25194 6452
rect 25682 6440 25688 6452
rect 25188 6412 25688 6440
rect 25188 6400 25194 6412
rect 25682 6400 25688 6412
rect 25740 6400 25746 6452
rect 27522 6440 27528 6452
rect 27483 6412 27528 6440
rect 27522 6400 27528 6412
rect 27580 6400 27586 6452
rect 29178 6440 29184 6452
rect 29139 6412 29184 6440
rect 29178 6400 29184 6412
rect 29236 6440 29242 6452
rect 30098 6440 30104 6452
rect 29236 6412 30104 6440
rect 29236 6400 29242 6412
rect 30098 6400 30104 6412
rect 30156 6400 30162 6452
rect 30374 6440 30380 6452
rect 30335 6412 30380 6440
rect 30374 6400 30380 6412
rect 30432 6400 30438 6452
rect 36081 6443 36139 6449
rect 36081 6409 36093 6443
rect 36127 6440 36139 6443
rect 37090 6440 37096 6452
rect 36127 6412 37096 6440
rect 36127 6409 36139 6412
rect 36081 6403 36139 6409
rect 37090 6400 37096 6412
rect 37148 6400 37154 6452
rect 38838 6400 38844 6452
rect 38896 6440 38902 6452
rect 39669 6443 39727 6449
rect 39669 6440 39681 6443
rect 38896 6412 39681 6440
rect 38896 6400 38902 6412
rect 39669 6409 39681 6412
rect 39715 6409 39727 6443
rect 39669 6403 39727 6409
rect 15933 6375 15991 6381
rect 15933 6341 15945 6375
rect 15979 6341 15991 6375
rect 17034 6372 17040 6384
rect 16995 6344 17040 6372
rect 15933 6335 15991 6341
rect 17034 6332 17040 6344
rect 17092 6332 17098 6384
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 22554 6372 22560 6384
rect 19392 6344 19564 6372
rect 19392 6332 19398 6344
rect 19536 6316 19564 6344
rect 22112 6344 22560 6372
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6273 13967 6307
rect 13909 6267 13967 6273
rect 14176 6307 14234 6313
rect 14176 6273 14188 6307
rect 14222 6304 14234 6307
rect 14458 6304 14464 6316
rect 14222 6276 14464 6304
rect 14222 6273 14234 6276
rect 14176 6267 14234 6273
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 16114 6304 16120 6316
rect 14700 6276 15976 6304
rect 16075 6276 16120 6304
rect 14700 6264 14706 6276
rect 15948 6236 15976 6276
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 19426 6304 19432 6316
rect 19387 6276 19432 6304
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19518 6264 19524 6316
rect 19576 6304 19582 6316
rect 22112 6313 22140 6344
rect 22554 6332 22560 6344
rect 22612 6372 22618 6384
rect 23293 6375 23351 6381
rect 23293 6372 23305 6375
rect 22612 6344 23305 6372
rect 22612 6332 22618 6344
rect 23293 6341 23305 6344
rect 23339 6341 23351 6375
rect 23293 6335 23351 6341
rect 23385 6375 23443 6381
rect 23385 6341 23397 6375
rect 23431 6372 23443 6375
rect 24394 6372 24400 6384
rect 23431 6344 24400 6372
rect 23431 6341 23443 6344
rect 23385 6335 23443 6341
rect 24394 6332 24400 6344
rect 24452 6332 24458 6384
rect 26421 6375 26479 6381
rect 26421 6341 26433 6375
rect 26467 6372 26479 6375
rect 27062 6372 27068 6384
rect 26467 6344 27068 6372
rect 26467 6341 26479 6344
rect 26421 6335 26479 6341
rect 27062 6332 27068 6344
rect 27120 6332 27126 6384
rect 27430 6332 27436 6384
rect 27488 6372 27494 6384
rect 31021 6375 31079 6381
rect 27488 6344 27936 6372
rect 27488 6332 27494 6344
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 19576 6276 19625 6304
rect 19576 6264 19582 6276
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 22097 6307 22155 6313
rect 22097 6273 22109 6307
rect 22143 6273 22155 6307
rect 22097 6267 22155 6273
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6273 23167 6307
rect 23109 6267 23167 6273
rect 18414 6236 18420 6248
rect 13004 6208 13952 6236
rect 15948 6208 18420 6236
rect 11793 6171 11851 6177
rect 11793 6137 11805 6171
rect 11839 6168 11851 6171
rect 13722 6168 13728 6180
rect 11839 6140 13728 6168
rect 11839 6137 11851 6140
rect 11793 6131 11851 6137
rect 13722 6128 13728 6140
rect 13780 6128 13786 6180
rect 9140 6072 10180 6100
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6100 10563 6103
rect 11054 6100 11060 6112
rect 10551 6072 11060 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 11054 6060 11060 6072
rect 11112 6100 11118 6112
rect 11422 6100 11428 6112
rect 11112 6072 11428 6100
rect 11112 6060 11118 6072
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 12894 6100 12900 6112
rect 12855 6072 12900 6100
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13446 6100 13452 6112
rect 13044 6072 13452 6100
rect 13044 6060 13050 6072
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13924 6100 13952 6208
rect 18414 6196 18420 6208
rect 18472 6236 18478 6248
rect 18598 6236 18604 6248
rect 18472 6208 18604 6236
rect 18472 6196 18478 6208
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 18785 6239 18843 6245
rect 18785 6205 18797 6239
rect 18831 6236 18843 6239
rect 19242 6236 19248 6248
rect 18831 6208 19248 6236
rect 18831 6205 18843 6208
rect 18785 6199 18843 6205
rect 19242 6196 19248 6208
rect 19300 6196 19306 6248
rect 21818 6236 21824 6248
rect 21779 6208 21824 6236
rect 21818 6196 21824 6208
rect 21876 6196 21882 6248
rect 18506 6128 18512 6180
rect 18564 6168 18570 6180
rect 23124 6168 23152 6267
rect 23198 6264 23204 6316
rect 23256 6304 23262 6316
rect 23477 6307 23535 6313
rect 23477 6304 23489 6307
rect 23256 6276 23489 6304
rect 23256 6264 23262 6276
rect 23477 6273 23489 6276
rect 23523 6273 23535 6307
rect 26970 6304 26976 6316
rect 26931 6276 26976 6304
rect 23477 6267 23535 6273
rect 26970 6264 26976 6276
rect 27028 6304 27034 6316
rect 27908 6313 27936 6344
rect 31021 6341 31033 6375
rect 31067 6372 31079 6375
rect 31067 6344 31754 6372
rect 31067 6341 31079 6344
rect 31021 6335 31079 6341
rect 27801 6307 27859 6313
rect 27801 6304 27813 6307
rect 27028 6276 27813 6304
rect 27028 6264 27034 6276
rect 27801 6273 27813 6276
rect 27847 6273 27859 6307
rect 27801 6267 27859 6273
rect 27893 6307 27951 6313
rect 27893 6273 27905 6307
rect 27939 6273 27951 6307
rect 27893 6267 27951 6273
rect 27982 6264 27988 6316
rect 28040 6304 28046 6316
rect 28040 6276 28085 6304
rect 28040 6264 28046 6276
rect 28166 6264 28172 6316
rect 28224 6304 28230 6316
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 28224 6276 29745 6304
rect 28224 6264 28230 6276
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 29748 6236 29776 6267
rect 29822 6264 29828 6316
rect 29880 6304 29886 6316
rect 29917 6310 29975 6316
rect 29917 6304 29929 6310
rect 29880 6276 29929 6304
rect 29963 6276 29975 6310
rect 30012 6310 30070 6316
rect 30012 6307 30024 6310
rect 29880 6264 29886 6276
rect 29917 6270 29975 6276
rect 30011 6276 30024 6307
rect 30058 6276 30070 6310
rect 30011 6270 30070 6276
rect 30011 6236 30039 6270
rect 30098 6264 30104 6316
rect 30156 6313 30162 6316
rect 30156 6307 30179 6313
rect 30167 6273 30179 6307
rect 31202 6304 31208 6316
rect 31163 6276 31208 6304
rect 30156 6267 30179 6273
rect 30156 6264 30162 6267
rect 31202 6264 31208 6276
rect 31260 6264 31266 6316
rect 31726 6304 31754 6344
rect 34790 6332 34796 6384
rect 34848 6372 34854 6384
rect 34946 6375 35004 6381
rect 34946 6372 34958 6375
rect 34848 6344 34958 6372
rect 34848 6332 34854 6344
rect 34946 6341 34958 6344
rect 34992 6341 35004 6375
rect 34946 6335 35004 6341
rect 36170 6332 36176 6384
rect 36228 6372 36234 6384
rect 36541 6375 36599 6381
rect 36541 6372 36553 6375
rect 36228 6344 36553 6372
rect 36228 6332 36234 6344
rect 36541 6341 36553 6344
rect 36587 6341 36599 6375
rect 38654 6372 38660 6384
rect 36541 6335 36599 6341
rect 37844 6344 38660 6372
rect 32030 6304 32036 6316
rect 31726 6276 32036 6304
rect 32030 6264 32036 6276
rect 32088 6264 32094 6316
rect 34698 6304 34704 6316
rect 34659 6276 34704 6304
rect 34698 6264 34704 6276
rect 34756 6264 34762 6316
rect 36078 6264 36084 6316
rect 36136 6304 36142 6316
rect 37844 6304 37872 6344
rect 38654 6332 38660 6344
rect 38712 6332 38718 6384
rect 36136 6276 37872 6304
rect 36136 6264 36142 6276
rect 37918 6264 37924 6316
rect 37976 6304 37982 6316
rect 38562 6313 38568 6316
rect 38289 6307 38347 6313
rect 38289 6304 38301 6307
rect 37976 6276 38301 6304
rect 37976 6264 37982 6276
rect 38289 6273 38301 6276
rect 38335 6273 38347 6307
rect 38556 6304 38568 6313
rect 38523 6276 38568 6304
rect 38289 6267 38347 6273
rect 38556 6267 38568 6276
rect 38562 6264 38568 6267
rect 38620 6264 38626 6316
rect 29748 6208 29868 6236
rect 30011 6208 30236 6236
rect 18564 6140 23152 6168
rect 29840 6168 29868 6208
rect 30098 6168 30104 6180
rect 29840 6140 30104 6168
rect 18564 6128 18570 6140
rect 30098 6128 30104 6140
rect 30156 6128 30162 6180
rect 14918 6100 14924 6112
rect 13924 6072 14924 6100
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15746 6100 15752 6112
rect 15707 6072 15752 6100
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 18230 6060 18236 6112
rect 18288 6100 18294 6112
rect 19245 6103 19303 6109
rect 19245 6100 19257 6103
rect 18288 6072 19257 6100
rect 18288 6060 18294 6072
rect 19245 6069 19257 6072
rect 19291 6069 19303 6103
rect 20254 6100 20260 6112
rect 20215 6072 20260 6100
rect 19245 6063 19303 6069
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 20806 6100 20812 6112
rect 20767 6072 20812 6100
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 30006 6060 30012 6112
rect 30064 6100 30070 6112
rect 30208 6100 30236 6208
rect 58158 6168 58164 6180
rect 58119 6140 58164 6168
rect 58158 6128 58164 6140
rect 58216 6128 58222 6180
rect 30064 6072 30236 6100
rect 30064 6060 30070 6072
rect 30374 6060 30380 6112
rect 30432 6100 30438 6112
rect 30837 6103 30895 6109
rect 30837 6100 30849 6103
rect 30432 6072 30849 6100
rect 30432 6060 30438 6072
rect 30837 6069 30849 6072
rect 30883 6069 30895 6103
rect 30837 6063 30895 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4062 5896 4068 5908
rect 4019 5868 4068 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 7650 5896 7656 5908
rect 4540 5868 7656 5896
rect 3237 5831 3295 5837
rect 3237 5797 3249 5831
rect 3283 5797 3295 5831
rect 3237 5791 3295 5797
rect 2866 5720 2872 5772
rect 2924 5760 2930 5772
rect 3252 5760 3280 5791
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 2924 5732 4261 5760
rect 2924 5720 2930 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 1854 5692 1860 5704
rect 1815 5664 1860 5692
rect 1854 5652 1860 5664
rect 1912 5692 1918 5704
rect 2498 5692 2504 5704
rect 1912 5664 2504 5692
rect 1912 5652 1918 5664
rect 2498 5652 2504 5664
rect 2556 5652 2562 5704
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 3878 5692 3884 5704
rect 3384 5664 3884 5692
rect 3384 5652 3390 5664
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5692 4215 5695
rect 4540 5692 4568 5868
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 14458 5896 14464 5908
rect 8168 5868 12434 5896
rect 14419 5868 14464 5896
rect 8168 5856 8174 5868
rect 6178 5788 6184 5840
rect 6236 5828 6242 5840
rect 6546 5828 6552 5840
rect 6236 5800 6552 5828
rect 6236 5788 6242 5800
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 6917 5831 6975 5837
rect 6917 5797 6929 5831
rect 6963 5828 6975 5831
rect 8202 5828 8208 5840
rect 6963 5800 8208 5828
rect 6963 5797 6975 5800
rect 6917 5791 6975 5797
rect 8202 5788 8208 5800
rect 8260 5828 8266 5840
rect 8260 5800 9812 5828
rect 8260 5788 8266 5800
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5760 4675 5763
rect 5718 5760 5724 5772
rect 4663 5732 5724 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 8662 5720 8668 5772
rect 8720 5760 8726 5772
rect 8720 5732 9168 5760
rect 8720 5720 8726 5732
rect 4203 5664 4568 5692
rect 4203 5661 4215 5664
rect 4157 5655 4215 5661
rect 4706 5652 4712 5704
rect 4764 5692 4770 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4764 5664 5457 5692
rect 4764 5652 4770 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5692 5687 5695
rect 5810 5692 5816 5704
rect 5675 5664 5816 5692
rect 5675 5661 5687 5664
rect 5629 5655 5687 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 6086 5692 6092 5704
rect 6047 5664 6092 5692
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6730 5692 6736 5704
rect 6227 5664 6736 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 7742 5692 7748 5704
rect 7423 5664 7748 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5692 8171 5695
rect 8294 5692 8300 5704
rect 8159 5664 8300 5692
rect 8159 5661 8171 5664
rect 8113 5655 8171 5661
rect 8294 5652 8300 5664
rect 8352 5692 8358 5704
rect 8938 5692 8944 5704
rect 8352 5664 8944 5692
rect 8352 5652 8358 5664
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9140 5701 9168 5732
rect 9784 5701 9812 5800
rect 12406 5760 12434 5868
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 18138 5896 18144 5908
rect 16592 5868 18144 5896
rect 12894 5788 12900 5840
rect 12952 5828 12958 5840
rect 16592 5828 16620 5868
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 18248 5868 18460 5896
rect 12952 5800 16620 5828
rect 12952 5788 12958 5800
rect 16666 5788 16672 5840
rect 16724 5828 16730 5840
rect 18248 5828 18276 5868
rect 16724 5800 18276 5828
rect 16724 5788 16730 5800
rect 18322 5788 18328 5840
rect 18380 5788 18386 5840
rect 14642 5760 14648 5772
rect 12406 5732 14648 5760
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 15746 5760 15752 5772
rect 14936 5732 15752 5760
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9769 5695 9827 5701
rect 9769 5661 9781 5695
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10502 5692 10508 5704
rect 10459 5664 10508 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 11054 5692 11060 5704
rect 11015 5664 11060 5692
rect 11054 5652 11060 5664
rect 11112 5652 11118 5704
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 11701 5695 11759 5701
rect 11701 5692 11713 5695
rect 11664 5664 11713 5692
rect 11664 5652 11670 5664
rect 11701 5661 11713 5664
rect 11747 5661 11759 5695
rect 11701 5655 11759 5661
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 12492 5664 12541 5692
rect 12492 5652 12498 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 13320 5664 13369 5692
rect 13320 5652 13326 5664
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 14734 5692 14740 5704
rect 14695 5664 14740 5692
rect 13357 5655 13415 5661
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 14936 5701 14964 5732
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 16022 5760 16028 5772
rect 15856 5732 16028 5760
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 14921 5695 14979 5701
rect 14921 5661 14933 5695
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15105 5695 15163 5701
rect 15105 5661 15117 5695
rect 15151 5692 15163 5695
rect 15286 5692 15292 5704
rect 15151 5664 15292 5692
rect 15151 5661 15163 5664
rect 15105 5655 15163 5661
rect 1670 5584 1676 5636
rect 1728 5624 1734 5636
rect 2102 5627 2160 5633
rect 2102 5624 2114 5627
rect 1728 5596 2114 5624
rect 1728 5584 1734 5596
rect 2102 5593 2114 5596
rect 2148 5593 2160 5627
rect 2102 5587 2160 5593
rect 6365 5627 6423 5633
rect 6365 5593 6377 5627
rect 6411 5624 6423 5627
rect 7926 5624 7932 5636
rect 6411 5596 7932 5624
rect 6411 5593 6423 5596
rect 6365 5587 6423 5593
rect 7926 5584 7932 5596
rect 7984 5624 7990 5636
rect 10870 5624 10876 5636
rect 7984 5596 10876 5624
rect 7984 5584 7990 5596
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 14844 5624 14872 5655
rect 15286 5652 15292 5664
rect 15344 5692 15350 5704
rect 15856 5692 15884 5732
rect 16022 5720 16028 5732
rect 16080 5760 16086 5772
rect 16080 5732 16988 5760
rect 16080 5720 16086 5732
rect 15344 5664 15884 5692
rect 16040 5664 16620 5692
rect 15344 5652 15350 5664
rect 15930 5624 15936 5636
rect 14844 5596 15936 5624
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 16040 5633 16068 5664
rect 16025 5627 16083 5633
rect 16025 5593 16037 5627
rect 16071 5593 16083 5627
rect 16025 5587 16083 5593
rect 16114 5584 16120 5636
rect 16172 5624 16178 5636
rect 16209 5627 16267 5633
rect 16209 5624 16221 5627
rect 16172 5596 16221 5624
rect 16172 5584 16178 5596
rect 16209 5593 16221 5596
rect 16255 5593 16267 5627
rect 16592 5624 16620 5664
rect 16666 5652 16672 5704
rect 16724 5692 16730 5704
rect 16960 5701 16988 5732
rect 16945 5695 17003 5701
rect 16724 5664 16769 5692
rect 16724 5652 16730 5664
rect 16945 5661 16957 5695
rect 16991 5692 17003 5695
rect 18046 5692 18052 5704
rect 16991 5664 18052 5692
rect 16991 5661 17003 5664
rect 16945 5655 17003 5661
rect 18046 5652 18052 5664
rect 18104 5652 18110 5704
rect 18230 5692 18236 5704
rect 18191 5664 18236 5692
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 18340 5701 18368 5788
rect 18432 5760 18460 5868
rect 19426 5856 19432 5908
rect 19484 5896 19490 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 19484 5868 20637 5896
rect 19484 5856 19490 5868
rect 20625 5865 20637 5868
rect 20671 5896 20683 5899
rect 20671 5868 22094 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 22066 5828 22094 5868
rect 23750 5856 23756 5908
rect 23808 5896 23814 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23808 5868 24409 5896
rect 23808 5856 23814 5868
rect 24397 5865 24409 5868
rect 24443 5865 24455 5899
rect 24397 5859 24455 5865
rect 29914 5856 29920 5908
rect 29972 5896 29978 5908
rect 30558 5896 30564 5908
rect 29972 5868 30564 5896
rect 29972 5856 29978 5868
rect 30558 5856 30564 5868
rect 30616 5856 30622 5908
rect 33870 5896 33876 5908
rect 33831 5868 33876 5896
rect 33870 5856 33876 5868
rect 33928 5856 33934 5908
rect 34977 5899 35035 5905
rect 34977 5865 34989 5899
rect 35023 5896 35035 5899
rect 35342 5896 35348 5908
rect 35023 5868 35348 5896
rect 35023 5865 35035 5868
rect 34977 5859 35035 5865
rect 35342 5856 35348 5868
rect 35400 5856 35406 5908
rect 35986 5896 35992 5908
rect 35947 5868 35992 5896
rect 35986 5856 35992 5868
rect 36044 5856 36050 5908
rect 27798 5828 27804 5840
rect 22066 5800 27804 5828
rect 27798 5788 27804 5800
rect 27856 5788 27862 5840
rect 30190 5788 30196 5840
rect 30248 5828 30254 5840
rect 31573 5831 31631 5837
rect 31573 5828 31585 5831
rect 30248 5800 31585 5828
rect 30248 5788 30254 5800
rect 31573 5797 31585 5800
rect 31619 5797 31631 5831
rect 31573 5791 31631 5797
rect 18432 5732 19380 5760
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5692 18475 5695
rect 18782 5692 18788 5704
rect 18463 5664 18788 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 19242 5692 19248 5704
rect 19203 5664 19248 5692
rect 19242 5652 19248 5664
rect 19300 5652 19306 5704
rect 19352 5692 19380 5732
rect 27338 5720 27344 5772
rect 27396 5760 27402 5772
rect 30006 5760 30012 5772
rect 27396 5732 30012 5760
rect 27396 5720 27402 5732
rect 30006 5720 30012 5732
rect 30064 5760 30070 5772
rect 30064 5732 30420 5760
rect 30064 5720 30070 5732
rect 25406 5692 25412 5704
rect 19352 5664 25412 5692
rect 25406 5652 25412 5664
rect 25464 5692 25470 5704
rect 25593 5695 25651 5701
rect 25593 5692 25605 5695
rect 25464 5664 25605 5692
rect 25464 5652 25470 5664
rect 25593 5661 25605 5664
rect 25639 5661 25651 5695
rect 25593 5655 25651 5661
rect 25869 5695 25927 5701
rect 25869 5661 25881 5695
rect 25915 5692 25927 5695
rect 25915 5664 27660 5692
rect 25915 5661 25927 5664
rect 25869 5655 25927 5661
rect 18506 5624 18512 5636
rect 16592 5596 18512 5624
rect 16209 5587 16267 5593
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 5350 5556 5356 5568
rect 4672 5528 5356 5556
rect 4672 5516 4678 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6178 5556 6184 5568
rect 6135 5528 6184 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7561 5559 7619 5565
rect 7561 5556 7573 5559
rect 6604 5528 7573 5556
rect 6604 5516 6610 5528
rect 7561 5525 7573 5528
rect 7607 5556 7619 5559
rect 8110 5556 8116 5568
rect 7607 5528 8116 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8478 5556 8484 5568
rect 8343 5528 8484 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8938 5556 8944 5568
rect 8899 5528 8944 5556
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9585 5559 9643 5565
rect 9585 5556 9597 5559
rect 9088 5528 9597 5556
rect 9088 5516 9094 5528
rect 9585 5525 9597 5528
rect 9631 5525 9643 5559
rect 9585 5519 9643 5525
rect 15470 5516 15476 5568
rect 15528 5556 15534 5568
rect 15841 5559 15899 5565
rect 15841 5556 15853 5559
rect 15528 5528 15853 5556
rect 15528 5516 15534 5528
rect 15841 5525 15853 5528
rect 15887 5525 15899 5559
rect 16224 5556 16252 5587
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 18693 5627 18751 5633
rect 18693 5593 18705 5627
rect 18739 5624 18751 5627
rect 19490 5627 19548 5633
rect 19490 5624 19502 5627
rect 18739 5596 19502 5624
rect 18739 5593 18751 5596
rect 18693 5587 18751 5593
rect 19490 5593 19502 5596
rect 19536 5593 19548 5627
rect 19490 5587 19548 5593
rect 23842 5584 23848 5636
rect 23900 5624 23906 5636
rect 24581 5627 24639 5633
rect 24581 5624 24593 5627
rect 23900 5596 24593 5624
rect 23900 5584 23906 5596
rect 24581 5593 24593 5596
rect 24627 5593 24639 5627
rect 24581 5587 24639 5593
rect 24765 5627 24823 5633
rect 24765 5593 24777 5627
rect 24811 5593 24823 5627
rect 24765 5587 24823 5593
rect 27525 5627 27583 5633
rect 27525 5593 27537 5627
rect 27571 5593 27583 5627
rect 27632 5624 27660 5664
rect 27706 5652 27712 5704
rect 27764 5692 27770 5704
rect 30098 5692 30104 5704
rect 27764 5664 27809 5692
rect 30059 5664 30104 5692
rect 27764 5652 27770 5664
rect 30098 5652 30104 5664
rect 30156 5652 30162 5704
rect 30190 5652 30196 5704
rect 30248 5686 30254 5704
rect 30392 5701 30420 5732
rect 30285 5695 30343 5701
rect 30285 5686 30297 5695
rect 30248 5661 30297 5686
rect 30331 5661 30343 5695
rect 30248 5658 30343 5661
rect 30248 5652 30254 5658
rect 30285 5655 30343 5658
rect 30380 5695 30438 5701
rect 30380 5661 30392 5695
rect 30426 5661 30438 5695
rect 30380 5655 30438 5661
rect 30469 5695 30527 5701
rect 30469 5661 30481 5695
rect 30515 5661 30527 5695
rect 30469 5655 30527 5661
rect 28166 5624 28172 5636
rect 27632 5596 28172 5624
rect 27525 5587 27583 5593
rect 19334 5556 19340 5568
rect 16224 5528 19340 5556
rect 15841 5519 15899 5525
rect 19334 5516 19340 5528
rect 19392 5516 19398 5568
rect 21634 5556 21640 5568
rect 21595 5528 21640 5556
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 22186 5556 22192 5568
rect 22147 5528 22192 5556
rect 22186 5516 22192 5528
rect 22244 5516 22250 5568
rect 22646 5556 22652 5568
rect 22607 5528 22652 5556
rect 22646 5516 22652 5528
rect 22704 5516 22710 5568
rect 23198 5556 23204 5568
rect 23159 5528 23204 5556
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 24302 5516 24308 5568
rect 24360 5556 24366 5568
rect 24780 5556 24808 5587
rect 24360 5528 24808 5556
rect 27341 5559 27399 5565
rect 24360 5516 24366 5528
rect 27341 5525 27353 5559
rect 27387 5556 27399 5559
rect 27430 5556 27436 5568
rect 27387 5528 27436 5556
rect 27387 5525 27399 5528
rect 27341 5519 27399 5525
rect 27430 5516 27436 5528
rect 27488 5516 27494 5568
rect 27540 5556 27568 5587
rect 28166 5584 28172 5596
rect 28224 5584 28230 5636
rect 30484 5624 30512 5655
rect 30650 5652 30656 5704
rect 30708 5692 30714 5704
rect 31662 5692 31668 5704
rect 30708 5664 31668 5692
rect 30708 5652 30714 5664
rect 31662 5652 31668 5664
rect 31720 5692 31726 5704
rect 32401 5695 32459 5701
rect 32401 5692 32413 5695
rect 31720 5664 32413 5692
rect 31720 5652 31726 5664
rect 32401 5661 32413 5664
rect 32447 5661 32459 5695
rect 32401 5655 32459 5661
rect 35161 5695 35219 5701
rect 35161 5661 35173 5695
rect 35207 5692 35219 5695
rect 35618 5692 35624 5704
rect 35207 5664 35624 5692
rect 35207 5661 35219 5664
rect 35161 5655 35219 5661
rect 35618 5652 35624 5664
rect 35676 5652 35682 5704
rect 36173 5695 36231 5701
rect 36173 5661 36185 5695
rect 36219 5692 36231 5695
rect 36262 5692 36268 5704
rect 36219 5664 36268 5692
rect 36219 5661 36231 5664
rect 36173 5655 36231 5661
rect 36262 5652 36268 5664
rect 36320 5652 36326 5704
rect 36357 5695 36415 5701
rect 36357 5661 36369 5695
rect 36403 5692 36415 5695
rect 38286 5692 38292 5704
rect 36403 5664 38292 5692
rect 36403 5661 36415 5664
rect 36357 5655 36415 5661
rect 38286 5652 38292 5664
rect 38344 5652 38350 5704
rect 30558 5624 30564 5636
rect 30484 5596 30564 5624
rect 30558 5584 30564 5596
rect 30616 5584 30622 5636
rect 31202 5624 31208 5636
rect 31163 5596 31208 5624
rect 31202 5584 31208 5596
rect 31260 5584 31266 5636
rect 31389 5627 31447 5633
rect 31389 5593 31401 5627
rect 31435 5624 31447 5627
rect 32122 5624 32128 5636
rect 31435 5596 32128 5624
rect 31435 5593 31447 5596
rect 31389 5587 31447 5593
rect 32122 5584 32128 5596
rect 32180 5584 32186 5636
rect 35345 5627 35403 5633
rect 35345 5593 35357 5627
rect 35391 5593 35403 5627
rect 35345 5587 35403 5593
rect 28534 5556 28540 5568
rect 27540 5528 28540 5556
rect 28534 5516 28540 5528
rect 28592 5516 28598 5568
rect 29546 5556 29552 5568
rect 29507 5528 29552 5556
rect 29546 5516 29552 5528
rect 29604 5556 29610 5568
rect 29914 5556 29920 5568
rect 29604 5528 29920 5556
rect 29604 5516 29610 5528
rect 29914 5516 29920 5528
rect 29972 5516 29978 5568
rect 30745 5559 30803 5565
rect 30745 5525 30757 5559
rect 30791 5556 30803 5559
rect 31110 5556 31116 5568
rect 30791 5528 31116 5556
rect 30791 5525 30803 5528
rect 30745 5519 30803 5525
rect 31110 5516 31116 5528
rect 31168 5516 31174 5568
rect 35360 5556 35388 5587
rect 37366 5556 37372 5568
rect 35360 5528 37372 5556
rect 37366 5516 37372 5528
rect 37424 5516 37430 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2409 5355 2467 5361
rect 2409 5352 2421 5355
rect 2372 5324 2421 5352
rect 2372 5312 2378 5324
rect 2409 5321 2421 5324
rect 2455 5321 2467 5355
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 2409 5315 2467 5321
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4614 5352 4620 5364
rect 4571 5324 4620 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5074 5352 5080 5364
rect 5031 5324 5080 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5534 5352 5540 5364
rect 5215 5324 5540 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 12713 5355 12771 5361
rect 12713 5321 12725 5355
rect 12759 5352 12771 5355
rect 21818 5352 21824 5364
rect 12759 5324 21824 5352
rect 12759 5321 12771 5324
rect 12713 5315 12771 5321
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 25406 5352 25412 5364
rect 25367 5324 25412 5352
rect 25406 5312 25412 5324
rect 25464 5312 25470 5364
rect 29086 5352 29092 5364
rect 25608 5324 29092 5352
rect 2222 5244 2228 5296
rect 2280 5284 2286 5296
rect 5721 5287 5779 5293
rect 2280 5256 4384 5284
rect 2280 5244 2286 5256
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3694 5216 3700 5228
rect 2832 5188 2877 5216
rect 3655 5188 3700 5216
rect 2832 5176 2838 5188
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 4356 5225 4384 5256
rect 5721 5253 5733 5287
rect 5767 5284 5779 5287
rect 5994 5284 6000 5296
rect 5767 5256 6000 5284
rect 5767 5253 5779 5256
rect 5721 5247 5779 5253
rect 5994 5244 6000 5256
rect 6052 5284 6058 5296
rect 6365 5287 6423 5293
rect 6365 5284 6377 5287
rect 6052 5256 6377 5284
rect 6052 5244 6058 5256
rect 6365 5253 6377 5256
rect 6411 5253 6423 5287
rect 6365 5247 6423 5253
rect 8389 5287 8447 5293
rect 8389 5253 8401 5287
rect 8435 5284 8447 5287
rect 8846 5284 8852 5296
rect 8435 5256 8852 5284
rect 8435 5253 8447 5256
rect 8389 5247 8447 5253
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 9766 5244 9772 5296
rect 9824 5284 9830 5296
rect 15930 5284 15936 5296
rect 9824 5256 12848 5284
rect 9824 5244 9830 5256
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 5350 5216 5356 5228
rect 4387 5188 5356 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5442 5176 5448 5228
rect 5500 5216 5506 5228
rect 6086 5216 6092 5228
rect 5500 5188 6092 5216
rect 5500 5176 5506 5188
rect 6086 5176 6092 5188
rect 6144 5216 6150 5228
rect 6549 5219 6607 5225
rect 6549 5216 6561 5219
rect 6144 5188 6561 5216
rect 6144 5176 6150 5188
rect 6549 5185 6561 5188
rect 6595 5185 6607 5219
rect 6730 5216 6736 5228
rect 6691 5188 6736 5216
rect 6549 5179 6607 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7558 5216 7564 5228
rect 7519 5188 7564 5216
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 8478 5216 8484 5228
rect 8036 5188 8484 5216
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5148 3111 5151
rect 3510 5148 3516 5160
rect 3099 5120 3516 5148
rect 3099 5117 3111 5120
rect 3053 5111 3111 5117
rect 3510 5108 3516 5120
rect 3568 5108 3574 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 7469 5151 7527 5157
rect 5307 5120 6592 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 6564 5092 6592 5120
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 7650 5148 7656 5160
rect 7515 5120 7656 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 8036 5157 8064 5188
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 9030 5216 9036 5228
rect 8991 5188 9036 5216
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 12820 5225 12848 5256
rect 15580 5256 15936 5284
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12406 5188 12633 5216
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5117 8079 5151
rect 8021 5111 8079 5117
rect 8110 5108 8116 5160
rect 8168 5148 8174 5160
rect 12406 5148 12434 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12805 5219 12863 5225
rect 12805 5185 12817 5219
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 14550 5216 14556 5228
rect 14332 5188 14556 5216
rect 14332 5176 14338 5188
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 15286 5216 15292 5228
rect 15247 5188 15292 5216
rect 15286 5176 15292 5188
rect 15344 5176 15350 5228
rect 15470 5216 15476 5228
rect 15431 5188 15476 5216
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 15580 5225 15608 5256
rect 15930 5244 15936 5256
rect 15988 5244 15994 5296
rect 19337 5287 19395 5293
rect 19337 5284 19349 5287
rect 18432 5256 19349 5284
rect 15565 5219 15623 5225
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 15565 5179 15623 5185
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15657 5179 15715 5185
rect 8168 5120 12434 5148
rect 8168 5108 8174 5120
rect 13446 5108 13452 5160
rect 13504 5148 13510 5160
rect 15672 5148 15700 5179
rect 18046 5176 18052 5228
rect 18104 5216 18110 5228
rect 18432 5225 18460 5256
rect 19337 5253 19349 5256
rect 19383 5253 19395 5287
rect 19337 5247 19395 5253
rect 19426 5244 19432 5296
rect 19484 5284 19490 5296
rect 19705 5287 19763 5293
rect 19705 5284 19717 5287
rect 19484 5256 19717 5284
rect 19484 5244 19490 5256
rect 19705 5253 19717 5256
rect 19751 5253 19763 5287
rect 19705 5247 19763 5253
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 18104 5188 18245 5216
rect 18104 5176 18110 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18417 5219 18475 5225
rect 18417 5185 18429 5219
rect 18463 5185 18475 5219
rect 18417 5179 18475 5185
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5185 18567 5219
rect 18509 5179 18567 5185
rect 13504 5120 15700 5148
rect 13504 5108 13510 5120
rect 18322 5108 18328 5160
rect 18380 5148 18386 5160
rect 18524 5148 18552 5179
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 19521 5219 19579 5225
rect 18656 5188 18701 5216
rect 18656 5176 18662 5188
rect 19521 5185 19533 5219
rect 19567 5216 19579 5219
rect 21358 5216 21364 5228
rect 19567 5188 21364 5216
rect 19567 5185 19579 5188
rect 19521 5179 19579 5185
rect 21358 5176 21364 5188
rect 21416 5176 21422 5228
rect 18380 5120 18552 5148
rect 18380 5108 18386 5120
rect 21082 5108 21088 5160
rect 21140 5148 21146 5160
rect 25608 5148 25636 5324
rect 29086 5312 29092 5324
rect 29144 5312 29150 5364
rect 29730 5352 29736 5364
rect 29643 5324 29736 5352
rect 29730 5312 29736 5324
rect 29788 5352 29794 5364
rect 30742 5352 30748 5364
rect 29788 5324 30748 5352
rect 29788 5312 29794 5324
rect 26418 5284 26424 5296
rect 26331 5256 26424 5284
rect 26418 5244 26424 5256
rect 26476 5284 26482 5296
rect 27890 5284 27896 5296
rect 26476 5256 27896 5284
rect 26476 5244 26482 5256
rect 27264 5225 27292 5256
rect 27890 5244 27896 5256
rect 27948 5244 27954 5296
rect 27249 5219 27307 5225
rect 27249 5185 27261 5219
rect 27295 5185 27307 5219
rect 27249 5179 27307 5185
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5185 27399 5219
rect 27341 5179 27399 5185
rect 21140 5120 25636 5148
rect 21140 5108 21146 5120
rect 27356 5092 27384 5179
rect 27430 5176 27436 5228
rect 27488 5216 27494 5228
rect 27617 5219 27675 5225
rect 27488 5188 27533 5216
rect 27488 5176 27494 5188
rect 27617 5185 27629 5219
rect 27663 5216 27675 5219
rect 28166 5216 28172 5228
rect 27663 5188 28172 5216
rect 27663 5185 27675 5188
rect 27617 5179 27675 5185
rect 28166 5176 28172 5188
rect 28224 5176 28230 5228
rect 30098 5176 30104 5228
rect 30156 5216 30162 5228
rect 30193 5219 30251 5225
rect 30193 5216 30205 5219
rect 30156 5188 30205 5216
rect 30156 5176 30162 5188
rect 30193 5185 30205 5188
rect 30239 5185 30251 5219
rect 30374 5216 30380 5228
rect 30335 5188 30380 5216
rect 30193 5179 30251 5185
rect 30374 5176 30380 5188
rect 30432 5176 30438 5228
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5185 30527 5219
rect 30469 5179 30527 5185
rect 30581 5219 30639 5225
rect 30581 5185 30593 5219
rect 30627 5216 30639 5219
rect 30668 5216 30696 5324
rect 30742 5312 30748 5324
rect 30800 5312 30806 5364
rect 31662 5312 31668 5364
rect 31720 5352 31726 5364
rect 32217 5355 32275 5361
rect 32217 5352 32229 5355
rect 31720 5324 32229 5352
rect 31720 5312 31726 5324
rect 32217 5321 32229 5324
rect 32263 5321 32275 5355
rect 32217 5315 32275 5321
rect 36262 5312 36268 5364
rect 36320 5352 36326 5364
rect 37277 5355 37335 5361
rect 37277 5352 37289 5355
rect 36320 5324 37289 5352
rect 36320 5312 36326 5324
rect 37277 5321 37289 5324
rect 37323 5321 37335 5355
rect 37277 5315 37335 5321
rect 37918 5244 37924 5296
rect 37976 5284 37982 5296
rect 37976 5256 38700 5284
rect 37976 5244 37982 5256
rect 30627 5188 30696 5216
rect 30627 5185 30639 5188
rect 30581 5179 30639 5185
rect 30006 5108 30012 5160
rect 30064 5148 30070 5160
rect 30484 5148 30512 5179
rect 38378 5176 38384 5228
rect 38436 5225 38442 5228
rect 38672 5225 38700 5256
rect 38436 5216 38448 5225
rect 38657 5219 38715 5225
rect 38436 5188 38481 5216
rect 38436 5179 38448 5188
rect 38657 5185 38669 5219
rect 38703 5185 38715 5219
rect 38657 5179 38715 5185
rect 38436 5176 38442 5179
rect 30064 5120 30512 5148
rect 30064 5108 30070 5120
rect 53742 5108 53748 5160
rect 53800 5148 53806 5160
rect 54389 5151 54447 5157
rect 54389 5148 54401 5151
rect 53800 5120 54401 5148
rect 53800 5108 53806 5120
rect 54389 5117 54401 5120
rect 54435 5117 54447 5151
rect 54389 5111 54447 5117
rect 5718 5080 5724 5092
rect 5679 5052 5724 5080
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 6546 5040 6552 5092
rect 6604 5040 6610 5092
rect 8849 5083 8907 5089
rect 8849 5080 8861 5083
rect 7944 5052 8861 5080
rect 1949 5015 2007 5021
rect 1949 4981 1961 5015
rect 1995 5012 2007 5015
rect 3510 5012 3516 5024
rect 1995 4984 3516 5012
rect 1995 4981 2007 4984
rect 1949 4975 2007 4981
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 3878 5012 3884 5024
rect 3839 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 7944 5021 7972 5052
rect 8849 5049 8861 5052
rect 8895 5049 8907 5083
rect 8849 5043 8907 5049
rect 15933 5083 15991 5089
rect 15933 5049 15945 5083
rect 15979 5080 15991 5083
rect 16942 5080 16948 5092
rect 15979 5052 16948 5080
rect 15979 5049 15991 5052
rect 15933 5043 15991 5049
rect 16942 5040 16948 5052
rect 17000 5040 17006 5092
rect 18877 5083 18935 5089
rect 18877 5049 18889 5083
rect 18923 5080 18935 5083
rect 19426 5080 19432 5092
rect 18923 5052 19432 5080
rect 18923 5049 18935 5052
rect 18877 5043 18935 5049
rect 19426 5040 19432 5052
rect 19484 5040 19490 5092
rect 22094 5040 22100 5092
rect 22152 5080 22158 5092
rect 23293 5083 23351 5089
rect 23293 5080 23305 5083
rect 22152 5052 23305 5080
rect 22152 5040 22158 5052
rect 23293 5049 23305 5052
rect 23339 5049 23351 5083
rect 23293 5043 23351 5049
rect 27338 5040 27344 5092
rect 27396 5040 27402 5092
rect 54110 5040 54116 5092
rect 54168 5080 54174 5092
rect 55033 5083 55091 5089
rect 55033 5080 55045 5083
rect 54168 5052 55045 5080
rect 54168 5040 54174 5052
rect 55033 5049 55045 5052
rect 55079 5049 55091 5083
rect 55033 5043 55091 5049
rect 7929 5015 7987 5021
rect 7929 5012 7941 5015
rect 6788 4984 7941 5012
rect 6788 4972 6794 4984
rect 7929 4981 7941 4984
rect 7975 4981 7987 5015
rect 7929 4975 7987 4981
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 10226 5012 10232 5024
rect 9723 4984 10232 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10778 5012 10784 5024
rect 10367 4984 10784 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 10965 5015 11023 5021
rect 10965 4981 10977 5015
rect 11011 5012 11023 5015
rect 11330 5012 11336 5024
rect 11011 4984 11336 5012
rect 11011 4981 11023 4984
rect 10965 4975 11023 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 11977 5015 12035 5021
rect 11977 5012 11989 5015
rect 11940 4984 11989 5012
rect 11940 4972 11946 4984
rect 11977 4981 11989 4984
rect 12023 4981 12035 5015
rect 11977 4975 12035 4981
rect 13449 5015 13507 5021
rect 13449 4981 13461 5015
rect 13495 5012 13507 5015
rect 13814 5012 13820 5024
rect 13495 4984 13820 5012
rect 13495 4981 13507 4984
rect 13449 4975 13507 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14090 5012 14096 5024
rect 14051 4984 14096 5012
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 14734 5012 14740 5024
rect 14695 4984 14740 5012
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 16758 4972 16764 5024
rect 16816 5012 16822 5024
rect 16853 5015 16911 5021
rect 16853 5012 16865 5015
rect 16816 4984 16865 5012
rect 16816 4972 16822 4984
rect 16853 4981 16865 4984
rect 16899 4981 16911 5015
rect 16853 4975 16911 4981
rect 17773 5015 17831 5021
rect 17773 4981 17785 5015
rect 17819 5012 17831 5015
rect 18414 5012 18420 5024
rect 17819 4984 18420 5012
rect 17819 4981 17831 4984
rect 17773 4975 17831 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 20165 5015 20223 5021
rect 20165 5012 20177 5015
rect 20128 4984 20177 5012
rect 20128 4972 20134 4984
rect 20165 4981 20177 4984
rect 20211 4981 20223 5015
rect 20165 4975 20223 4981
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20956 4984 21005 5012
rect 20956 4972 20962 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 21726 4972 21732 5024
rect 21784 5012 21790 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21784 4984 21833 5012
rect 21784 4972 21790 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 21821 4975 21879 4981
rect 22554 4972 22560 5024
rect 22612 5012 22618 5024
rect 22649 5015 22707 5021
rect 22649 5012 22661 5015
rect 22612 4984 22661 5012
rect 22612 4972 22618 4984
rect 22649 4981 22661 4984
rect 22695 4981 22707 5015
rect 22649 4975 22707 4981
rect 23474 4972 23480 5024
rect 23532 5012 23538 5024
rect 23845 5015 23903 5021
rect 23845 5012 23857 5015
rect 23532 4984 23857 5012
rect 23532 4972 23538 4984
rect 23845 4981 23857 4984
rect 23891 4981 23903 5015
rect 23845 4975 23903 4981
rect 26973 5015 27031 5021
rect 26973 4981 26985 5015
rect 27019 5012 27031 5015
rect 27246 5012 27252 5024
rect 27019 4984 27252 5012
rect 27019 4981 27031 4984
rect 26973 4975 27031 4981
rect 27246 4972 27252 4984
rect 27304 4972 27310 5024
rect 30834 5012 30840 5024
rect 30795 4984 30840 5012
rect 30834 4972 30840 4984
rect 30892 4972 30898 5024
rect 53650 4972 53656 5024
rect 53708 5012 53714 5024
rect 53745 5015 53803 5021
rect 53745 5012 53757 5015
rect 53708 4984 53757 5012
rect 53708 4972 53714 4984
rect 53745 4981 53757 4984
rect 53791 4981 53803 5015
rect 58158 5012 58164 5024
rect 58119 4984 58164 5012
rect 53745 4975 53803 4981
rect 58158 4972 58164 4984
rect 58216 4972 58222 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 2746 4780 6040 4808
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 2746 4740 2774 4780
rect 2363 4712 2774 4740
rect 4985 4743 5043 4749
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 4985 4709 4997 4743
rect 5031 4740 5043 4743
rect 5902 4740 5908 4752
rect 5031 4712 5908 4740
rect 5031 4709 5043 4712
rect 4985 4703 5043 4709
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 6012 4740 6040 4780
rect 6086 4768 6092 4820
rect 6144 4808 6150 4820
rect 7466 4808 7472 4820
rect 6144 4780 6189 4808
rect 7427 4780 7472 4808
rect 6144 4768 6150 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7745 4811 7803 4817
rect 7745 4777 7757 4811
rect 7791 4808 7803 4811
rect 8110 4808 8116 4820
rect 7791 4780 8116 4808
rect 7791 4777 7803 4780
rect 7745 4771 7803 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 8220 4780 8953 4808
rect 7006 4740 7012 4752
rect 6012 4712 7012 4740
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 7484 4740 7512 4768
rect 8220 4740 8248 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 9398 4808 9404 4820
rect 9359 4780 9404 4808
rect 8941 4771 8999 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 9824 4780 10241 4808
rect 9824 4768 9830 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 10229 4771 10287 4777
rect 22465 4811 22523 4817
rect 22465 4777 22477 4811
rect 22511 4808 22523 4811
rect 23842 4808 23848 4820
rect 22511 4780 23848 4808
rect 22511 4777 22523 4780
rect 22465 4771 22523 4777
rect 23842 4768 23848 4780
rect 23900 4768 23906 4820
rect 24394 4808 24400 4820
rect 24355 4780 24400 4808
rect 24394 4768 24400 4780
rect 24452 4768 24458 4820
rect 46750 4808 46756 4820
rect 24504 4780 46756 4808
rect 7484 4712 8248 4740
rect 8389 4743 8447 4749
rect 8389 4709 8401 4743
rect 8435 4740 8447 4743
rect 9858 4740 9864 4752
rect 8435 4712 9864 4740
rect 8435 4709 8447 4712
rect 8389 4703 8447 4709
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 10134 4700 10140 4752
rect 10192 4740 10198 4752
rect 10597 4743 10655 4749
rect 10597 4740 10609 4743
rect 10192 4712 10609 4740
rect 10192 4700 10198 4712
rect 10597 4709 10609 4712
rect 10643 4709 10655 4743
rect 10597 4703 10655 4709
rect 16761 4743 16819 4749
rect 16761 4709 16773 4743
rect 16807 4740 16819 4743
rect 18138 4740 18144 4752
rect 16807 4712 18144 4740
rect 16807 4709 16819 4712
rect 16761 4703 16819 4709
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 21361 4743 21419 4749
rect 21361 4709 21373 4743
rect 21407 4740 21419 4743
rect 22002 4740 22008 4752
rect 21407 4712 22008 4740
rect 21407 4709 21419 4712
rect 21361 4703 21419 4709
rect 22002 4700 22008 4712
rect 22060 4700 22066 4752
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 7469 4675 7527 4681
rect 7469 4672 7481 4675
rect 5776 4644 7481 4672
rect 5776 4632 5782 4644
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3007 4576 3985 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5258 4604 5264 4616
rect 5215 4576 5264 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 1765 4539 1823 4545
rect 1765 4505 1777 4539
rect 1811 4536 1823 4539
rect 4172 4536 4200 4567
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 6012 4613 6040 4644
rect 7469 4641 7481 4644
rect 7515 4672 7527 4675
rect 8478 4672 8484 4684
rect 7515 4644 8484 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 8478 4632 8484 4644
rect 8536 4672 8542 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8536 4644 9045 4672
rect 8536 4632 8542 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 10505 4675 10563 4681
rect 10505 4672 10517 4675
rect 10468 4644 10517 4672
rect 10468 4632 10474 4644
rect 10505 4641 10517 4644
rect 10551 4641 10563 4675
rect 10505 4635 10563 4641
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4672 12955 4675
rect 13446 4672 13452 4684
rect 12943 4644 13452 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 18966 4672 18972 4684
rect 18095 4644 18972 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 24504 4672 24532 4780
rect 46750 4768 46756 4780
rect 46808 4768 46814 4820
rect 32122 4700 32128 4752
rect 32180 4740 32186 4752
rect 32401 4743 32459 4749
rect 32401 4740 32413 4743
rect 32180 4712 32413 4740
rect 32180 4700 32186 4712
rect 32401 4709 32413 4712
rect 32447 4709 32459 4743
rect 32401 4703 32459 4709
rect 52178 4700 52184 4752
rect 52236 4740 52242 4752
rect 52825 4743 52883 4749
rect 52825 4740 52837 4743
rect 52236 4712 52837 4740
rect 52236 4700 52242 4712
rect 52825 4709 52837 4712
rect 52871 4709 52883 4743
rect 52825 4703 52883 4709
rect 53926 4700 53932 4752
rect 53984 4740 53990 4752
rect 55309 4743 55367 4749
rect 55309 4740 55321 4743
rect 53984 4712 55321 4740
rect 53984 4700 53990 4712
rect 55309 4709 55321 4712
rect 55355 4709 55367 4743
rect 55309 4703 55367 4709
rect 23768 4644 24532 4672
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5592 4576 5641 4604
rect 5592 4564 5598 4576
rect 5629 4573 5641 4576
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4573 6055 4607
rect 6178 4604 6184 4616
rect 6139 4576 6184 4604
rect 5997 4567 6055 4573
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 6788 4576 7113 4604
rect 6788 4564 6794 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7558 4604 7564 4616
rect 7519 4576 7564 4604
rect 7101 4567 7159 4573
rect 6546 4536 6552 4548
rect 1811 4508 4108 4536
rect 4172 4508 6552 4536
rect 1811 4505 1823 4508
rect 1765 4499 1823 4505
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 4080 4468 4108 4508
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 6822 4496 6828 4548
rect 6880 4536 6886 4548
rect 7116 4536 7144 4567
rect 7558 4564 7564 4576
rect 7616 4604 7622 4616
rect 9122 4604 9128 4616
rect 7616 4576 9128 4604
rect 7616 4564 7622 4576
rect 9122 4564 9128 4576
rect 9180 4604 9186 4616
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 9180 4576 9229 4604
rect 9180 4564 9186 4576
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 10726 4607 10784 4613
rect 10726 4604 10738 4607
rect 9217 4567 9275 4573
rect 9600 4576 10738 4604
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 6880 4508 7052 4536
rect 7116 4508 8953 4536
rect 6880 4496 6886 4508
rect 5258 4468 5264 4480
rect 2832 4440 2877 4468
rect 4080 4440 5264 4468
rect 2832 4428 2838 4440
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 5813 4471 5871 4477
rect 5813 4437 5825 4471
rect 5859 4468 5871 4471
rect 6914 4468 6920 4480
rect 5859 4440 6920 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7024 4468 7052 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 9600 4468 9628 4576
rect 10726 4573 10738 4576
rect 10772 4604 10784 4607
rect 10962 4604 10968 4616
rect 10772 4576 10968 4604
rect 10772 4573 10784 4576
rect 10726 4567 10784 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4604 11667 4607
rect 12158 4604 12164 4616
rect 11655 4576 12164 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 12253 4607 12311 4613
rect 12253 4573 12265 4607
rect 12299 4604 12311 4607
rect 12986 4604 12992 4616
rect 12299 4576 12992 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13357 4607 13415 4613
rect 13357 4573 13369 4607
rect 13403 4604 13415 4607
rect 13906 4604 13912 4616
rect 13403 4576 13912 4604
rect 13403 4573 13415 4576
rect 13357 4567 13415 4573
rect 13906 4564 13912 4576
rect 13964 4604 13970 4616
rect 14182 4604 14188 4616
rect 13964 4576 14188 4604
rect 13964 4564 13970 4576
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4604 14887 4607
rect 15378 4604 15384 4616
rect 14875 4576 15384 4604
rect 14875 4573 14887 4576
rect 14829 4567 14887 4573
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4604 15531 4607
rect 16022 4604 16028 4616
rect 15519 4576 16028 4604
rect 15519 4573 15531 4576
rect 15473 4567 15531 4573
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 16117 4607 16175 4613
rect 16117 4573 16129 4607
rect 16163 4604 16175 4607
rect 16482 4604 16488 4616
rect 16163 4576 16488 4604
rect 16163 4573 16175 4576
rect 16117 4567 16175 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 17402 4604 17408 4616
rect 17363 4576 17408 4604
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 19150 4604 19156 4616
rect 18739 4576 19156 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19392 4576 19441 4604
rect 19392 4564 19398 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4604 20131 4607
rect 20622 4604 20628 4616
rect 20119 4576 20628 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 20717 4607 20775 4613
rect 20717 4573 20729 4607
rect 20763 4604 20775 4607
rect 21174 4604 21180 4616
rect 20763 4576 21180 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 21174 4564 21180 4576
rect 21232 4564 21238 4616
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 22278 4604 22284 4616
rect 22051 4576 22284 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22278 4564 22284 4576
rect 22336 4564 22342 4616
rect 23566 4564 23572 4616
rect 23624 4613 23630 4616
rect 23624 4604 23636 4613
rect 23624 4576 23669 4604
rect 23624 4567 23636 4576
rect 23624 4564 23630 4567
rect 10594 4496 10600 4548
rect 10652 4536 10658 4548
rect 10870 4536 10876 4548
rect 10652 4508 10876 4536
rect 10652 4496 10658 4508
rect 10870 4496 10876 4508
rect 10928 4496 10934 4548
rect 22370 4496 22376 4548
rect 22428 4536 22434 4548
rect 23768 4536 23796 4644
rect 53190 4632 53196 4684
rect 53248 4672 53254 4684
rect 54113 4675 54171 4681
rect 54113 4672 54125 4675
rect 53248 4644 54125 4672
rect 53248 4632 53254 4644
rect 54113 4641 54125 4644
rect 54159 4641 54171 4675
rect 54113 4635 54171 4641
rect 54294 4632 54300 4684
rect 54352 4672 54358 4684
rect 55953 4675 56011 4681
rect 55953 4672 55965 4675
rect 54352 4644 55965 4672
rect 54352 4632 54358 4644
rect 55953 4641 55965 4644
rect 55999 4641 56011 4675
rect 55953 4635 56011 4641
rect 23845 4607 23903 4613
rect 23845 4573 23857 4607
rect 23891 4604 23903 4607
rect 25130 4604 25136 4616
rect 23891 4576 25136 4604
rect 23891 4573 23903 4576
rect 23845 4567 23903 4573
rect 25130 4564 25136 4576
rect 25188 4604 25194 4616
rect 25774 4604 25780 4616
rect 25188 4576 25780 4604
rect 25188 4564 25194 4576
rect 25774 4564 25780 4576
rect 25832 4564 25838 4616
rect 30926 4564 30932 4616
rect 30984 4604 30990 4616
rect 31021 4607 31079 4613
rect 31021 4604 31033 4607
rect 30984 4576 31033 4604
rect 30984 4564 30990 4576
rect 31021 4573 31033 4576
rect 31067 4573 31079 4607
rect 31021 4567 31079 4573
rect 31110 4564 31116 4616
rect 31168 4604 31174 4616
rect 31277 4607 31335 4613
rect 31277 4604 31289 4607
rect 31168 4576 31289 4604
rect 31168 4564 31174 4576
rect 31277 4573 31289 4576
rect 31323 4573 31335 4607
rect 31277 4567 31335 4573
rect 52086 4564 52092 4616
rect 52144 4604 52150 4616
rect 52181 4607 52239 4613
rect 52181 4604 52193 4607
rect 52144 4576 52193 4604
rect 52144 4564 52150 4576
rect 52181 4573 52193 4576
rect 52227 4573 52239 4607
rect 52181 4567 52239 4573
rect 52638 4564 52644 4616
rect 52696 4604 52702 4616
rect 53469 4607 53527 4613
rect 53469 4604 53481 4607
rect 52696 4576 53481 4604
rect 52696 4564 52702 4576
rect 53469 4573 53481 4576
rect 53515 4573 53527 4607
rect 53469 4567 53527 4573
rect 22428 4508 23796 4536
rect 22428 4496 22434 4508
rect 25038 4496 25044 4548
rect 25096 4536 25102 4548
rect 25510 4539 25568 4545
rect 25510 4536 25522 4539
rect 25096 4508 25522 4536
rect 25096 4496 25102 4508
rect 25510 4505 25522 4508
rect 25556 4505 25568 4539
rect 25510 4499 25568 4505
rect 7024 4440 9628 4468
rect 13541 4471 13599 4477
rect 13541 4437 13553 4471
rect 13587 4468 13599 4471
rect 13998 4468 14004 4480
rect 13587 4440 14004 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 14185 4471 14243 4477
rect 14185 4437 14197 4471
rect 14231 4468 14243 4471
rect 18322 4468 18328 4480
rect 14231 4440 18328 4468
rect 14231 4437 14243 4440
rect 14185 4431 14243 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 3602 4224 3608 4276
rect 3660 4264 3666 4276
rect 4062 4264 4068 4276
rect 3660 4236 4068 4264
rect 3660 4224 3666 4236
rect 4062 4224 4068 4236
rect 4120 4264 4126 4276
rect 6270 4264 6276 4276
rect 4120 4236 6276 4264
rect 4120 4224 4126 4236
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 6733 4267 6791 4273
rect 6733 4233 6745 4267
rect 6779 4264 6791 4267
rect 7098 4264 7104 4276
rect 6779 4236 7104 4264
rect 6779 4233 6791 4236
rect 6733 4227 6791 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 9398 4224 9404 4276
rect 9456 4264 9462 4276
rect 29730 4264 29736 4276
rect 9456 4236 29736 4264
rect 9456 4224 9462 4236
rect 29730 4224 29736 4236
rect 29788 4224 29794 4276
rect 3878 4156 3884 4208
rect 3936 4196 3942 4208
rect 6365 4199 6423 4205
rect 6365 4196 6377 4199
rect 3936 4168 6377 4196
rect 3936 4156 3942 4168
rect 6365 4165 6377 4168
rect 6411 4165 6423 4199
rect 6546 4196 6552 4208
rect 6507 4168 6552 4196
rect 6365 4159 6423 4165
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 10520 4168 10732 4196
rect 1762 4088 1768 4140
rect 1820 4128 1826 4140
rect 2590 4128 2596 4140
rect 1820 4100 2596 4128
rect 1820 4088 1826 4100
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3786 4128 3792 4140
rect 3559 4100 3792 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 4062 4128 4068 4140
rect 4023 4100 4068 4128
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4614 4128 4620 4140
rect 4295 4100 4620 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 4614 4088 4620 4100
rect 4672 4088 4678 4140
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 7466 4128 7472 4140
rect 5859 4100 7472 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2130 3924 2136 3936
rect 2091 3896 2136 3924
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 2777 3927 2835 3933
rect 2777 3893 2789 3927
rect 2823 3924 2835 3927
rect 3234 3924 3240 3936
rect 2823 3896 3240 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3329 3927 3387 3933
rect 3329 3893 3341 3927
rect 3375 3924 3387 3927
rect 4614 3924 4620 3936
rect 3375 3896 4620 3924
rect 3375 3893 3387 3896
rect 3329 3887 3387 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4798 3924 4804 3936
rect 4759 3896 4804 3924
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5000 3924 5028 4091
rect 7466 4088 7472 4100
rect 7524 4128 7530 4140
rect 7837 4131 7895 4137
rect 7837 4128 7849 4131
rect 7524 4100 7849 4128
rect 7524 4088 7530 4100
rect 7837 4097 7849 4100
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6822 4060 6828 4072
rect 5767 4032 6828 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 8386 4060 8392 4072
rect 7432 4032 7604 4060
rect 8347 4032 8392 4060
rect 7432 4020 7438 4032
rect 7466 3992 7472 4004
rect 5828 3964 7472 3992
rect 5074 3924 5080 3936
rect 5000 3896 5080 3924
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5445 3927 5503 3933
rect 5445 3893 5457 3927
rect 5491 3924 5503 3927
rect 5534 3924 5540 3936
rect 5491 3896 5540 3924
rect 5491 3893 5503 3896
rect 5445 3887 5503 3893
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5828 3933 5856 3964
rect 7466 3952 7472 3964
rect 7524 3952 7530 4004
rect 7576 3936 7604 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8570 4060 8576 4072
rect 8531 4032 8576 4060
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9508 4060 9536 4091
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 10008 4100 10057 4128
rect 10008 4088 10014 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10520 4128 10548 4168
rect 10045 4091 10103 4097
rect 10336 4100 10548 4128
rect 10704 4128 10732 4168
rect 16776 4168 17080 4196
rect 11514 4128 11520 4140
rect 10704 4100 11520 4128
rect 10336 4060 10364 4100
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 11698 4128 11704 4140
rect 11659 4100 11704 4128
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 12069 4131 12127 4137
rect 12069 4128 12081 4131
rect 11808 4100 12081 4128
rect 9508 4032 10364 4060
rect 10410 4020 10416 4072
rect 10468 4060 10474 4072
rect 10962 4060 10968 4072
rect 10468 4032 10513 4060
rect 10923 4032 10968 4060
rect 10468 4020 10474 4032
rect 10962 4020 10968 4032
rect 11020 4060 11026 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11020 4032 11621 4060
rect 11020 4020 11026 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 11609 4023 11667 4029
rect 8294 3992 8300 4004
rect 8255 3964 8300 3992
rect 8294 3952 8300 3964
rect 8352 3952 8358 4004
rect 10594 3992 10600 4004
rect 10555 3964 10600 3992
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 10686 3952 10692 4004
rect 10744 3992 10750 4004
rect 11808 3992 11836 4100
rect 12069 4097 12081 4100
rect 12115 4097 12127 4131
rect 12069 4091 12127 4097
rect 12250 4088 12256 4140
rect 12308 4128 12314 4140
rect 13357 4131 13415 4137
rect 13357 4128 13369 4131
rect 12308 4100 13369 4128
rect 12308 4088 12314 4100
rect 13357 4097 13369 4100
rect 13403 4128 13415 4131
rect 14274 4128 14280 4140
rect 13403 4100 14280 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 15562 4088 15568 4140
rect 15620 4128 15626 4140
rect 16669 4131 16727 4137
rect 16669 4128 16681 4131
rect 15620 4100 16681 4128
rect 15620 4088 15626 4100
rect 16669 4097 16681 4100
rect 16715 4128 16727 4131
rect 16776 4128 16804 4168
rect 16942 4137 16948 4140
rect 16936 4128 16948 4137
rect 16715 4100 16804 4128
rect 16903 4100 16948 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 16936 4091 16948 4100
rect 16942 4088 16948 4091
rect 17000 4088 17006 4140
rect 17052 4128 17080 4168
rect 19426 4156 19432 4208
rect 19484 4196 19490 4208
rect 27246 4205 27252 4208
rect 27240 4196 27252 4205
rect 19484 4168 19656 4196
rect 27207 4168 27252 4196
rect 19484 4156 19490 4168
rect 19242 4128 19248 4140
rect 17052 4100 19248 4128
rect 19242 4088 19248 4100
rect 19300 4128 19306 4140
rect 19521 4131 19579 4137
rect 19521 4128 19533 4131
rect 19300 4100 19533 4128
rect 19300 4088 19306 4100
rect 19521 4097 19533 4100
rect 19567 4097 19579 4131
rect 19628 4128 19656 4168
rect 27240 4159 27252 4168
rect 27246 4156 27252 4159
rect 27304 4156 27310 4208
rect 19777 4131 19835 4137
rect 19777 4128 19789 4131
rect 19628 4100 19789 4128
rect 19521 4091 19579 4097
rect 19777 4097 19789 4100
rect 19823 4097 19835 4131
rect 19777 4091 19835 4097
rect 25774 4088 25780 4140
rect 25832 4128 25838 4140
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 25832 4100 26985 4128
rect 25832 4088 25838 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 30926 4088 30932 4140
rect 30984 4128 30990 4140
rect 33870 4128 33876 4140
rect 30984 4100 33876 4128
rect 30984 4088 30990 4100
rect 33870 4088 33876 4100
rect 33928 4128 33934 4140
rect 34609 4131 34667 4137
rect 34609 4128 34621 4131
rect 33928 4100 34621 4128
rect 33928 4088 33934 4100
rect 34609 4097 34621 4100
rect 34655 4097 34667 4131
rect 34609 4091 34667 4097
rect 34698 4088 34704 4140
rect 34756 4128 34762 4140
rect 34865 4131 34923 4137
rect 34865 4128 34877 4131
rect 34756 4100 34877 4128
rect 34756 4088 34762 4100
rect 34865 4097 34877 4100
rect 34911 4097 34923 4131
rect 34865 4091 34923 4097
rect 53006 4088 53012 4140
rect 53064 4128 53070 4140
rect 54665 4131 54723 4137
rect 54665 4128 54677 4131
rect 53064 4100 54677 4128
rect 53064 4088 53070 4100
rect 54665 4097 54677 4100
rect 54711 4097 54723 4131
rect 54665 4091 54723 4097
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4060 14887 4063
rect 16206 4060 16212 4072
rect 14875 4032 16212 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 51810 4020 51816 4072
rect 51868 4060 51874 4072
rect 52733 4063 52791 4069
rect 52733 4060 52745 4063
rect 51868 4032 52745 4060
rect 51868 4020 51874 4032
rect 52733 4029 52745 4032
rect 52779 4029 52791 4063
rect 52733 4023 52791 4029
rect 54018 4020 54024 4072
rect 54076 4060 54082 4072
rect 55953 4063 56011 4069
rect 55953 4060 55965 4063
rect 54076 4032 55965 4060
rect 54076 4020 54082 4032
rect 55953 4029 55965 4032
rect 55999 4029 56011 4063
rect 55953 4023 56011 4029
rect 10744 3964 11836 3992
rect 12897 3995 12955 4001
rect 10744 3952 10750 3964
rect 12897 3961 12909 3995
rect 12943 3992 12955 3995
rect 14185 3995 14243 4001
rect 12943 3964 14136 3992
rect 12943 3961 12955 3964
rect 12897 3955 12955 3961
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3893 5871 3927
rect 5813 3887 5871 3893
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3924 6607 3927
rect 6638 3924 6644 3936
rect 6595 3896 6644 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 6638 3884 6644 3896
rect 6696 3884 6702 3936
rect 7374 3924 7380 3936
rect 7335 3896 7380 3924
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 7558 3884 7564 3936
rect 7616 3884 7622 3936
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 8478 3924 8484 3936
rect 8251 3896 8484 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 8478 3884 8484 3896
rect 8536 3924 8542 3936
rect 9030 3924 9036 3936
rect 8536 3896 9036 3924
rect 8536 3884 8542 3896
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9122 3884 9128 3936
rect 9180 3924 9186 3936
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 9180 3896 9321 3924
rect 9180 3884 9186 3896
rect 9309 3893 9321 3896
rect 9355 3893 9367 3927
rect 9309 3887 9367 3893
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10192 3896 10517 3924
rect 10192 3884 10198 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10505 3887 10563 3893
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 12032 3896 12081 3924
rect 12032 3884 12038 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12069 3887 12127 3893
rect 12253 3927 12311 3933
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 13170 3924 13176 3936
rect 12299 3896 13176 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 13538 3924 13544 3936
rect 13499 3896 13544 3924
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 14108 3924 14136 3964
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 15194 3992 15200 4004
rect 14231 3964 15200 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 15473 3995 15531 4001
rect 15473 3961 15485 3995
rect 15519 3992 15531 3995
rect 16666 3992 16672 4004
rect 15519 3964 16672 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 18049 3995 18107 4001
rect 18049 3961 18061 3995
rect 18095 3992 18107 3995
rect 18506 3992 18512 4004
rect 18095 3964 18512 3992
rect 18095 3961 18107 3964
rect 18049 3955 18107 3961
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 20901 3995 20959 4001
rect 20901 3961 20913 3995
rect 20947 3992 20959 3995
rect 21358 3992 21364 4004
rect 20947 3964 21364 3992
rect 20947 3961 20959 3964
rect 20901 3955 20959 3961
rect 21358 3952 21364 3964
rect 21416 3952 21422 4004
rect 22462 3952 22468 4004
rect 22520 3992 22526 4004
rect 24949 3995 25007 4001
rect 24949 3992 24961 3995
rect 22520 3964 24961 3992
rect 22520 3952 22526 3964
rect 24949 3961 24961 3964
rect 24995 3961 25007 3995
rect 24949 3955 25007 3961
rect 28353 3995 28411 4001
rect 28353 3961 28365 3995
rect 28399 3992 28411 3995
rect 28534 3992 28540 4004
rect 28399 3964 28540 3992
rect 28399 3961 28411 3964
rect 28353 3955 28411 3961
rect 28534 3952 28540 3964
rect 28592 3952 28598 4004
rect 35618 3952 35624 4004
rect 35676 3992 35682 4004
rect 35989 3995 36047 4001
rect 35989 3992 36001 3995
rect 35676 3964 36001 3992
rect 35676 3952 35682 3964
rect 35989 3961 36001 3964
rect 36035 3961 36047 3995
rect 35989 3955 36047 3961
rect 52822 3952 52828 4004
rect 52880 3992 52886 4004
rect 52880 3964 54064 3992
rect 52880 3952 52886 3964
rect 15930 3924 15936 3936
rect 14108 3896 15936 3924
rect 15930 3884 15936 3896
rect 15988 3884 15994 3936
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 17678 3924 17684 3936
rect 16163 3896 17684 3924
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3924 19119 3927
rect 19426 3924 19432 3936
rect 19107 3896 19432 3924
rect 19107 3893 19119 3896
rect 19061 3887 19119 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 22373 3927 22431 3933
rect 22373 3893 22385 3927
rect 22419 3924 22431 3927
rect 22922 3924 22928 3936
rect 22419 3896 22928 3924
rect 22419 3893 22431 3896
rect 22373 3887 22431 3893
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 23017 3927 23075 3933
rect 23017 3893 23029 3927
rect 23063 3924 23075 3927
rect 23106 3924 23112 3936
rect 23063 3896 23112 3924
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 23106 3884 23112 3896
rect 23164 3884 23170 3936
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 23477 3927 23535 3933
rect 23477 3924 23489 3927
rect 23440 3896 23489 3924
rect 23440 3884 23446 3896
rect 23477 3893 23489 3896
rect 23523 3893 23535 3927
rect 23477 3887 23535 3893
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 24305 3927 24363 3933
rect 24305 3924 24317 3927
rect 24268 3896 24317 3924
rect 24268 3884 24274 3896
rect 24305 3893 24317 3896
rect 24351 3893 24363 3927
rect 25498 3924 25504 3936
rect 25459 3896 25504 3924
rect 24305 3887 24363 3893
rect 25498 3884 25504 3896
rect 25556 3884 25562 3936
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 51169 3927 51227 3933
rect 51169 3924 51181 3927
rect 51132 3896 51181 3924
rect 51132 3884 51138 3896
rect 51169 3893 51181 3896
rect 51215 3893 51227 3927
rect 51169 3887 51227 3893
rect 51350 3884 51356 3936
rect 51408 3924 51414 3936
rect 51813 3927 51871 3933
rect 51813 3924 51825 3927
rect 51408 3896 51825 3924
rect 51408 3884 51414 3896
rect 51813 3893 51825 3896
rect 51859 3893 51871 3927
rect 51813 3887 51871 3893
rect 52454 3884 52460 3936
rect 52512 3924 52518 3936
rect 54036 3933 54064 3964
rect 53377 3927 53435 3933
rect 53377 3924 53389 3927
rect 52512 3896 53389 3924
rect 52512 3884 52518 3896
rect 53377 3893 53389 3896
rect 53423 3893 53435 3927
rect 53377 3887 53435 3893
rect 54021 3927 54079 3933
rect 54021 3893 54033 3927
rect 54067 3893 54079 3927
rect 55306 3924 55312 3936
rect 55267 3896 55312 3924
rect 54021 3887 54079 3893
rect 55306 3884 55312 3896
rect 55364 3884 55370 3936
rect 58161 3927 58219 3933
rect 58161 3893 58173 3927
rect 58207 3924 58219 3927
rect 58434 3924 58440 3936
rect 58207 3896 58440 3924
rect 58207 3893 58219 3896
rect 58161 3887 58219 3893
rect 58434 3884 58440 3896
rect 58492 3884 58498 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 7006 3720 7012 3732
rect 4856 3692 7012 3720
rect 4856 3680 4862 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8294 3720 8300 3732
rect 7975 3692 8300 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9033 3723 9091 3729
rect 9033 3689 9045 3723
rect 9079 3720 9091 3723
rect 9306 3720 9312 3732
rect 9079 3692 9312 3720
rect 9079 3689 9091 3692
rect 9033 3683 9091 3689
rect 9306 3680 9312 3692
rect 9364 3680 9370 3732
rect 9766 3720 9772 3732
rect 9727 3692 9772 3720
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 12066 3720 12072 3732
rect 10735 3692 12072 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 12066 3680 12072 3692
rect 12124 3680 12130 3732
rect 12897 3723 12955 3729
rect 12897 3689 12909 3723
rect 12943 3720 12955 3723
rect 14642 3720 14648 3732
rect 12943 3692 14648 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 14642 3680 14648 3692
rect 14700 3680 14706 3732
rect 17034 3720 17040 3732
rect 16995 3692 17040 3720
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 18601 3723 18659 3729
rect 18601 3689 18613 3723
rect 18647 3720 18659 3723
rect 18874 3720 18880 3732
rect 18647 3692 18880 3720
rect 18647 3689 18659 3692
rect 18601 3683 18659 3689
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 20257 3723 20315 3729
rect 20257 3689 20269 3723
rect 20303 3720 20315 3723
rect 20438 3720 20444 3732
rect 20303 3692 20444 3720
rect 20303 3689 20315 3692
rect 20257 3683 20315 3689
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 21082 3720 21088 3732
rect 21043 3692 21088 3720
rect 21082 3680 21088 3692
rect 21140 3680 21146 3732
rect 21910 3720 21916 3732
rect 21871 3692 21916 3720
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 32030 3680 32036 3732
rect 32088 3720 32094 3732
rect 32309 3723 32367 3729
rect 32309 3720 32321 3723
rect 32088 3692 32321 3720
rect 32088 3680 32094 3692
rect 32309 3689 32321 3692
rect 32355 3689 32367 3723
rect 32309 3683 32367 3689
rect 52730 3680 52736 3732
rect 52788 3720 52794 3732
rect 52788 3692 55214 3720
rect 52788 3680 52794 3692
rect 2958 3612 2964 3664
rect 3016 3652 3022 3664
rect 3602 3652 3608 3664
rect 3016 3624 3608 3652
rect 3016 3612 3022 3624
rect 3602 3612 3608 3624
rect 3660 3652 3666 3664
rect 3789 3655 3847 3661
rect 3789 3652 3801 3655
rect 3660 3624 3801 3652
rect 3660 3612 3666 3624
rect 3789 3621 3801 3624
rect 3835 3621 3847 3655
rect 3789 3615 3847 3621
rect 6270 3612 6276 3664
rect 6328 3652 6334 3664
rect 6730 3652 6736 3664
rect 6328 3624 6736 3652
rect 6328 3612 6334 3624
rect 6730 3612 6736 3624
rect 6788 3612 6794 3664
rect 7466 3652 7472 3664
rect 7427 3624 7472 3652
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 7837 3655 7895 3661
rect 7837 3621 7849 3655
rect 7883 3652 7895 3655
rect 8478 3652 8484 3664
rect 7883 3624 8484 3652
rect 7883 3621 7895 3624
rect 7837 3615 7895 3621
rect 8478 3612 8484 3624
rect 8536 3612 8542 3664
rect 10873 3655 10931 3661
rect 10873 3652 10885 3655
rect 10152 3624 10885 3652
rect 10152 3596 10180 3624
rect 10873 3621 10885 3624
rect 10919 3621 10931 3655
rect 10873 3615 10931 3621
rect 6178 3584 6184 3596
rect 6139 3556 6184 3584
rect 6178 3544 6184 3556
rect 6236 3544 6242 3596
rect 8018 3584 8024 3596
rect 7979 3556 8024 3584
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8754 3584 8760 3596
rect 8435 3556 8760 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8754 3544 8760 3556
rect 8812 3544 8818 3596
rect 10134 3584 10140 3596
rect 9048 3556 10140 3584
rect 1854 3516 1860 3528
rect 1767 3488 1860 3516
rect 1854 3476 1860 3488
rect 1912 3516 1918 3528
rect 2406 3516 2412 3528
rect 1912 3488 2412 3516
rect 1912 3476 1918 3488
rect 2406 3476 2412 3488
rect 2464 3516 2470 3528
rect 5169 3519 5227 3525
rect 5169 3516 5181 3519
rect 2464 3488 4016 3516
rect 2464 3476 2470 3488
rect 2124 3451 2182 3457
rect 2124 3417 2136 3451
rect 2170 3448 2182 3451
rect 3418 3448 3424 3460
rect 2170 3420 3424 3448
rect 2170 3417 2182 3420
rect 2124 3411 2182 3417
rect 3418 3408 3424 3420
rect 3476 3408 3482 3460
rect 3988 3448 4016 3488
rect 4264 3488 5181 3516
rect 4264 3448 4292 3488
rect 5169 3485 5181 3488
rect 5215 3485 5227 3519
rect 5169 3479 5227 3485
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 6457 3519 6515 3525
rect 6457 3516 6469 3519
rect 5868 3488 6469 3516
rect 5868 3476 5874 3488
rect 6457 3485 6469 3488
rect 6503 3516 6515 3519
rect 9048 3516 9076 3556
rect 10134 3544 10140 3556
rect 10192 3544 10198 3596
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 10686 3584 10692 3596
rect 10468 3556 10692 3584
rect 10468 3544 10474 3556
rect 10686 3544 10692 3556
rect 10744 3584 10750 3596
rect 10781 3587 10839 3593
rect 10781 3584 10793 3587
rect 10744 3556 10793 3584
rect 10744 3544 10750 3556
rect 10781 3553 10793 3556
rect 10827 3553 10839 3587
rect 10888 3584 10916 3615
rect 10962 3612 10968 3664
rect 11020 3652 11026 3664
rect 13541 3655 13599 3661
rect 11020 3624 11065 3652
rect 11020 3612 11026 3624
rect 13541 3621 13553 3655
rect 13587 3652 13599 3655
rect 14185 3655 14243 3661
rect 14185 3652 14197 3655
rect 13587 3624 14197 3652
rect 13587 3621 13599 3624
rect 13541 3615 13599 3621
rect 14185 3621 14197 3624
rect 14231 3621 14243 3655
rect 14185 3615 14243 3621
rect 16209 3655 16267 3661
rect 16209 3621 16221 3655
rect 16255 3652 16267 3655
rect 16390 3652 16396 3664
rect 16255 3624 16396 3652
rect 16255 3621 16267 3624
rect 16209 3615 16267 3621
rect 16390 3612 16396 3624
rect 16448 3612 16454 3664
rect 17862 3652 17868 3664
rect 17823 3624 17868 3652
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 25498 3652 25504 3664
rect 19116 3624 25504 3652
rect 19116 3612 19122 3624
rect 25498 3612 25504 3624
rect 25556 3612 25562 3664
rect 46290 3612 46296 3664
rect 46348 3652 46354 3664
rect 46937 3655 46995 3661
rect 46937 3652 46949 3655
rect 46348 3624 46949 3652
rect 46348 3612 46354 3624
rect 46937 3621 46949 3624
rect 46983 3621 46995 3655
rect 46937 3615 46995 3621
rect 51442 3612 51448 3664
rect 51500 3652 51506 3664
rect 52825 3655 52883 3661
rect 52825 3652 52837 3655
rect 51500 3624 52837 3652
rect 51500 3612 51506 3624
rect 52825 3621 52837 3624
rect 52871 3621 52883 3655
rect 55186 3652 55214 3692
rect 55309 3655 55367 3661
rect 55309 3652 55321 3655
rect 55186 3624 55321 3652
rect 52825 3615 52883 3621
rect 55309 3621 55321 3624
rect 55355 3621 55367 3655
rect 55309 3615 55367 3621
rect 11974 3584 11980 3596
rect 10888 3556 11980 3584
rect 10781 3547 10839 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 12253 3587 12311 3593
rect 12253 3553 12265 3587
rect 12299 3584 12311 3587
rect 14366 3584 14372 3596
rect 12299 3556 14372 3584
rect 12299 3553 12311 3556
rect 12253 3547 12311 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 14734 3584 14740 3596
rect 14695 3556 14740 3584
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 15930 3544 15936 3596
rect 15988 3584 15994 3596
rect 15988 3556 16988 3584
rect 15988 3544 15994 3556
rect 9214 3516 9220 3528
rect 6503 3488 9076 3516
rect 9175 3488 9220 3516
rect 6503 3485 6515 3488
rect 6457 3479 6515 3485
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9640 3488 9965 3516
rect 9640 3476 9646 3488
rect 9953 3485 9965 3488
rect 9999 3516 10011 3519
rect 10318 3516 10324 3528
rect 9999 3488 10324 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 11333 3519 11391 3525
rect 11333 3516 11345 3519
rect 10652 3488 11345 3516
rect 10652 3476 10658 3488
rect 11333 3485 11345 3488
rect 11379 3516 11391 3519
rect 11698 3516 11704 3528
rect 11379 3488 11704 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 13906 3516 13912 3528
rect 13403 3488 13912 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 3988 3420 4292 3448
rect 4924 3451 4982 3457
rect 4924 3417 4936 3451
rect 4970 3448 4982 3451
rect 5074 3448 5080 3460
rect 4970 3420 5080 3448
rect 4970 3417 4982 3420
rect 4924 3411 4982 3417
rect 5074 3408 5080 3420
rect 5132 3408 5138 3460
rect 5721 3451 5779 3457
rect 5721 3417 5733 3451
rect 5767 3448 5779 3451
rect 5767 3420 12434 3448
rect 5767 3417 5779 3420
rect 5721 3411 5779 3417
rect 3237 3383 3295 3389
rect 3237 3349 3249 3383
rect 3283 3380 3295 3383
rect 3326 3380 3332 3392
rect 3283 3352 3332 3380
rect 3283 3349 3295 3352
rect 3237 3343 3295 3349
rect 3326 3340 3332 3352
rect 3384 3340 3390 3392
rect 3510 3340 3516 3392
rect 3568 3380 3574 3392
rect 8478 3380 8484 3392
rect 3568 3352 8484 3380
rect 3568 3340 3574 3352
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 9398 3380 9404 3392
rect 8628 3352 9404 3380
rect 8628 3340 8634 3352
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 12406 3380 12434 3420
rect 13372 3380 13400 3479
rect 13906 3476 13912 3488
rect 13964 3476 13970 3528
rect 13998 3476 14004 3528
rect 14056 3516 14062 3528
rect 14645 3519 14703 3525
rect 14645 3516 14657 3519
rect 14056 3488 14657 3516
rect 14056 3476 14062 3488
rect 14645 3485 14657 3488
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15746 3516 15752 3528
rect 14976 3488 15752 3516
rect 14976 3476 14982 3488
rect 15746 3476 15752 3488
rect 15804 3516 15810 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15804 3488 16037 3516
rect 15804 3476 15810 3488
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 16850 3516 16856 3528
rect 16811 3488 16856 3516
rect 16025 3479 16083 3485
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 16960 3516 16988 3556
rect 17402 3544 17408 3596
rect 17460 3584 17466 3596
rect 18690 3584 18696 3596
rect 17460 3556 18696 3584
rect 17460 3544 17466 3556
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 19613 3587 19671 3593
rect 19613 3553 19625 3587
rect 19659 3584 19671 3587
rect 21450 3584 21456 3596
rect 19659 3556 21456 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 30926 3584 30932 3596
rect 30887 3556 30932 3584
rect 30926 3544 30932 3556
rect 30984 3544 30990 3596
rect 50798 3544 50804 3596
rect 50856 3584 50862 3596
rect 51537 3587 51595 3593
rect 51537 3584 51549 3587
rect 50856 3556 51549 3584
rect 50856 3544 50862 3556
rect 51537 3553 51549 3556
rect 51583 3553 51595 3587
rect 51537 3547 51595 3553
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 53469 3587 53527 3593
rect 53469 3584 53481 3587
rect 51684 3556 53481 3584
rect 51684 3544 51690 3556
rect 53469 3553 53481 3556
rect 53515 3553 53527 3587
rect 53469 3547 53527 3553
rect 53834 3544 53840 3596
rect 53892 3584 53898 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 53892 3556 56609 3584
rect 53892 3544 53898 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 17494 3516 17500 3528
rect 16960 3488 17500 3516
rect 17494 3476 17500 3488
rect 17552 3516 17558 3528
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17552 3488 17693 3516
rect 17552 3476 17558 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18417 3519 18475 3525
rect 18417 3516 18429 3519
rect 18380 3488 18429 3516
rect 18380 3476 18386 3488
rect 18417 3485 18429 3488
rect 18463 3485 18475 3519
rect 18417 3479 18475 3485
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 19576 3488 20085 3516
rect 19576 3476 19582 3488
rect 20073 3485 20085 3488
rect 20119 3485 20131 3519
rect 20073 3479 20131 3485
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 20901 3519 20959 3525
rect 20901 3516 20913 3519
rect 20864 3488 20913 3516
rect 20864 3476 20870 3488
rect 20901 3485 20913 3488
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 21634 3476 21640 3528
rect 21692 3516 21698 3528
rect 21729 3519 21787 3525
rect 21729 3516 21741 3519
rect 21692 3488 21741 3516
rect 21692 3476 21698 3488
rect 21729 3485 21741 3488
rect 21775 3485 21787 3519
rect 21729 3479 21787 3485
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 23658 3516 23664 3528
rect 23247 3488 23664 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 23934 3516 23940 3528
rect 23891 3488 23940 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 23934 3476 23940 3488
rect 23992 3476 23998 3528
rect 24762 3476 24768 3528
rect 24820 3516 24826 3528
rect 24857 3519 24915 3525
rect 24857 3516 24869 3519
rect 24820 3488 24869 3516
rect 24820 3476 24826 3488
rect 24857 3485 24869 3488
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 25590 3476 25596 3528
rect 25648 3516 25654 3528
rect 25685 3519 25743 3525
rect 25685 3516 25697 3519
rect 25648 3488 25697 3516
rect 25648 3476 25654 3488
rect 25685 3485 25697 3488
rect 25731 3485 25743 3519
rect 25685 3479 25743 3485
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 26789 3519 26847 3525
rect 26789 3516 26801 3519
rect 26752 3488 26801 3516
rect 26752 3476 26758 3488
rect 26789 3485 26801 3488
rect 26835 3485 26847 3519
rect 26789 3479 26847 3485
rect 27522 3476 27528 3528
rect 27580 3516 27586 3528
rect 27617 3519 27675 3525
rect 27617 3516 27629 3519
rect 27580 3488 27629 3516
rect 27580 3476 27586 3488
rect 27617 3485 27629 3488
rect 27663 3485 27675 3519
rect 27617 3479 27675 3485
rect 28626 3476 28632 3528
rect 28684 3516 28690 3528
rect 28721 3519 28779 3525
rect 28721 3516 28733 3519
rect 28684 3488 28733 3516
rect 28684 3476 28690 3488
rect 28721 3485 28733 3488
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 30834 3476 30840 3528
rect 30892 3516 30898 3528
rect 31185 3519 31243 3525
rect 31185 3516 31197 3519
rect 30892 3488 31197 3516
rect 30892 3476 30898 3488
rect 31185 3485 31197 3488
rect 31231 3485 31243 3519
rect 31185 3479 31243 3485
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34793 3519 34851 3525
rect 34793 3516 34805 3519
rect 34756 3488 34805 3516
rect 34756 3476 34762 3488
rect 34793 3485 34805 3488
rect 34839 3485 34851 3519
rect 34793 3479 34851 3485
rect 35342 3476 35348 3528
rect 35400 3516 35406 3528
rect 35437 3519 35495 3525
rect 35437 3516 35449 3519
rect 35400 3488 35449 3516
rect 35400 3476 35406 3488
rect 35437 3485 35449 3488
rect 35483 3485 35495 3519
rect 35437 3479 35495 3485
rect 35802 3476 35808 3528
rect 35860 3516 35866 3528
rect 36081 3519 36139 3525
rect 36081 3516 36093 3519
rect 35860 3488 36093 3516
rect 35860 3476 35866 3488
rect 36081 3485 36093 3488
rect 36127 3485 36139 3519
rect 36081 3479 36139 3485
rect 36630 3476 36636 3528
rect 36688 3516 36694 3528
rect 36725 3519 36783 3525
rect 36725 3516 36737 3519
rect 36688 3488 36737 3516
rect 36688 3476 36694 3488
rect 36725 3485 36737 3488
rect 36771 3485 36783 3519
rect 36725 3479 36783 3485
rect 37458 3476 37464 3528
rect 37516 3516 37522 3528
rect 37553 3519 37611 3525
rect 37553 3516 37565 3519
rect 37516 3488 37565 3516
rect 37516 3476 37522 3488
rect 37553 3485 37565 3488
rect 37599 3485 37611 3519
rect 37553 3479 37611 3485
rect 38562 3476 38568 3528
rect 38620 3516 38626 3528
rect 38657 3519 38715 3525
rect 38657 3516 38669 3519
rect 38620 3488 38669 3516
rect 38620 3476 38626 3488
rect 38657 3485 38669 3488
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 40000 3488 40049 3516
rect 40000 3476 40006 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40494 3476 40500 3528
rect 40552 3516 40558 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40552 3488 40693 3516
rect 40552 3476 40558 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 40681 3479 40739 3485
rect 41046 3476 41052 3528
rect 41104 3516 41110 3528
rect 41325 3519 41383 3525
rect 41325 3516 41337 3519
rect 41104 3488 41337 3516
rect 41104 3476 41110 3488
rect 41325 3485 41337 3488
rect 41371 3485 41383 3519
rect 41325 3479 41383 3485
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 42521 3519 42579 3525
rect 42521 3516 42533 3519
rect 42484 3488 42533 3516
rect 42484 3476 42490 3488
rect 42521 3485 42533 3488
rect 42567 3485 42579 3519
rect 42521 3479 42579 3485
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 43165 3519 43223 3525
rect 43165 3516 43177 3519
rect 42760 3488 43177 3516
rect 42760 3476 42766 3488
rect 43165 3485 43177 3488
rect 43211 3485 43223 3519
rect 43165 3479 43223 3485
rect 44358 3476 44364 3528
rect 44416 3516 44422 3528
rect 45005 3519 45063 3525
rect 45005 3516 45017 3519
rect 44416 3488 45017 3516
rect 44416 3476 44422 3488
rect 45005 3485 45017 3488
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 45186 3476 45192 3528
rect 45244 3516 45250 3528
rect 45649 3519 45707 3525
rect 45649 3516 45661 3519
rect 45244 3488 45661 3516
rect 45244 3476 45250 3488
rect 45649 3485 45661 3488
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 46014 3476 46020 3528
rect 46072 3516 46078 3528
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 46072 3488 46305 3516
rect 46072 3476 46078 3488
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 47670 3476 47676 3528
rect 47728 3516 47734 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47728 3488 47777 3516
rect 47728 3476 47734 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 48222 3476 48228 3528
rect 48280 3516 48286 3528
rect 48409 3519 48467 3525
rect 48409 3516 48421 3519
rect 48280 3488 48421 3516
rect 48280 3476 48286 3488
rect 48409 3485 48421 3488
rect 48455 3485 48467 3519
rect 48409 3479 48467 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50249 3519 50307 3525
rect 50249 3516 50261 3519
rect 50212 3488 50261 3516
rect 50212 3476 50218 3488
rect 50249 3485 50261 3488
rect 50295 3485 50307 3519
rect 50249 3479 50307 3485
rect 50614 3476 50620 3528
rect 50672 3516 50678 3528
rect 50893 3519 50951 3525
rect 50893 3516 50905 3519
rect 50672 3488 50905 3516
rect 50672 3476 50678 3488
rect 50893 3485 50905 3488
rect 50939 3485 50951 3519
rect 50893 3479 50951 3485
rect 51166 3476 51172 3528
rect 51224 3516 51230 3528
rect 52181 3519 52239 3525
rect 52181 3516 52193 3519
rect 51224 3488 52193 3516
rect 51224 3476 51230 3488
rect 52181 3485 52193 3488
rect 52227 3485 52239 3519
rect 52181 3479 52239 3485
rect 52270 3476 52276 3528
rect 52328 3516 52334 3528
rect 54113 3519 54171 3525
rect 54113 3516 54125 3519
rect 52328 3488 54125 3516
rect 52328 3476 52334 3488
rect 54113 3485 54125 3488
rect 54159 3485 54171 3519
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 54113 3479 54171 3485
rect 55186 3488 55965 3516
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 14185 3451 14243 3457
rect 14185 3448 14197 3451
rect 13596 3420 14197 3448
rect 13596 3408 13602 3420
rect 14185 3417 14197 3420
rect 14231 3417 14243 3451
rect 14185 3411 14243 3417
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 15286 3448 15292 3460
rect 14884 3420 15292 3448
rect 14884 3408 14890 3420
rect 15286 3408 15292 3420
rect 15344 3408 15350 3460
rect 17770 3408 17776 3460
rect 17828 3448 17834 3460
rect 23474 3448 23480 3460
rect 17828 3420 23480 3448
rect 17828 3408 17834 3420
rect 23474 3408 23480 3420
rect 23532 3408 23538 3460
rect 53282 3408 53288 3460
rect 53340 3448 53346 3460
rect 55186 3448 55214 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 57514 3516 57520 3528
rect 57475 3488 57520 3516
rect 55953 3479 56011 3485
rect 57514 3476 57520 3488
rect 57572 3476 57578 3528
rect 58158 3516 58164 3528
rect 58119 3488 58164 3516
rect 58158 3476 58164 3488
rect 58216 3476 58222 3528
rect 53340 3420 55214 3448
rect 53340 3408 53346 3420
rect 14918 3380 14924 3392
rect 12406 3352 13400 3380
rect 14879 3352 14924 3380
rect 14918 3340 14924 3352
rect 14976 3340 14982 3392
rect 15473 3383 15531 3389
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 19518 3380 19524 3392
rect 15519 3352 19524 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 19518 3340 19524 3352
rect 19576 3340 19582 3392
rect 22557 3383 22615 3389
rect 22557 3349 22569 3383
rect 22603 3380 22615 3383
rect 22830 3380 22836 3392
rect 22603 3352 22836 3380
rect 22603 3349 22615 3352
rect 22557 3343 22615 3349
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 3786 3176 3792 3188
rect 3747 3148 3792 3176
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5655 3179 5713 3185
rect 4764 3148 5580 3176
rect 4764 3136 4770 3148
rect 1946 3108 1952 3120
rect 1907 3080 1952 3108
rect 1946 3068 1952 3080
rect 2004 3068 2010 3120
rect 2676 3111 2734 3117
rect 2676 3077 2688 3111
rect 2722 3108 2734 3111
rect 2774 3108 2780 3120
rect 2722 3080 2780 3108
rect 2722 3077 2734 3080
rect 2676 3071 2734 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 3234 3068 3240 3120
rect 3292 3108 3298 3120
rect 5445 3111 5503 3117
rect 5445 3108 5457 3111
rect 3292 3080 5457 3108
rect 3292 3068 3298 3080
rect 5445 3077 5457 3080
rect 5491 3077 5503 3111
rect 5552 3108 5580 3148
rect 5655 3145 5667 3179
rect 5701 3176 5713 3179
rect 6822 3176 6828 3188
rect 5701 3148 6828 3176
rect 5701 3145 5713 3148
rect 5655 3139 5713 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 8018 3176 8024 3188
rect 6972 3148 8024 3176
rect 6972 3136 6978 3148
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8570 3176 8576 3188
rect 8343 3148 8576 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8570 3136 8576 3148
rect 8628 3136 8634 3188
rect 8846 3136 8852 3188
rect 8904 3176 8910 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 8904 3148 11621 3176
rect 8904 3136 8910 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 14458 3176 14464 3188
rect 14419 3148 14464 3176
rect 11609 3139 11667 3145
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 14936 3148 16620 3176
rect 5552 3080 6868 3108
rect 5445 3071 5503 3077
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1544 3012 1777 3040
rect 1544 3000 1550 3012
rect 1765 3009 1777 3012
rect 1811 3009 1823 3043
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 1765 3003 1823 3009
rect 1780 2972 1808 3003
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 4798 3040 4804 3052
rect 2516 3012 4804 3040
rect 2516 2972 2544 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5258 3040 5264 3052
rect 5031 3012 5264 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6840 3049 6868 3080
rect 7374 3068 7380 3120
rect 7432 3108 7438 3120
rect 13722 3108 13728 3120
rect 7432 3080 13728 3108
rect 7432 3068 7438 3080
rect 13722 3068 13728 3080
rect 13780 3068 13786 3120
rect 14936 3108 14964 3148
rect 15102 3108 15108 3120
rect 13924 3080 14964 3108
rect 15063 3080 15108 3108
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6512 3012 6561 3040
rect 6512 3000 6518 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 1780 2944 2544 2972
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 6086 2972 6092 2984
rect 3752 2944 6092 2972
rect 3752 2932 3758 2944
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 6840 2972 6868 3003
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7616 3012 8033 3040
rect 7616 3000 7622 3012
rect 8021 3009 8033 3012
rect 8067 3040 8079 3043
rect 8202 3040 8208 3052
rect 8067 3012 8208 3040
rect 8067 3009 8079 3012
rect 8021 3003 8079 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8754 3040 8760 3052
rect 8536 3012 8760 3040
rect 8536 3000 8542 3012
rect 8754 3000 8760 3012
rect 8812 3040 8818 3052
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8812 3012 8953 3040
rect 8812 3000 8818 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 8941 3003 8999 3009
rect 9048 3012 9873 3040
rect 9048 2972 9076 3012
rect 9861 3009 9873 3012
rect 9907 3009 9919 3043
rect 10686 3040 10692 3052
rect 10647 3012 10692 3040
rect 9861 3003 9919 3009
rect 10686 3000 10692 3012
rect 10744 3000 10750 3052
rect 11790 3040 11796 3052
rect 11751 3012 11796 3040
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 13924 3049 13952 3080
rect 15102 3068 15108 3080
rect 15160 3068 15166 3120
rect 16117 3111 16175 3117
rect 16117 3077 16129 3111
rect 16163 3108 16175 3111
rect 16298 3108 16304 3120
rect 16163 3080 16304 3108
rect 16163 3077 16175 3080
rect 16117 3071 16175 3077
rect 16298 3068 16304 3080
rect 16356 3068 16362 3120
rect 16592 3108 16620 3148
rect 16666 3136 16672 3188
rect 16724 3176 16730 3188
rect 17034 3176 17040 3188
rect 16724 3148 17040 3176
rect 16724 3136 16730 3148
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 18230 3176 18236 3188
rect 18191 3148 18236 3176
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18874 3176 18880 3188
rect 18835 3148 18880 3176
rect 18874 3136 18880 3148
rect 18932 3136 18938 3188
rect 20346 3176 20352 3188
rect 20307 3148 20352 3176
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 21082 3176 21088 3188
rect 21043 3148 21088 3176
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 21266 3136 21272 3188
rect 21324 3176 21330 3188
rect 22646 3176 22652 3188
rect 21324 3148 22652 3176
rect 21324 3136 21330 3148
rect 22646 3136 22652 3148
rect 22704 3136 22710 3188
rect 23014 3176 23020 3188
rect 22975 3148 23020 3176
rect 23014 3136 23020 3148
rect 23072 3136 23078 3188
rect 17310 3108 17316 3120
rect 16592 3080 17316 3108
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 17586 3108 17592 3120
rect 17547 3080 17592 3108
rect 17586 3068 17592 3080
rect 17644 3068 17650 3120
rect 18892 3080 20116 3108
rect 18892 3052 18920 3080
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 14826 3040 14832 3052
rect 14599 3012 14832 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 15010 3000 15016 3052
rect 15068 3040 15074 3052
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 15068 3012 15301 3040
rect 15068 3000 15074 3012
rect 15289 3009 15301 3012
rect 15335 3040 15347 3043
rect 15562 3040 15568 3052
rect 15335 3012 15568 3040
rect 15335 3009 15347 3012
rect 15289 3003 15347 3009
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3040 15991 3043
rect 16574 3040 16580 3052
rect 15979 3012 16580 3040
rect 15979 3009 15991 3012
rect 15933 3003 15991 3009
rect 16574 3000 16580 3012
rect 16632 3000 16638 3052
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3040 17463 3043
rect 17770 3040 17776 3052
rect 17451 3012 17776 3040
rect 17451 3009 17463 3012
rect 17405 3003 17463 3009
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 18012 3012 18061 3040
rect 18012 3000 18018 3012
rect 18049 3009 18061 3012
rect 18095 3040 18107 3043
rect 18598 3040 18604 3052
rect 18095 3012 18604 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18874 3000 18880 3052
rect 18932 3000 18938 3052
rect 19058 3040 19064 3052
rect 19019 3012 19064 3040
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19797 3043 19855 3049
rect 19797 3009 19809 3043
rect 19843 3040 19855 3043
rect 19978 3040 19984 3052
rect 19843 3012 19984 3040
rect 19843 3009 19855 3012
rect 19797 3003 19855 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 20088 3040 20116 3080
rect 20254 3068 20260 3120
rect 20312 3108 20318 3120
rect 20441 3111 20499 3117
rect 20441 3108 20453 3111
rect 20312 3080 20453 3108
rect 20312 3068 20318 3080
rect 20441 3077 20453 3080
rect 20487 3108 20499 3111
rect 20530 3108 20536 3120
rect 20487 3080 20536 3108
rect 20487 3077 20499 3080
rect 20441 3071 20499 3077
rect 20530 3068 20536 3080
rect 20588 3068 20594 3120
rect 22186 3108 22192 3120
rect 21376 3080 22192 3108
rect 21376 3052 21404 3080
rect 22186 3068 22192 3080
rect 22244 3068 22250 3120
rect 51902 3068 51908 3120
rect 51960 3108 51966 3120
rect 51960 3080 54708 3108
rect 51960 3068 51966 3080
rect 21269 3043 21327 3049
rect 20088 3012 21128 3040
rect 10410 2972 10416 2984
rect 6840 2944 7972 2972
rect 5350 2904 5356 2916
rect 4080 2876 5356 2904
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 4080 2836 4108 2876
rect 5350 2864 5356 2876
rect 5408 2864 5414 2916
rect 7742 2904 7748 2916
rect 5460 2876 7748 2904
rect 2648 2808 4108 2836
rect 4801 2839 4859 2845
rect 2648 2796 2654 2808
rect 4801 2805 4813 2839
rect 4847 2836 4859 2839
rect 5460 2836 5488 2876
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 5626 2836 5632 2848
rect 4847 2808 5488 2836
rect 5587 2808 5632 2836
rect 4847 2805 4859 2808
rect 4801 2799 4859 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 5813 2839 5871 2845
rect 5813 2805 5825 2839
rect 5859 2836 5871 2839
rect 6546 2836 6552 2848
rect 5859 2808 6552 2836
rect 5859 2805 5871 2808
rect 5813 2799 5871 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 7944 2836 7972 2944
rect 8036 2944 9076 2972
rect 9140 2944 10416 2972
rect 8036 2916 8064 2944
rect 8018 2864 8024 2916
rect 8076 2864 8082 2916
rect 9140 2836 9168 2944
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 13265 2975 13323 2981
rect 13265 2941 13277 2975
rect 13311 2972 13323 2975
rect 15654 2972 15660 2984
rect 13311 2944 15660 2972
rect 13311 2941 13323 2944
rect 13265 2935 13323 2941
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 21100 2972 21128 3012
rect 21269 3009 21281 3043
rect 21315 3040 21327 3043
rect 21358 3040 21364 3052
rect 21315 3012 21364 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 21358 3000 21364 3012
rect 21416 3000 21422 3052
rect 22094 3000 22100 3052
rect 22152 3040 22158 3052
rect 22830 3040 22836 3052
rect 22152 3012 22197 3040
rect 22791 3012 22836 3040
rect 22152 3000 22158 3012
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 34514 3040 34520 3052
rect 31726 3012 34520 3040
rect 23198 2972 23204 2984
rect 21100 2944 23204 2972
rect 23198 2932 23204 2944
rect 23256 2932 23262 2984
rect 23845 2975 23903 2981
rect 23845 2941 23857 2975
rect 23891 2972 23903 2975
rect 24486 2972 24492 2984
rect 23891 2944 24492 2972
rect 23891 2941 23903 2944
rect 23845 2935 23903 2941
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 9398 2864 9404 2916
rect 9456 2904 9462 2916
rect 10873 2907 10931 2913
rect 10873 2904 10885 2907
rect 9456 2876 10885 2904
rect 9456 2864 9462 2876
rect 10873 2873 10885 2876
rect 10919 2873 10931 2907
rect 10873 2867 10931 2873
rect 12621 2907 12679 2913
rect 12621 2873 12633 2907
rect 12667 2904 12679 2907
rect 14918 2904 14924 2916
rect 12667 2876 14924 2904
rect 12667 2873 12679 2876
rect 12621 2867 12679 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 17862 2904 17868 2916
rect 15028 2876 17868 2904
rect 7944 2808 9168 2836
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9490 2836 9496 2848
rect 9263 2808 9496 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 9953 2839 10011 2845
rect 9953 2836 9965 2839
rect 9732 2808 9965 2836
rect 9732 2796 9738 2808
rect 9953 2805 9965 2808
rect 9999 2805 10011 2839
rect 9953 2799 10011 2805
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 15028 2836 15056 2876
rect 17862 2864 17868 2876
rect 17920 2864 17926 2916
rect 17954 2864 17960 2916
rect 18012 2904 18018 2916
rect 18874 2904 18880 2916
rect 18012 2876 18880 2904
rect 18012 2864 18018 2876
rect 18874 2864 18880 2876
rect 18932 2864 18938 2916
rect 19613 2907 19671 2913
rect 19613 2873 19625 2907
rect 19659 2904 19671 2907
rect 31726 2904 31754 3012
rect 34514 3000 34520 3012
rect 34572 3000 34578 3052
rect 51718 3000 51724 3052
rect 51776 3040 51782 3052
rect 54680 3049 54708 3080
rect 54021 3043 54079 3049
rect 54021 3040 54033 3043
rect 51776 3012 54033 3040
rect 51776 3000 51782 3012
rect 54021 3009 54033 3012
rect 54067 3009 54079 3043
rect 54021 3003 54079 3009
rect 54665 3043 54723 3049
rect 54665 3009 54677 3043
rect 54711 3009 54723 3043
rect 54665 3003 54723 3009
rect 54754 3000 54760 3052
rect 54812 3040 54818 3052
rect 55309 3043 55367 3049
rect 55309 3040 55321 3043
rect 54812 3012 55321 3040
rect 54812 3000 54818 3012
rect 55309 3009 55321 3012
rect 55355 3009 55367 3043
rect 55309 3003 55367 3009
rect 32766 2932 32772 2984
rect 32824 2972 32830 2984
rect 33413 2975 33471 2981
rect 33413 2972 33425 2975
rect 32824 2944 33425 2972
rect 32824 2932 32830 2944
rect 33413 2941 33425 2944
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 38286 2932 38292 2984
rect 38344 2972 38350 2984
rect 39209 2975 39267 2981
rect 39209 2972 39221 2975
rect 38344 2944 39221 2972
rect 38344 2932 38350 2944
rect 39209 2941 39221 2944
rect 39255 2941 39267 2975
rect 39209 2935 39267 2941
rect 42150 2932 42156 2984
rect 42208 2972 42214 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 42208 2944 43085 2972
rect 42208 2932 42214 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 53098 2932 53104 2984
rect 53156 2972 53162 2984
rect 55953 2975 56011 2981
rect 55953 2972 55965 2975
rect 53156 2944 55965 2972
rect 53156 2932 53162 2944
rect 55953 2941 55965 2944
rect 55999 2941 56011 2975
rect 56594 2972 56600 2984
rect 56555 2944 56600 2972
rect 55953 2935 56011 2941
rect 56594 2932 56600 2944
rect 56652 2932 56658 2984
rect 19659 2876 31754 2904
rect 19659 2873 19671 2876
rect 19613 2867 19671 2873
rect 33870 2864 33876 2916
rect 33928 2904 33934 2916
rect 34701 2907 34759 2913
rect 34701 2904 34713 2907
rect 33928 2876 34713 2904
rect 33928 2864 33934 2876
rect 34701 2873 34713 2876
rect 34747 2873 34759 2907
rect 34701 2867 34759 2873
rect 37182 2864 37188 2916
rect 37240 2904 37246 2916
rect 37921 2907 37979 2913
rect 37921 2904 37933 2907
rect 37240 2876 37933 2904
rect 37240 2864 37246 2876
rect 37921 2873 37933 2876
rect 37967 2873 37979 2907
rect 37921 2867 37979 2873
rect 39114 2864 39120 2916
rect 39172 2904 39178 2916
rect 39853 2907 39911 2913
rect 39853 2904 39865 2907
rect 39172 2876 39865 2904
rect 39172 2864 39178 2876
rect 39853 2873 39865 2876
rect 39899 2873 39911 2907
rect 39853 2867 39911 2873
rect 40218 2864 40224 2916
rect 40276 2904 40282 2916
rect 41141 2907 41199 2913
rect 41141 2904 41153 2907
rect 40276 2876 41153 2904
rect 40276 2864 40282 2876
rect 41141 2873 41153 2876
rect 41187 2873 41199 2907
rect 41141 2867 41199 2873
rect 42978 2864 42984 2916
rect 43036 2904 43042 2916
rect 43717 2907 43775 2913
rect 43717 2904 43729 2907
rect 43036 2876 43729 2904
rect 43036 2864 43042 2876
rect 43717 2873 43729 2876
rect 43763 2873 43775 2907
rect 43717 2867 43775 2873
rect 44082 2864 44088 2916
rect 44140 2904 44146 2916
rect 45005 2907 45063 2913
rect 45005 2904 45017 2907
rect 44140 2876 45017 2904
rect 44140 2864 44146 2876
rect 45005 2873 45017 2876
rect 45051 2873 45063 2907
rect 45649 2907 45707 2913
rect 45649 2904 45661 2907
rect 45005 2867 45063 2873
rect 45112 2876 45661 2904
rect 14792 2808 15056 2836
rect 16853 2839 16911 2845
rect 14792 2796 14798 2808
rect 16853 2805 16865 2839
rect 16899 2836 16911 2839
rect 19426 2836 19432 2848
rect 16899 2808 19432 2836
rect 16899 2805 16911 2808
rect 16853 2799 16911 2805
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 22281 2839 22339 2845
rect 22281 2805 22293 2839
rect 22327 2836 22339 2839
rect 22370 2836 22376 2848
rect 22327 2808 22376 2836
rect 22327 2805 22339 2808
rect 22281 2799 22339 2805
rect 22370 2796 22376 2808
rect 22428 2796 22434 2848
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 25038 2836 25044 2848
rect 24535 2808 25044 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2836 25191 2839
rect 25314 2836 25320 2848
rect 25179 2808 25320 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 25314 2796 25320 2808
rect 25372 2796 25378 2848
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 26142 2836 26148 2848
rect 25823 2808 26148 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 26142 2796 26148 2808
rect 26200 2796 26206 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 26878 2836 26884 2848
rect 26467 2808 26884 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 26878 2796 26884 2808
rect 26936 2796 26942 2848
rect 27617 2839 27675 2845
rect 27617 2805 27629 2839
rect 27663 2836 27675 2839
rect 27798 2836 27804 2848
rect 27663 2808 27804 2836
rect 27663 2805 27675 2808
rect 27617 2799 27675 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28074 2836 28080 2848
rect 28035 2808 28080 2836
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 28905 2839 28963 2845
rect 28905 2805 28917 2839
rect 28951 2836 28963 2839
rect 29178 2836 29184 2848
rect 28951 2808 29184 2836
rect 28951 2805 28963 2808
rect 28905 2799 28963 2805
rect 29178 2796 29184 2808
rect 29236 2796 29242 2848
rect 29549 2839 29607 2845
rect 29549 2805 29561 2839
rect 29595 2836 29607 2839
rect 29730 2836 29736 2848
rect 29595 2808 29736 2836
rect 29595 2805 29607 2808
rect 29549 2799 29607 2805
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 30006 2836 30012 2848
rect 29967 2808 30012 2836
rect 30006 2796 30012 2808
rect 30064 2796 30070 2848
rect 30558 2796 30564 2848
rect 30616 2836 30622 2848
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 30616 2808 30665 2836
rect 30616 2796 30622 2808
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 31662 2796 31668 2848
rect 31720 2836 31726 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31720 2808 32137 2836
rect 31720 2796 31726 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 32769 2839 32827 2845
rect 32769 2836 32781 2839
rect 32272 2808 32781 2836
rect 32272 2796 32278 2808
rect 32769 2805 32781 2808
rect 32815 2805 32827 2839
rect 32769 2799 32827 2805
rect 33318 2796 33324 2848
rect 33376 2836 33382 2848
rect 34057 2839 34115 2845
rect 34057 2836 34069 2839
rect 33376 2808 34069 2836
rect 33376 2796 33382 2808
rect 34057 2805 34069 2808
rect 34103 2805 34115 2839
rect 34057 2799 34115 2805
rect 34422 2796 34428 2848
rect 34480 2836 34486 2848
rect 35345 2839 35403 2845
rect 35345 2836 35357 2839
rect 34480 2808 35357 2836
rect 34480 2796 34486 2808
rect 35345 2805 35357 2808
rect 35391 2805 35403 2839
rect 35345 2799 35403 2805
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35989 2839 36047 2845
rect 35989 2836 36001 2839
rect 35492 2808 36001 2836
rect 35492 2796 35498 2808
rect 35989 2805 36001 2808
rect 36035 2805 36047 2839
rect 35989 2799 36047 2805
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36412 2808 37289 2836
rect 36412 2796 36418 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37734 2796 37740 2848
rect 37792 2836 37798 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 37792 2808 38577 2836
rect 37792 2796 37798 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 39666 2796 39672 2848
rect 39724 2836 39730 2848
rect 40497 2839 40555 2845
rect 40497 2836 40509 2839
rect 39724 2808 40509 2836
rect 39724 2796 39730 2808
rect 40497 2805 40509 2808
rect 40543 2805 40555 2839
rect 40497 2799 40555 2805
rect 41598 2796 41604 2848
rect 41656 2836 41662 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41656 2808 42441 2836
rect 41656 2796 41662 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 43530 2796 43536 2848
rect 43588 2836 43594 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 43588 2808 44373 2836
rect 43588 2796 43594 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 44910 2796 44916 2848
rect 44968 2836 44974 2848
rect 45112 2836 45140 2876
rect 45649 2873 45661 2876
rect 45695 2873 45707 2907
rect 45649 2867 45707 2873
rect 47394 2864 47400 2916
rect 47452 2904 47458 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 47452 2876 48237 2904
rect 47452 2864 47458 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 48774 2864 48780 2916
rect 48832 2904 48838 2916
rect 49513 2907 49571 2913
rect 49513 2904 49525 2907
rect 48832 2876 49525 2904
rect 48832 2864 48838 2876
rect 49513 2873 49525 2876
rect 49559 2873 49571 2907
rect 49513 2867 49571 2873
rect 49878 2864 49884 2916
rect 49936 2904 49942 2916
rect 50801 2907 50859 2913
rect 50801 2904 50813 2907
rect 49936 2876 50813 2904
rect 49936 2864 49942 2876
rect 50801 2873 50813 2876
rect 50847 2873 50859 2907
rect 50801 2867 50859 2873
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 52733 2907 52791 2913
rect 52733 2904 52745 2907
rect 51040 2876 52745 2904
rect 51040 2864 51046 2876
rect 52733 2873 52745 2876
rect 52779 2873 52791 2907
rect 52733 2867 52791 2873
rect 54202 2864 54208 2916
rect 54260 2904 54266 2916
rect 57885 2907 57943 2913
rect 57885 2904 57897 2907
rect 54260 2876 57897 2904
rect 54260 2864 54266 2876
rect 57885 2873 57897 2876
rect 57931 2873 57943 2907
rect 57885 2867 57943 2873
rect 44968 2808 45140 2836
rect 44968 2796 44974 2808
rect 45462 2796 45468 2848
rect 45520 2836 45526 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45520 2808 46305 2836
rect 45520 2796 45526 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 46842 2796 46848 2848
rect 46900 2836 46906 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46900 2808 47593 2836
rect 46900 2796 46906 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 47946 2796 47952 2848
rect 48004 2836 48010 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48004 2808 48881 2836
rect 48004 2796 48010 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49326 2796 49332 2848
rect 49384 2836 49390 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49384 2808 50169 2836
rect 49384 2796 49390 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 50706 2796 50712 2848
rect 50764 2836 50770 2848
rect 51445 2839 51503 2845
rect 51445 2836 51457 2839
rect 50764 2808 51457 2836
rect 50764 2796 50770 2808
rect 51445 2805 51457 2808
rect 51491 2805 51503 2839
rect 51445 2799 51503 2805
rect 51534 2796 51540 2848
rect 51592 2836 51598 2848
rect 53377 2839 53435 2845
rect 53377 2836 53389 2839
rect 51592 2808 53389 2836
rect 51592 2796 51598 2808
rect 53377 2805 53389 2808
rect 53423 2805 53435 2839
rect 53377 2799 53435 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 6270 2632 6276 2644
rect 1627 2604 6276 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 8628 2604 12357 2632
rect 8628 2592 8634 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 12345 2595 12403 2601
rect 13541 2635 13599 2641
rect 13541 2601 13553 2635
rect 13587 2632 13599 2635
rect 14734 2632 14740 2644
rect 13587 2604 14740 2632
rect 13587 2601 13599 2604
rect 13541 2595 13599 2601
rect 14734 2592 14740 2604
rect 14792 2592 14798 2644
rect 15838 2632 15844 2644
rect 14844 2604 15844 2632
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 2682 2564 2688 2576
rect 2455 2536 2688 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 2682 2524 2688 2536
rect 2740 2524 2746 2576
rect 3145 2567 3203 2573
rect 3145 2533 3157 2567
rect 3191 2564 3203 2567
rect 7374 2564 7380 2576
rect 3191 2536 7380 2564
rect 3191 2533 3203 2536
rect 3145 2527 3203 2533
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 9674 2524 9680 2576
rect 9732 2564 9738 2576
rect 11701 2567 11759 2573
rect 11701 2564 11713 2567
rect 9732 2536 11713 2564
rect 9732 2524 9738 2536
rect 11701 2533 11713 2536
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 14369 2567 14427 2573
rect 14369 2533 14381 2567
rect 14415 2564 14427 2567
rect 14550 2564 14556 2576
rect 14415 2536 14556 2564
rect 14415 2533 14427 2536
rect 14369 2527 14427 2533
rect 14550 2524 14556 2536
rect 14608 2524 14614 2576
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7650 2496 7656 2508
rect 7239 2468 7656 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 12618 2496 12624 2508
rect 8435 2468 12624 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 14844 2496 14872 2604
rect 15838 2592 15844 2604
rect 15896 2632 15902 2644
rect 16114 2632 16120 2644
rect 15896 2604 16120 2632
rect 15896 2592 15902 2604
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 17126 2632 17132 2644
rect 17087 2604 17132 2632
rect 17126 2592 17132 2604
rect 17184 2592 17190 2644
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 17773 2635 17831 2641
rect 17773 2632 17785 2635
rect 17736 2604 17785 2632
rect 17736 2592 17742 2604
rect 17773 2601 17785 2604
rect 17819 2601 17831 2635
rect 17773 2595 17831 2601
rect 19610 2592 19616 2644
rect 19668 2632 19674 2644
rect 20438 2632 20444 2644
rect 19668 2604 20444 2632
rect 19668 2592 19674 2604
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 21085 2635 21143 2641
rect 21085 2601 21097 2635
rect 21131 2632 21143 2635
rect 27338 2632 27344 2644
rect 21131 2604 27344 2632
rect 21131 2601 21143 2604
rect 21085 2595 21143 2601
rect 27338 2592 27344 2604
rect 27396 2592 27402 2644
rect 28966 2604 35572 2632
rect 15381 2567 15439 2573
rect 15381 2533 15393 2567
rect 15427 2564 15439 2567
rect 16298 2564 16304 2576
rect 15427 2536 16304 2564
rect 15427 2533 15439 2536
rect 15381 2527 15439 2533
rect 16298 2524 16304 2536
rect 16356 2524 16362 2576
rect 18506 2564 18512 2576
rect 18467 2536 18512 2564
rect 18506 2524 18512 2536
rect 18564 2524 18570 2576
rect 19797 2567 19855 2573
rect 19797 2533 19809 2567
rect 19843 2564 19855 2567
rect 20346 2564 20352 2576
rect 19843 2536 20352 2564
rect 19843 2533 19855 2536
rect 19797 2527 19855 2533
rect 20346 2524 20352 2536
rect 20404 2524 20410 2576
rect 22005 2567 22063 2573
rect 22005 2533 22017 2567
rect 22051 2564 22063 2567
rect 22646 2564 22652 2576
rect 22051 2536 22652 2564
rect 22051 2533 22063 2536
rect 22005 2527 22063 2533
rect 22646 2524 22652 2536
rect 22704 2524 22710 2576
rect 22741 2567 22799 2573
rect 22741 2533 22753 2567
rect 22787 2533 22799 2567
rect 23566 2564 23572 2576
rect 23527 2536 23572 2564
rect 22741 2527 22799 2533
rect 17218 2496 17224 2508
rect 14200 2468 14872 2496
rect 15856 2468 17224 2496
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 1765 2391 1823 2397
rect 1780 2360 1808 2391
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2958 2428 2964 2440
rect 2919 2400 2964 2428
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3050 2388 3056 2440
rect 3108 2428 3114 2440
rect 4062 2428 4068 2440
rect 3108 2400 4068 2428
rect 3108 2388 3114 2400
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 5077 2431 5135 2437
rect 5077 2428 5089 2431
rect 5040 2400 5089 2428
rect 5040 2388 5046 2400
rect 5077 2397 5089 2400
rect 5123 2397 5135 2431
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5077 2391 5135 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7098 2428 7104 2440
rect 6963 2400 7104 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 11514 2428 11520 2440
rect 8588 2400 10548 2428
rect 11475 2400 11520 2428
rect 3694 2360 3700 2372
rect 1780 2332 3700 2360
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 6457 2363 6515 2369
rect 4908 2332 6408 2360
rect 4246 2292 4252 2304
rect 4207 2264 4252 2292
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 4908 2301 4936 2332
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2261 4951 2295
rect 4893 2255 4951 2261
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2292 5687 2295
rect 5810 2292 5816 2304
rect 5675 2264 5816 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 6380 2292 6408 2332
rect 6457 2329 6469 2363
rect 6503 2360 6515 2363
rect 8588 2360 8616 2400
rect 6503 2332 8616 2360
rect 6503 2329 6515 2332
rect 6457 2323 6515 2329
rect 8662 2320 8668 2372
rect 8720 2360 8726 2372
rect 9030 2360 9036 2372
rect 8720 2332 9036 2360
rect 8720 2320 8726 2332
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 9214 2320 9220 2372
rect 9272 2360 9278 2372
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 9272 2332 10149 2360
rect 9272 2320 9278 2332
rect 10137 2329 10149 2332
rect 10183 2329 10195 2363
rect 10520 2360 10548 2400
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2428 12587 2431
rect 12710 2428 12716 2440
rect 12575 2400 12716 2428
rect 12575 2397 12587 2400
rect 12529 2391 12587 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 14200 2437 14228 2468
rect 15856 2437 15884 2468
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 19978 2456 19984 2508
rect 20036 2496 20042 2508
rect 20162 2496 20168 2508
rect 20036 2468 20168 2496
rect 20036 2456 20042 2468
rect 20162 2456 20168 2468
rect 20220 2456 20226 2508
rect 20990 2496 20996 2508
rect 20272 2468 20996 2496
rect 14185 2431 14243 2437
rect 14185 2397 14197 2431
rect 14231 2397 14243 2431
rect 15841 2431 15899 2437
rect 15841 2428 15853 2431
rect 14185 2391 14243 2397
rect 14292 2400 15853 2428
rect 14292 2360 14320 2400
rect 15841 2397 15853 2400
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2397 17003 2431
rect 17954 2428 17960 2440
rect 17915 2400 17960 2428
rect 16945 2391 17003 2397
rect 10520 2332 14320 2360
rect 15197 2363 15255 2369
rect 10137 2323 10195 2329
rect 15197 2329 15209 2363
rect 15243 2360 15255 2363
rect 15470 2360 15476 2372
rect 15243 2332 15476 2360
rect 15243 2329 15255 2332
rect 15197 2323 15255 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 16960 2360 16988 2391
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18693 2431 18751 2437
rect 18693 2397 18705 2431
rect 18739 2428 18751 2431
rect 19518 2428 19524 2440
rect 18739 2400 19524 2428
rect 18739 2397 18751 2400
rect 18693 2391 18751 2397
rect 19518 2388 19524 2400
rect 19576 2428 19582 2440
rect 20272 2428 20300 2468
rect 20990 2456 20996 2468
rect 21048 2456 21054 2508
rect 22756 2496 22784 2527
rect 23566 2524 23572 2536
rect 23624 2524 23630 2576
rect 25777 2567 25835 2573
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 26418 2564 26424 2576
rect 25823 2536 26424 2564
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 26418 2524 26424 2536
rect 26476 2524 26482 2576
rect 27709 2567 27767 2573
rect 27709 2533 27721 2567
rect 27755 2564 27767 2567
rect 28350 2564 28356 2576
rect 27755 2536 28356 2564
rect 27755 2533 27767 2536
rect 27709 2527 27767 2533
rect 28350 2524 28356 2536
rect 28408 2524 28414 2576
rect 28966 2496 28994 2604
rect 35544 2564 35572 2604
rect 35618 2592 35624 2644
rect 35676 2632 35682 2644
rect 37277 2635 37335 2641
rect 37277 2632 37289 2635
rect 35676 2604 37289 2632
rect 35676 2592 35682 2604
rect 37277 2601 37289 2604
rect 37323 2601 37335 2635
rect 42886 2632 42892 2644
rect 37277 2595 37335 2601
rect 37384 2604 42892 2632
rect 36722 2564 36728 2576
rect 35544 2536 36728 2564
rect 36722 2524 36728 2536
rect 36780 2524 36786 2576
rect 37384 2564 37412 2604
rect 42886 2592 42892 2604
rect 42944 2592 42950 2644
rect 51994 2592 52000 2644
rect 52052 2632 52058 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 52052 2604 55321 2632
rect 52052 2592 52058 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 36832 2536 37412 2564
rect 22756 2468 28994 2496
rect 31938 2456 31944 2508
rect 31996 2496 32002 2508
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 31996 2468 32781 2496
rect 31996 2456 32002 2468
rect 32769 2465 32781 2468
rect 32815 2465 32827 2499
rect 32769 2459 32827 2465
rect 33042 2456 33048 2508
rect 33100 2496 33106 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 33100 2468 34713 2496
rect 33100 2456 33106 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 35618 2456 35624 2508
rect 35676 2496 35682 2508
rect 36832 2496 36860 2536
rect 38010 2524 38016 2576
rect 38068 2564 38074 2576
rect 39853 2567 39911 2573
rect 39853 2564 39865 2567
rect 38068 2536 39865 2564
rect 38068 2524 38074 2536
rect 39853 2533 39865 2536
rect 39899 2533 39911 2567
rect 39853 2527 39911 2533
rect 41874 2524 41880 2576
rect 41932 2564 41938 2576
rect 43717 2567 43775 2573
rect 43717 2564 43729 2567
rect 41932 2536 43729 2564
rect 41932 2524 41938 2536
rect 43717 2533 43729 2536
rect 43763 2533 43775 2567
rect 43717 2527 43775 2533
rect 45738 2524 45744 2576
rect 45796 2564 45802 2576
rect 47581 2567 47639 2573
rect 47581 2564 47593 2567
rect 45796 2536 47593 2564
rect 45796 2524 45802 2536
rect 47581 2533 47593 2536
rect 47627 2533 47639 2567
rect 47581 2527 47639 2533
rect 49602 2524 49608 2576
rect 49660 2564 49666 2576
rect 51445 2567 51503 2573
rect 51445 2564 51457 2567
rect 49660 2536 51457 2564
rect 49660 2524 49666 2536
rect 51445 2533 51457 2536
rect 51491 2533 51503 2567
rect 54021 2567 54079 2573
rect 54021 2564 54033 2567
rect 51445 2527 51503 2533
rect 51552 2536 54033 2564
rect 35676 2468 36860 2496
rect 35676 2456 35682 2468
rect 36906 2456 36912 2508
rect 36964 2496 36970 2508
rect 38565 2499 38623 2505
rect 38565 2496 38577 2499
rect 36964 2468 38577 2496
rect 36964 2456 36970 2468
rect 38565 2465 38577 2468
rect 38611 2465 38623 2499
rect 38565 2459 38623 2465
rect 38838 2456 38844 2508
rect 38896 2496 38902 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 38896 2468 40509 2496
rect 38896 2456 38902 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 40770 2456 40776 2508
rect 40828 2496 40834 2508
rect 42429 2499 42487 2505
rect 42429 2496 42441 2499
rect 40828 2468 42441 2496
rect 40828 2456 40834 2468
rect 42429 2465 42441 2468
rect 42475 2465 42487 2499
rect 42429 2459 42487 2465
rect 43254 2456 43260 2508
rect 43312 2496 43318 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 43312 2468 45017 2496
rect 43312 2456 43318 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45005 2459 45063 2465
rect 46566 2456 46572 2508
rect 46624 2496 46630 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 46624 2468 48237 2496
rect 46624 2456 46630 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 48498 2456 48504 2508
rect 48556 2496 48562 2508
rect 50157 2499 50215 2505
rect 50157 2496 50169 2499
rect 48556 2468 50169 2496
rect 48556 2456 48562 2468
rect 50157 2465 50169 2468
rect 50203 2465 50215 2499
rect 50157 2459 50215 2465
rect 51258 2456 51264 2508
rect 51316 2496 51322 2508
rect 51552 2496 51580 2536
rect 54021 2533 54033 2536
rect 54067 2533 54079 2567
rect 54021 2527 54079 2533
rect 54386 2524 54392 2576
rect 54444 2564 54450 2576
rect 56597 2567 56655 2573
rect 56597 2564 56609 2567
rect 54444 2536 56609 2564
rect 54444 2524 54450 2536
rect 56597 2533 56609 2536
rect 56643 2533 56655 2567
rect 56597 2527 56655 2533
rect 51316 2468 51580 2496
rect 51316 2456 51322 2468
rect 52546 2456 52552 2508
rect 52604 2496 52610 2508
rect 53377 2499 53435 2505
rect 53377 2496 53389 2499
rect 52604 2468 53389 2496
rect 52604 2456 52610 2468
rect 53377 2465 53389 2468
rect 53423 2465 53435 2499
rect 53377 2459 53435 2465
rect 53558 2456 53564 2508
rect 53616 2496 53622 2508
rect 57885 2499 57943 2505
rect 57885 2496 57897 2499
rect 53616 2468 57897 2496
rect 53616 2456 53622 2468
rect 57885 2465 57897 2468
rect 57931 2465 57943 2499
rect 57885 2459 57943 2465
rect 19576 2400 20300 2428
rect 20533 2431 20591 2437
rect 19576 2388 19582 2400
rect 20533 2397 20545 2431
rect 20579 2428 20591 2431
rect 20714 2428 20720 2440
rect 20579 2400 20720 2428
rect 20579 2397 20591 2400
rect 20533 2391 20591 2397
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 21266 2428 21272 2440
rect 21227 2400 21272 2428
rect 21266 2388 21272 2400
rect 21324 2388 21330 2440
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22462 2428 22468 2440
rect 22235 2400 22468 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22462 2388 22468 2400
rect 22520 2388 22526 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 18046 2360 18052 2372
rect 16960 2332 18052 2360
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 19613 2363 19671 2369
rect 19613 2329 19625 2363
rect 19659 2360 19671 2363
rect 20254 2360 20260 2372
rect 19659 2332 20260 2360
rect 19659 2329 19671 2332
rect 19613 2323 19671 2329
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 8018 2292 8024 2304
rect 6380 2264 8024 2292
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 10042 2292 10048 2304
rect 9355 2264 10048 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 10042 2252 10048 2264
rect 10100 2252 10106 2304
rect 10410 2292 10416 2304
rect 10371 2264 10416 2292
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 16022 2292 16028 2304
rect 15983 2264 16028 2292
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 20346 2292 20352 2304
rect 20307 2264 20352 2292
rect 20346 2252 20352 2264
rect 20404 2252 20410 2304
rect 22940 2292 22968 2391
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 23348 2400 23397 2428
rect 23348 2388 23354 2400
rect 23385 2397 23397 2400
rect 23431 2428 23443 2431
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23431 2400 24409 2428
rect 23431 2397 23443 2400
rect 23385 2391 23443 2397
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2428 25191 2431
rect 25866 2428 25872 2440
rect 25179 2400 25872 2428
rect 25179 2397 25191 2400
rect 25133 2391 25191 2397
rect 25866 2388 25872 2400
rect 25924 2388 25930 2440
rect 26421 2431 26479 2437
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 27246 2428 27252 2440
rect 26467 2400 27252 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 27246 2388 27252 2400
rect 27304 2388 27310 2440
rect 27338 2388 27344 2440
rect 27396 2428 27402 2440
rect 28353 2431 28411 2437
rect 27396 2400 27752 2428
rect 27396 2388 27402 2400
rect 23566 2320 23572 2372
rect 23624 2360 23630 2372
rect 27724 2360 27752 2400
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28902 2428 28908 2440
rect 28399 2400 28908 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28902 2388 28908 2400
rect 28960 2388 28966 2440
rect 28997 2431 29055 2437
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 29454 2428 29460 2440
rect 29043 2400 29460 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29454 2388 29460 2400
rect 29512 2388 29518 2440
rect 30101 2431 30159 2437
rect 30101 2397 30113 2431
rect 30147 2428 30159 2431
rect 30282 2428 30288 2440
rect 30147 2400 30288 2428
rect 30147 2397 30159 2400
rect 30101 2391 30159 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2428 30803 2431
rect 30834 2428 30840 2440
rect 30791 2400 30840 2428
rect 30791 2397 30803 2400
rect 30745 2391 30803 2397
rect 30834 2388 30840 2400
rect 30892 2388 30898 2440
rect 31110 2388 31116 2440
rect 31168 2428 31174 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 31168 2400 31217 2428
rect 31168 2388 31174 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31444 2400 32137 2428
rect 31444 2388 31450 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32490 2388 32496 2440
rect 32548 2428 32554 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 32548 2400 33425 2428
rect 32548 2388 32554 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 33594 2388 33600 2440
rect 33652 2428 33658 2440
rect 35345 2431 35403 2437
rect 35345 2428 35357 2431
rect 33652 2400 35357 2428
rect 33652 2388 33658 2400
rect 35345 2397 35357 2400
rect 35391 2397 35403 2431
rect 35345 2391 35403 2397
rect 35710 2388 35716 2440
rect 35768 2428 35774 2440
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 35768 2400 36001 2428
rect 35768 2388 35774 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37921 2431 37979 2437
rect 37921 2428 37933 2431
rect 36136 2400 37933 2428
rect 36136 2388 36142 2400
rect 37921 2397 37933 2400
rect 37967 2397 37979 2431
rect 37921 2391 37979 2397
rect 39390 2388 39396 2440
rect 39448 2428 39454 2440
rect 41141 2431 41199 2437
rect 41141 2428 41153 2431
rect 39448 2400 41153 2428
rect 39448 2388 39454 2400
rect 41141 2397 41153 2400
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 41322 2388 41328 2440
rect 41380 2428 41386 2440
rect 43073 2431 43131 2437
rect 43073 2428 43085 2431
rect 41380 2400 43085 2428
rect 41380 2388 41386 2400
rect 43073 2397 43085 2400
rect 43119 2397 43131 2431
rect 43073 2391 43131 2397
rect 43806 2388 43812 2440
rect 43864 2428 43870 2440
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 43864 2400 45661 2428
rect 43864 2388 43870 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 46293 2431 46351 2437
rect 46293 2397 46305 2431
rect 46339 2397 46351 2431
rect 46293 2391 46351 2397
rect 36538 2360 36544 2372
rect 23624 2332 27108 2360
rect 27724 2332 36544 2360
rect 23624 2320 23630 2332
rect 23014 2292 23020 2304
rect 22927 2264 23020 2292
rect 23014 2252 23020 2264
rect 23072 2292 23078 2304
rect 26973 2295 27031 2301
rect 26973 2292 26985 2295
rect 23072 2264 26985 2292
rect 23072 2252 23078 2264
rect 26973 2261 26985 2264
rect 27019 2261 27031 2295
rect 27080 2292 27108 2332
rect 36538 2320 36544 2332
rect 36596 2320 36602 2372
rect 36722 2320 36728 2372
rect 36780 2360 36786 2372
rect 43162 2360 43168 2372
rect 36780 2332 43168 2360
rect 36780 2320 36786 2332
rect 43162 2320 43168 2332
rect 43220 2320 43226 2372
rect 44634 2320 44640 2372
rect 44692 2360 44698 2372
rect 46308 2360 46336 2391
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 48869 2431 48927 2437
rect 48869 2428 48881 2431
rect 47176 2400 48881 2428
rect 47176 2388 47182 2400
rect 48869 2397 48881 2400
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 49050 2388 49056 2440
rect 49108 2428 49114 2440
rect 50801 2431 50859 2437
rect 50801 2428 50813 2431
rect 49108 2400 50813 2428
rect 49108 2388 49114 2400
rect 50801 2397 50813 2400
rect 50847 2397 50859 2431
rect 50801 2391 50859 2397
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 50948 2400 52745 2428
rect 50948 2388 50954 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 52733 2391 52791 2397
rect 55953 2431 56011 2437
rect 55953 2397 55965 2431
rect 55999 2397 56011 2431
rect 55953 2391 56011 2397
rect 44692 2332 46336 2360
rect 44692 2320 44698 2332
rect 52362 2320 52368 2372
rect 52420 2360 52426 2372
rect 55968 2360 55996 2391
rect 52420 2332 55996 2360
rect 52420 2320 52426 2332
rect 56318 2292 56324 2304
rect 27080 2264 56324 2292
rect 26973 2255 27031 2261
rect 56318 2252 56324 2264
rect 56376 2252 56382 2304
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 5810 2048 5816 2100
rect 5868 2088 5874 2100
rect 8294 2088 8300 2100
rect 5868 2060 8300 2088
rect 5868 2048 5874 2060
rect 8294 2048 8300 2060
rect 8352 2048 8358 2100
rect 18782 2088 18788 2100
rect 8404 2060 18788 2088
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 7650 2020 7656 2032
rect 4120 1992 7656 2020
rect 4120 1980 4126 1992
rect 7650 1980 7656 1992
rect 7708 1980 7714 2032
rect 6822 1912 6828 1964
rect 6880 1952 6886 1964
rect 7098 1952 7104 1964
rect 6880 1924 7104 1952
rect 6880 1912 6886 1924
rect 7098 1912 7104 1924
rect 7156 1912 7162 1964
rect 4246 1844 4252 1896
rect 4304 1884 4310 1896
rect 8404 1884 8432 2060
rect 18782 2048 18788 2060
rect 18840 2048 18846 2100
rect 22646 2048 22652 2100
rect 22704 2088 22710 2100
rect 35618 2088 35624 2100
rect 22704 2060 35624 2088
rect 22704 2048 22710 2060
rect 35618 2048 35624 2060
rect 35676 2048 35682 2100
rect 36538 2048 36544 2100
rect 36596 2088 36602 2100
rect 44726 2088 44732 2100
rect 36596 2060 44732 2088
rect 36596 2048 36602 2060
rect 44726 2048 44732 2060
rect 44784 2048 44790 2100
rect 52730 2048 52736 2100
rect 52788 2048 52794 2100
rect 52914 2048 52920 2100
rect 52972 2088 52978 2100
rect 54386 2088 54392 2100
rect 52972 2060 54392 2088
rect 52972 2048 52978 2060
rect 54386 2048 54392 2060
rect 54444 2048 54450 2100
rect 10042 1980 10048 2032
rect 10100 2020 10106 2032
rect 12894 2020 12900 2032
rect 10100 1992 12900 2020
rect 10100 1980 10106 1992
rect 12894 1980 12900 1992
rect 12952 1980 12958 2032
rect 20346 1980 20352 2032
rect 20404 2020 20410 2032
rect 43438 2020 43444 2032
rect 20404 1992 43444 2020
rect 20404 1980 20410 1992
rect 43438 1980 43444 1992
rect 43496 1980 43502 2032
rect 4304 1856 8432 1884
rect 4304 1844 4310 1856
rect 10410 1844 10416 1896
rect 10468 1884 10474 1896
rect 29546 1884 29552 1896
rect 10468 1856 29552 1884
rect 10468 1844 10474 1856
rect 29546 1844 29552 1856
rect 29604 1844 29610 1896
rect 5902 1776 5908 1828
rect 5960 1816 5966 1828
rect 6638 1816 6644 1828
rect 5960 1788 6644 1816
rect 5960 1776 5966 1788
rect 6638 1776 6644 1788
rect 6696 1776 6702 1828
rect 15470 1708 15476 1760
rect 15528 1748 15534 1760
rect 16390 1748 16396 1760
rect 15528 1720 16396 1748
rect 15528 1708 15534 1720
rect 16390 1708 16396 1720
rect 16448 1708 16454 1760
rect 20714 1708 20720 1760
rect 20772 1748 20778 1760
rect 21082 1748 21088 1760
rect 20772 1720 21088 1748
rect 20772 1708 20778 1720
rect 21082 1708 21088 1720
rect 21140 1708 21146 1760
rect 21266 1708 21272 1760
rect 21324 1748 21330 1760
rect 21910 1748 21916 1760
rect 21324 1720 21916 1748
rect 21324 1708 21330 1720
rect 21910 1708 21916 1720
rect 21968 1708 21974 1760
rect 5350 1572 5356 1624
rect 5408 1612 5414 1624
rect 5902 1612 5908 1624
rect 5408 1584 5908 1612
rect 5408 1572 5414 1584
rect 5902 1572 5908 1584
rect 5960 1572 5966 1624
rect 13998 1436 14004 1488
rect 14056 1476 14062 1488
rect 15010 1476 15016 1488
rect 14056 1448 15016 1476
rect 14056 1436 14062 1448
rect 15010 1436 15016 1448
rect 15068 1436 15074 1488
rect 19334 1436 19340 1488
rect 19392 1476 19398 1488
rect 19794 1476 19800 1488
rect 19392 1448 19800 1476
rect 19392 1436 19398 1448
rect 19794 1436 19800 1448
rect 19852 1436 19858 1488
rect 4614 1368 4620 1420
rect 4672 1408 4678 1420
rect 5718 1408 5724 1420
rect 4672 1380 5724 1408
rect 4672 1368 4678 1380
rect 5718 1368 5724 1380
rect 5776 1368 5782 1420
rect 14274 1368 14280 1420
rect 14332 1408 14338 1420
rect 14734 1408 14740 1420
rect 14332 1380 14740 1408
rect 14332 1368 14338 1380
rect 14734 1368 14740 1380
rect 14792 1368 14798 1420
rect 19702 1368 19708 1420
rect 19760 1408 19766 1420
rect 20162 1408 20168 1420
rect 19760 1380 20168 1408
rect 19760 1368 19766 1380
rect 20162 1368 20168 1380
rect 20220 1368 20226 1420
rect 34146 1368 34152 1420
rect 34204 1408 34210 1420
rect 35710 1408 35716 1420
rect 34204 1380 35716 1408
rect 34204 1368 34210 1380
rect 35710 1368 35716 1380
rect 35768 1368 35774 1420
rect 4798 1300 4804 1352
rect 4856 1340 4862 1352
rect 6178 1340 6184 1352
rect 4856 1312 6184 1340
rect 4856 1300 4862 1312
rect 6178 1300 6184 1312
rect 6236 1300 6242 1352
rect 19426 1300 19432 1352
rect 19484 1340 19490 1352
rect 19610 1340 19616 1352
rect 19484 1312 19616 1340
rect 19484 1300 19490 1312
rect 19610 1300 19616 1312
rect 19668 1300 19674 1352
rect 52748 1340 52776 2048
rect 52822 1436 52828 1488
rect 52880 1476 52886 1488
rect 53006 1476 53012 1488
rect 52880 1448 53012 1476
rect 52880 1436 52886 1448
rect 53006 1436 53012 1448
rect 53064 1436 53070 1488
rect 53006 1340 53012 1352
rect 52748 1312 53012 1340
rect 53006 1300 53012 1312
rect 53064 1300 53070 1352
rect 52546 1136 52552 1148
rect 51000 1108 52552 1136
rect 51000 944 51028 1108
rect 52546 1096 52552 1108
rect 52604 1096 52610 1148
rect 52546 960 52552 1012
rect 52604 1000 52610 1012
rect 54754 1000 54760 1012
rect 52604 972 54760 1000
rect 52604 960 52610 972
rect 54754 960 54760 972
rect 54812 960 54818 1012
rect 50982 892 50988 944
rect 51040 892 51046 944
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 12716 57536 12768 57588
rect 14280 57536 14332 57588
rect 15844 57536 15896 57588
rect 17408 57536 17460 57588
rect 19340 57536 19392 57588
rect 20720 57536 20772 57588
rect 22100 57536 22152 57588
rect 23664 57536 23716 57588
rect 25228 57536 25280 57588
rect 26792 57536 26844 57588
rect 28356 57536 28408 57588
rect 29920 57536 29972 57588
rect 31484 57536 31536 57588
rect 33140 57536 33192 57588
rect 34612 57536 34664 57588
rect 36176 57536 36228 57588
rect 37740 57536 37792 57588
rect 39304 57536 39356 57588
rect 40868 57536 40920 57588
rect 42432 57536 42484 57588
rect 44180 57536 44232 57588
rect 45560 57536 45612 57588
rect 47124 57536 47176 57588
rect 48688 57536 48740 57588
rect 50160 57536 50212 57588
rect 51816 57536 51868 57588
rect 53380 57536 53432 57588
rect 54944 57536 54996 57588
rect 56600 57536 56652 57588
rect 58072 57579 58124 57588
rect 58072 57545 58081 57579
rect 58081 57545 58115 57579
rect 58115 57545 58124 57579
rect 58072 57536 58124 57545
rect 20904 57468 20956 57520
rect 1768 57400 1820 57452
rect 3332 57400 3384 57452
rect 4896 57400 4948 57452
rect 6460 57400 6512 57452
rect 8024 57400 8076 57452
rect 9680 57443 9732 57452
rect 9680 57409 9689 57443
rect 9689 57409 9723 57443
rect 9723 57409 9732 57443
rect 9680 57400 9732 57409
rect 11152 57400 11204 57452
rect 13084 57443 13136 57452
rect 13084 57409 13093 57443
rect 13093 57409 13127 57443
rect 13127 57409 13136 57443
rect 13084 57400 13136 57409
rect 14648 57443 14700 57452
rect 14648 57409 14657 57443
rect 14657 57409 14691 57443
rect 14691 57409 14700 57443
rect 14648 57400 14700 57409
rect 16672 57443 16724 57452
rect 16672 57409 16681 57443
rect 16681 57409 16715 57443
rect 16715 57409 16724 57443
rect 16672 57400 16724 57409
rect 17500 57443 17552 57452
rect 17500 57409 17509 57443
rect 17509 57409 17543 57443
rect 17543 57409 17552 57443
rect 17500 57400 17552 57409
rect 19248 57443 19300 57452
rect 19248 57409 19257 57443
rect 19257 57409 19291 57443
rect 19291 57409 19300 57443
rect 19248 57400 19300 57409
rect 20628 57443 20680 57452
rect 20628 57409 20637 57443
rect 20637 57409 20671 57443
rect 20671 57409 20680 57443
rect 20628 57400 20680 57409
rect 22192 57443 22244 57452
rect 22192 57409 22201 57443
rect 22201 57409 22235 57443
rect 22235 57409 22244 57443
rect 22192 57400 22244 57409
rect 24400 57443 24452 57452
rect 24400 57409 24409 57443
rect 24409 57409 24443 57443
rect 24443 57409 24452 57443
rect 24400 57400 24452 57409
rect 31760 57468 31812 57520
rect 28448 57443 28500 57452
rect 19340 57332 19392 57384
rect 28448 57409 28457 57443
rect 28457 57409 28491 57443
rect 28491 57409 28500 57443
rect 28448 57400 28500 57409
rect 29000 57400 29052 57452
rect 32128 57443 32180 57452
rect 32128 57409 32137 57443
rect 32137 57409 32171 57443
rect 32171 57409 32180 57443
rect 32128 57400 32180 57409
rect 33140 57443 33192 57452
rect 33140 57409 33149 57443
rect 33149 57409 33183 57443
rect 33183 57409 33192 57443
rect 33140 57400 33192 57409
rect 34704 57443 34756 57452
rect 34704 57409 34713 57443
rect 34713 57409 34747 57443
rect 34747 57409 34756 57443
rect 34704 57400 34756 57409
rect 46204 57468 46256 57520
rect 37832 57443 37884 57452
rect 37832 57409 37841 57443
rect 37841 57409 37875 57443
rect 37875 57409 37884 57443
rect 37832 57400 37884 57409
rect 39856 57443 39908 57452
rect 39856 57409 39865 57443
rect 39865 57409 39899 57443
rect 39899 57409 39908 57443
rect 39856 57400 39908 57409
rect 42524 57443 42576 57452
rect 22284 57196 22336 57248
rect 40776 57332 40828 57384
rect 42524 57409 42533 57443
rect 42533 57409 42567 57443
rect 42567 57409 42576 57443
rect 42524 57400 42576 57409
rect 44088 57443 44140 57452
rect 44088 57409 44097 57443
rect 44097 57409 44131 57443
rect 44131 57409 44140 57443
rect 44088 57400 44140 57409
rect 44180 57400 44232 57452
rect 47584 57443 47636 57452
rect 47584 57409 47593 57443
rect 47593 57409 47627 57443
rect 47627 57409 47636 57443
rect 47584 57400 47636 57409
rect 47676 57400 47728 57452
rect 53472 57443 53524 57452
rect 48320 57332 48372 57384
rect 53472 57409 53481 57443
rect 53481 57409 53515 57443
rect 53515 57409 53524 57443
rect 53472 57400 53524 57409
rect 55312 57443 55364 57452
rect 55312 57409 55321 57443
rect 55321 57409 55355 57443
rect 55355 57409 55364 57443
rect 55312 57400 55364 57409
rect 56048 57400 56100 57452
rect 57796 57400 57848 57452
rect 56048 57239 56100 57248
rect 56048 57205 56057 57239
rect 56057 57205 56091 57239
rect 56091 57205 56100 57239
rect 56048 57196 56100 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 21088 56992 21140 57044
rect 40776 57035 40828 57044
rect 40776 57001 40785 57035
rect 40785 57001 40819 57035
rect 40819 57001 40828 57035
rect 40776 56992 40828 57001
rect 57520 57035 57572 57044
rect 57520 57001 57529 57035
rect 57529 57001 57563 57035
rect 57563 57001 57572 57035
rect 57520 56992 57572 57001
rect 42524 56924 42576 56976
rect 57888 56788 57940 56840
rect 16488 56652 16540 56704
rect 28080 56695 28132 56704
rect 28080 56661 28089 56695
rect 28089 56661 28123 56695
rect 28123 56661 28132 56695
rect 28080 56652 28132 56661
rect 29184 56652 29236 56704
rect 45468 56652 45520 56704
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 13084 56448 13136 56500
rect 14648 56448 14700 56500
rect 16672 56448 16724 56500
rect 17500 56448 17552 56500
rect 20628 56448 20680 56500
rect 22284 56491 22336 56500
rect 22284 56457 22293 56491
rect 22293 56457 22327 56491
rect 22327 56457 22336 56491
rect 22284 56448 22336 56457
rect 24400 56448 24452 56500
rect 28448 56448 28500 56500
rect 32128 56448 32180 56500
rect 33140 56448 33192 56500
rect 34704 56448 34756 56500
rect 37832 56448 37884 56500
rect 19340 56380 19392 56432
rect 21088 56423 21140 56432
rect 21088 56389 21097 56423
rect 21097 56389 21131 56423
rect 21131 56389 21140 56423
rect 21088 56380 21140 56389
rect 14188 56312 14240 56364
rect 15108 56312 15160 56364
rect 16488 56312 16540 56364
rect 16580 56312 16632 56364
rect 17224 56312 17276 56364
rect 17868 56312 17920 56364
rect 18604 56355 18656 56364
rect 18604 56321 18613 56355
rect 18613 56321 18647 56355
rect 18647 56321 18656 56355
rect 18604 56312 18656 56321
rect 19064 56312 19116 56364
rect 20352 56312 20404 56364
rect 21916 56312 21968 56364
rect 23112 56355 23164 56364
rect 23112 56321 23121 56355
rect 23121 56321 23155 56355
rect 23155 56321 23164 56355
rect 23112 56312 23164 56321
rect 20168 56244 20220 56296
rect 28080 56380 28132 56432
rect 44180 56448 44232 56500
rect 46204 56448 46256 56500
rect 47584 56448 47636 56500
rect 53472 56380 53524 56432
rect 19248 56176 19300 56228
rect 20904 56176 20956 56228
rect 20352 56151 20404 56160
rect 20352 56117 20361 56151
rect 20361 56117 20395 56151
rect 20395 56117 20404 56151
rect 20352 56108 20404 56117
rect 23572 56108 23624 56160
rect 29184 56355 29236 56364
rect 29184 56321 29193 56355
rect 29193 56321 29227 56355
rect 29227 56321 29236 56355
rect 29184 56312 29236 56321
rect 30012 56312 30064 56364
rect 30840 56312 30892 56364
rect 32128 56355 32180 56364
rect 32128 56321 32137 56355
rect 32137 56321 32171 56355
rect 32171 56321 32180 56355
rect 32128 56312 32180 56321
rect 33600 56355 33652 56364
rect 33600 56321 33609 56355
rect 33609 56321 33643 56355
rect 33643 56321 33652 56355
rect 33600 56312 33652 56321
rect 35808 56355 35860 56364
rect 35808 56321 35817 56355
rect 35817 56321 35851 56355
rect 35851 56321 35860 56355
rect 35808 56312 35860 56321
rect 42892 56355 42944 56364
rect 42892 56321 42901 56355
rect 42901 56321 42935 56355
rect 42935 56321 42944 56355
rect 42892 56312 42944 56321
rect 43536 56355 43588 56364
rect 43536 56321 43545 56355
rect 43545 56321 43579 56355
rect 43579 56321 43588 56355
rect 43536 56312 43588 56321
rect 43996 56312 44048 56364
rect 44732 56312 44784 56364
rect 45468 56355 45520 56364
rect 45468 56321 45477 56355
rect 45477 56321 45511 56355
rect 45511 56321 45520 56355
rect 45468 56312 45520 56321
rect 46112 56355 46164 56364
rect 46112 56321 46121 56355
rect 46121 56321 46155 56355
rect 46155 56321 46164 56355
rect 46112 56312 46164 56321
rect 46756 56355 46808 56364
rect 46756 56321 46765 56355
rect 46765 56321 46799 56355
rect 46799 56321 46808 56355
rect 46756 56312 46808 56321
rect 58440 56312 58492 56364
rect 29000 56176 29052 56228
rect 44088 56176 44140 56228
rect 55312 56244 55364 56296
rect 48320 56176 48372 56228
rect 30840 56151 30892 56160
rect 30840 56117 30849 56151
rect 30849 56117 30883 56151
rect 30883 56117 30892 56151
rect 30840 56108 30892 56117
rect 31760 56108 31812 56160
rect 47676 56108 47728 56160
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 17868 55947 17920 55956
rect 17868 55913 17877 55947
rect 17877 55913 17911 55947
rect 17911 55913 17920 55947
rect 17868 55904 17920 55913
rect 22192 55904 22244 55956
rect 16396 55632 16448 55684
rect 18604 55632 18656 55684
rect 27620 55743 27672 55752
rect 27620 55709 27629 55743
rect 27629 55709 27663 55743
rect 27663 55709 27672 55743
rect 27620 55700 27672 55709
rect 14188 55607 14240 55616
rect 14188 55573 14197 55607
rect 14197 55573 14231 55607
rect 14231 55573 14240 55607
rect 14188 55564 14240 55573
rect 15108 55607 15160 55616
rect 15108 55573 15117 55607
rect 15117 55573 15151 55607
rect 15151 55573 15160 55607
rect 15108 55564 15160 55573
rect 16580 55607 16632 55616
rect 16580 55573 16589 55607
rect 16589 55573 16623 55607
rect 16623 55573 16632 55607
rect 17224 55607 17276 55616
rect 16580 55564 16632 55573
rect 17224 55573 17233 55607
rect 17233 55573 17267 55607
rect 17267 55573 17276 55607
rect 17224 55564 17276 55573
rect 19064 55564 19116 55616
rect 20444 55607 20496 55616
rect 20444 55573 20453 55607
rect 20453 55573 20487 55607
rect 20487 55573 20496 55607
rect 20444 55564 20496 55573
rect 21916 55607 21968 55616
rect 21916 55573 21925 55607
rect 21925 55573 21959 55607
rect 21959 55573 21968 55607
rect 21916 55564 21968 55573
rect 39856 55632 39908 55684
rect 30012 55607 30064 55616
rect 30012 55573 30021 55607
rect 30021 55573 30055 55607
rect 30055 55573 30064 55607
rect 30012 55564 30064 55573
rect 42892 55564 42944 55616
rect 43536 55564 43588 55616
rect 43996 55607 44048 55616
rect 43996 55573 44005 55607
rect 44005 55573 44039 55607
rect 44039 55573 44048 55607
rect 43996 55564 44048 55573
rect 44732 55564 44784 55616
rect 46112 55564 46164 55616
rect 46756 55564 46808 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 23940 55360 23992 55412
rect 43996 55360 44048 55412
rect 58164 55131 58216 55140
rect 58164 55097 58173 55131
rect 58173 55097 58207 55131
rect 58207 55097 58216 55131
rect 58164 55088 58216 55097
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 57888 53932 57940 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 57888 52436 57940 52488
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 43168 51391 43220 51400
rect 43168 51357 43177 51391
rect 43177 51357 43211 51391
rect 43211 51357 43220 51391
rect 43168 51348 43220 51357
rect 58164 51391 58216 51400
rect 58164 51357 58173 51391
rect 58173 51357 58207 51391
rect 58207 51357 58216 51391
rect 58164 51348 58216 51357
rect 56048 51212 56100 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 58164 49759 58216 49768
rect 58164 49725 58173 49759
rect 58173 49725 58207 49759
rect 58207 49725 58216 49759
rect 58164 49716 58216 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 58164 48535 58216 48544
rect 58164 48501 58173 48535
rect 58173 48501 58207 48535
rect 58207 48501 58216 48535
rect 58164 48492 58216 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 58164 47039 58216 47048
rect 58164 47005 58173 47039
rect 58173 47005 58207 47039
rect 58207 47005 58216 47039
rect 58164 46996 58216 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 58164 45951 58216 45960
rect 58164 45917 58173 45951
rect 58173 45917 58207 45951
rect 58207 45917 58216 45951
rect 58164 45908 58216 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 56324 45475 56376 45484
rect 56324 45441 56333 45475
rect 56333 45441 56367 45475
rect 56367 45441 56376 45475
rect 56324 45432 56376 45441
rect 57796 45296 57848 45348
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 58164 44251 58216 44260
rect 58164 44217 58173 44251
rect 58173 44217 58207 44251
rect 58207 44217 58216 44251
rect 58164 44208 58216 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 58164 43095 58216 43104
rect 58164 43061 58173 43095
rect 58173 43061 58207 43095
rect 58207 43061 58216 43095
rect 58164 43052 58216 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 16948 42712 17000 42764
rect 20444 42712 20496 42764
rect 17224 42508 17276 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 12532 42168 12584 42220
rect 15016 42211 15068 42220
rect 15016 42177 15025 42211
rect 15025 42177 15059 42211
rect 15059 42177 15068 42211
rect 15016 42168 15068 42177
rect 15200 42211 15252 42220
rect 15200 42177 15209 42211
rect 15209 42177 15243 42211
rect 15243 42177 15252 42211
rect 15200 42168 15252 42177
rect 12716 42100 12768 42152
rect 17224 42168 17276 42220
rect 15568 42100 15620 42152
rect 12440 42032 12492 42084
rect 12808 41964 12860 42016
rect 15660 42007 15712 42016
rect 15660 41973 15669 42007
rect 15669 41973 15703 42007
rect 15703 41973 15712 42007
rect 15660 41964 15712 41973
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 15200 41760 15252 41812
rect 11520 41735 11572 41744
rect 11520 41701 11529 41735
rect 11529 41701 11563 41735
rect 11563 41701 11572 41735
rect 11520 41692 11572 41701
rect 12716 41692 12768 41744
rect 12900 41624 12952 41676
rect 11704 41531 11756 41540
rect 11704 41497 11713 41531
rect 11713 41497 11747 41531
rect 11747 41497 11756 41531
rect 11704 41488 11756 41497
rect 12992 41599 13044 41608
rect 12992 41565 13001 41599
rect 13001 41565 13035 41599
rect 13035 41565 13044 41599
rect 12992 41556 13044 41565
rect 14740 41556 14792 41608
rect 15016 41556 15068 41608
rect 16580 41624 16632 41676
rect 13820 41488 13872 41540
rect 9680 41463 9732 41472
rect 9680 41429 9689 41463
rect 9689 41429 9723 41463
rect 9723 41429 9732 41463
rect 9680 41420 9732 41429
rect 12348 41463 12400 41472
rect 12348 41429 12357 41463
rect 12357 41429 12391 41463
rect 12391 41429 12400 41463
rect 12348 41420 12400 41429
rect 12440 41420 12492 41472
rect 15200 41488 15252 41540
rect 15568 41488 15620 41540
rect 14556 41420 14608 41472
rect 16764 41488 16816 41540
rect 19892 41692 19944 41744
rect 17224 41556 17276 41608
rect 20352 41624 20404 41676
rect 19892 41599 19944 41608
rect 19340 41488 19392 41540
rect 19892 41565 19901 41599
rect 19901 41565 19935 41599
rect 19935 41565 19944 41599
rect 19892 41556 19944 41565
rect 58164 41599 58216 41608
rect 58164 41565 58173 41599
rect 58173 41565 58207 41599
rect 58207 41565 58216 41599
rect 58164 41556 58216 41565
rect 19432 41420 19484 41472
rect 20168 41488 20220 41540
rect 24400 41420 24452 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 9956 41216 10008 41268
rect 18512 41216 18564 41268
rect 23020 41216 23072 41268
rect 9864 41148 9916 41200
rect 14648 41148 14700 41200
rect 9404 41123 9456 41132
rect 9404 41089 9413 41123
rect 9413 41089 9447 41123
rect 9447 41089 9456 41123
rect 9404 41080 9456 41089
rect 9680 41012 9732 41064
rect 10324 41080 10376 41132
rect 10876 41080 10928 41132
rect 10416 40944 10468 40996
rect 12808 41123 12860 41132
rect 12808 41089 12822 41123
rect 12822 41089 12856 41123
rect 12856 41089 12860 41123
rect 12808 41080 12860 41089
rect 12992 41123 13044 41132
rect 12992 41089 13001 41123
rect 13001 41089 13035 41123
rect 13035 41089 13044 41123
rect 14740 41123 14792 41132
rect 12992 41080 13044 41089
rect 14740 41089 14749 41123
rect 14749 41089 14783 41123
rect 14783 41089 14792 41123
rect 14740 41080 14792 41089
rect 17776 41148 17828 41200
rect 19432 41191 19484 41200
rect 19432 41157 19450 41191
rect 19450 41157 19484 41191
rect 19432 41148 19484 41157
rect 24768 41148 24820 41200
rect 12900 41012 12952 41064
rect 15568 41012 15620 41064
rect 14740 40944 14792 40996
rect 15016 40944 15068 40996
rect 20076 41080 20128 41132
rect 20720 41080 20772 41132
rect 22100 41080 22152 41132
rect 23388 41080 23440 41132
rect 8944 40919 8996 40928
rect 8944 40885 8953 40919
rect 8953 40885 8987 40919
rect 8987 40885 8996 40919
rect 8944 40876 8996 40885
rect 10140 40876 10192 40928
rect 11796 40876 11848 40928
rect 15384 40919 15436 40928
rect 15384 40885 15393 40919
rect 15393 40885 15427 40919
rect 15427 40885 15436 40919
rect 15384 40876 15436 40885
rect 17960 40876 18012 40928
rect 19340 40876 19392 40928
rect 20628 40944 20680 40996
rect 19800 40876 19852 40928
rect 22652 40876 22704 40928
rect 23020 40876 23072 40928
rect 26608 40876 26660 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 14648 40672 14700 40724
rect 20168 40672 20220 40724
rect 4896 40604 4948 40656
rect 9680 40604 9732 40656
rect 14280 40604 14332 40656
rect 19524 40604 19576 40656
rect 12992 40536 13044 40588
rect 4252 40511 4304 40520
rect 4252 40477 4266 40511
rect 4266 40477 4300 40511
rect 4300 40477 4304 40511
rect 4252 40468 4304 40477
rect 4804 40468 4856 40520
rect 6092 40511 6144 40520
rect 6092 40477 6101 40511
rect 6101 40477 6135 40511
rect 6135 40477 6144 40511
rect 6092 40468 6144 40477
rect 9956 40511 10008 40520
rect 9956 40477 9965 40511
rect 9965 40477 9999 40511
rect 9999 40477 10008 40511
rect 9956 40468 10008 40477
rect 3792 40375 3844 40384
rect 3792 40341 3801 40375
rect 3801 40341 3835 40375
rect 3835 40341 3844 40375
rect 3792 40332 3844 40341
rect 4896 40443 4948 40452
rect 4896 40409 4905 40443
rect 4905 40409 4939 40443
rect 4939 40409 4948 40443
rect 4896 40400 4948 40409
rect 5816 40400 5868 40452
rect 5448 40332 5500 40384
rect 5724 40332 5776 40384
rect 7196 40400 7248 40452
rect 9864 40400 9916 40452
rect 10140 40511 10192 40520
rect 10140 40477 10149 40511
rect 10149 40477 10183 40511
rect 10183 40477 10192 40511
rect 10140 40468 10192 40477
rect 10416 40468 10468 40520
rect 10876 40468 10928 40520
rect 14464 40468 14516 40520
rect 16120 40468 16172 40520
rect 17960 40468 18012 40520
rect 19432 40468 19484 40520
rect 19984 40604 20036 40656
rect 20352 40604 20404 40656
rect 20628 40536 20680 40588
rect 10508 40400 10560 40452
rect 6920 40332 6972 40384
rect 8116 40332 8168 40384
rect 9680 40375 9732 40384
rect 9680 40341 9689 40375
rect 9689 40341 9723 40375
rect 9723 40341 9732 40375
rect 9680 40332 9732 40341
rect 10784 40375 10836 40384
rect 10784 40341 10793 40375
rect 10793 40341 10827 40375
rect 10827 40341 10836 40375
rect 10784 40332 10836 40341
rect 11060 40332 11112 40384
rect 13176 40400 13228 40452
rect 14740 40443 14792 40452
rect 14740 40409 14749 40443
rect 14749 40409 14783 40443
rect 14783 40409 14792 40443
rect 14740 40400 14792 40409
rect 15660 40443 15712 40452
rect 15660 40409 15694 40443
rect 15694 40409 15712 40443
rect 15660 40400 15712 40409
rect 19800 40468 19852 40520
rect 19892 40511 19944 40520
rect 19892 40477 19901 40511
rect 19901 40477 19935 40511
rect 19935 40477 19944 40511
rect 19892 40468 19944 40477
rect 20444 40468 20496 40520
rect 22284 40468 22336 40520
rect 22744 40511 22796 40520
rect 22744 40477 22753 40511
rect 22753 40477 22787 40511
rect 22787 40477 22796 40511
rect 22744 40468 22796 40477
rect 16764 40375 16816 40384
rect 16764 40341 16773 40375
rect 16773 40341 16807 40375
rect 16807 40341 16816 40375
rect 16764 40332 16816 40341
rect 19248 40375 19300 40384
rect 19248 40341 19257 40375
rect 19257 40341 19291 40375
rect 19291 40341 19300 40375
rect 19248 40332 19300 40341
rect 20352 40400 20404 40452
rect 21364 40400 21416 40452
rect 21916 40400 21968 40452
rect 23020 40468 23072 40520
rect 27252 40511 27304 40520
rect 27252 40477 27261 40511
rect 27261 40477 27295 40511
rect 27295 40477 27304 40511
rect 27252 40468 27304 40477
rect 58164 40511 58216 40520
rect 58164 40477 58173 40511
rect 58173 40477 58207 40511
rect 58207 40477 58216 40511
rect 58164 40468 58216 40477
rect 27160 40400 27212 40452
rect 20720 40332 20772 40384
rect 22560 40332 22612 40384
rect 23480 40332 23532 40384
rect 23664 40375 23716 40384
rect 23664 40341 23673 40375
rect 23673 40341 23707 40375
rect 23707 40341 23716 40375
rect 23664 40332 23716 40341
rect 28172 40332 28224 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 3792 40060 3844 40112
rect 4252 40128 4304 40180
rect 5816 40171 5868 40180
rect 4988 40060 5040 40112
rect 5816 40137 5825 40171
rect 5825 40137 5859 40171
rect 5859 40137 5868 40171
rect 5816 40128 5868 40137
rect 12532 40128 12584 40180
rect 12900 40171 12952 40180
rect 12900 40137 12909 40171
rect 12909 40137 12943 40171
rect 12943 40137 12952 40171
rect 12900 40128 12952 40137
rect 13544 40128 13596 40180
rect 14740 40171 14792 40180
rect 14740 40137 14749 40171
rect 14749 40137 14783 40171
rect 14783 40137 14792 40171
rect 14740 40128 14792 40137
rect 19248 40128 19300 40180
rect 19524 40128 19576 40180
rect 6920 40060 6972 40112
rect 9864 40060 9916 40112
rect 4712 40035 4764 40044
rect 4712 40001 4721 40035
rect 4721 40001 4755 40035
rect 4755 40001 4764 40035
rect 4712 39992 4764 40001
rect 4804 39992 4856 40044
rect 5448 40035 5500 40044
rect 5448 40001 5460 40035
rect 5460 40001 5494 40035
rect 5494 40001 5500 40035
rect 5448 39992 5500 40001
rect 5724 39992 5776 40044
rect 6736 40035 6788 40044
rect 6736 40001 6745 40035
rect 6745 40001 6779 40035
rect 6779 40001 6788 40035
rect 6736 39992 6788 40001
rect 8944 39992 8996 40044
rect 10784 40060 10836 40112
rect 11796 40103 11848 40112
rect 11796 40069 11830 40103
rect 11830 40069 11848 40103
rect 11796 40060 11848 40069
rect 15384 40060 15436 40112
rect 17408 40060 17460 40112
rect 22100 40128 22152 40180
rect 22192 40128 22244 40180
rect 10416 40035 10468 40044
rect 1860 39924 1912 39976
rect 6092 39924 6144 39976
rect 10416 40001 10425 40035
rect 10425 40001 10459 40035
rect 10459 40001 10468 40035
rect 10416 39992 10468 40001
rect 16120 40035 16172 40044
rect 16120 40001 16129 40035
rect 16129 40001 16163 40035
rect 16163 40001 16172 40035
rect 16120 39992 16172 40001
rect 22560 40060 22612 40112
rect 22284 39992 22336 40044
rect 22652 40035 22704 40044
rect 22652 40001 22661 40035
rect 22661 40001 22695 40035
rect 22695 40001 22704 40035
rect 22652 39992 22704 40001
rect 23664 40128 23716 40180
rect 30840 40128 30892 40180
rect 28172 40103 28224 40112
rect 28172 40069 28181 40103
rect 28181 40069 28215 40103
rect 28215 40069 28224 40103
rect 28172 40060 28224 40069
rect 29184 40060 29236 40112
rect 8576 39831 8628 39840
rect 8576 39797 8585 39831
rect 8585 39797 8619 39831
rect 8619 39797 8628 39831
rect 8576 39788 8628 39797
rect 9772 39831 9824 39840
rect 9772 39797 9781 39831
rect 9781 39797 9815 39831
rect 9815 39797 9824 39831
rect 9772 39788 9824 39797
rect 10968 39831 11020 39840
rect 10968 39797 10977 39831
rect 10977 39797 11011 39831
rect 11011 39797 11020 39831
rect 10968 39788 11020 39797
rect 21916 39924 21968 39976
rect 30564 40035 30616 40044
rect 30564 40001 30573 40035
rect 30573 40001 30607 40035
rect 30607 40001 30616 40035
rect 30564 39992 30616 40001
rect 25044 39924 25096 39976
rect 31024 39992 31076 40044
rect 31116 39856 31168 39908
rect 12624 39788 12676 39840
rect 17408 39831 17460 39840
rect 17408 39797 17417 39831
rect 17417 39797 17451 39831
rect 17451 39797 17460 39831
rect 17408 39788 17460 39797
rect 19248 39831 19300 39840
rect 19248 39797 19257 39831
rect 19257 39797 19291 39831
rect 19291 39797 19300 39831
rect 19248 39788 19300 39797
rect 20352 39788 20404 39840
rect 21824 39788 21876 39840
rect 23388 39788 23440 39840
rect 27620 39788 27672 39840
rect 30012 39831 30064 39840
rect 30012 39797 30021 39831
rect 30021 39797 30055 39831
rect 30055 39797 30064 39831
rect 30012 39788 30064 39797
rect 31024 39788 31076 39840
rect 31300 39788 31352 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 5816 39448 5868 39500
rect 11060 39584 11112 39636
rect 11704 39584 11756 39636
rect 15476 39627 15528 39636
rect 15476 39593 15485 39627
rect 15485 39593 15519 39627
rect 15519 39593 15528 39627
rect 15476 39584 15528 39593
rect 21364 39627 21416 39636
rect 21364 39593 21373 39627
rect 21373 39593 21407 39627
rect 21407 39593 21416 39627
rect 21364 39584 21416 39593
rect 32680 39584 32732 39636
rect 1860 39380 1912 39432
rect 6092 39380 6144 39432
rect 9036 39380 9088 39432
rect 9772 39380 9824 39432
rect 12348 39423 12400 39432
rect 12348 39389 12366 39423
rect 12366 39389 12400 39423
rect 12348 39380 12400 39389
rect 12624 39423 12676 39432
rect 12624 39389 12633 39423
rect 12633 39389 12667 39423
rect 12667 39389 12676 39423
rect 12624 39380 12676 39389
rect 13268 39380 13320 39432
rect 16120 39380 16172 39432
rect 18144 39380 18196 39432
rect 19248 39423 19300 39432
rect 19248 39389 19257 39423
rect 19257 39389 19291 39423
rect 19291 39389 19300 39423
rect 19248 39380 19300 39389
rect 19524 39423 19576 39432
rect 19524 39389 19558 39423
rect 19558 39389 19576 39423
rect 19524 39380 19576 39389
rect 21640 39423 21692 39432
rect 21640 39389 21649 39423
rect 21649 39389 21683 39423
rect 21683 39389 21692 39423
rect 21640 39380 21692 39389
rect 5172 39312 5224 39364
rect 16580 39355 16632 39364
rect 16580 39321 16598 39355
rect 16598 39321 16632 39355
rect 16580 39312 16632 39321
rect 21824 39423 21876 39432
rect 21824 39389 21833 39423
rect 21833 39389 21867 39423
rect 21867 39389 21876 39423
rect 21824 39380 21876 39389
rect 22284 39380 22336 39432
rect 25044 39380 25096 39432
rect 27252 39380 27304 39432
rect 31300 39423 31352 39432
rect 31300 39389 31334 39423
rect 31334 39389 31352 39423
rect 31300 39380 31352 39389
rect 21916 39312 21968 39364
rect 23480 39312 23532 39364
rect 27528 39312 27580 39364
rect 30564 39312 30616 39364
rect 31024 39312 31076 39364
rect 6644 39244 6696 39296
rect 10508 39287 10560 39296
rect 10508 39253 10517 39287
rect 10517 39253 10551 39287
rect 10551 39253 10560 39287
rect 10508 39244 10560 39253
rect 20076 39244 20128 39296
rect 22652 39244 22704 39296
rect 28816 39244 28868 39296
rect 29000 39244 29052 39296
rect 30380 39287 30432 39296
rect 30380 39253 30389 39287
rect 30389 39253 30423 39287
rect 30423 39253 30432 39287
rect 30380 39244 30432 39253
rect 31300 39244 31352 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 5172 39083 5224 39092
rect 5172 39049 5181 39083
rect 5181 39049 5215 39083
rect 5215 39049 5224 39083
rect 5172 39040 5224 39049
rect 5264 39040 5316 39092
rect 3053 38947 3105 38956
rect 3053 38913 3080 38947
rect 3080 38913 3105 38947
rect 3053 38904 3105 38913
rect 3148 38947 3200 38956
rect 3148 38913 3162 38947
rect 3162 38913 3196 38947
rect 3196 38913 3200 38947
rect 3332 38947 3384 38956
rect 3148 38904 3200 38913
rect 3332 38913 3341 38947
rect 3341 38913 3375 38947
rect 3375 38913 3384 38947
rect 3332 38904 3384 38913
rect 6000 38972 6052 39024
rect 6092 38972 6144 39024
rect 5816 38947 5868 38956
rect 5816 38913 5825 38947
rect 5825 38913 5859 38947
rect 5859 38913 5868 38947
rect 5816 38904 5868 38913
rect 6644 38904 6696 38956
rect 6736 38947 6788 38956
rect 6736 38913 6745 38947
rect 6745 38913 6779 38947
rect 6779 38913 6788 38947
rect 9036 38972 9088 39024
rect 9680 38972 9732 39024
rect 12440 39040 12492 39092
rect 22100 39040 22152 39092
rect 22744 39040 22796 39092
rect 27160 39083 27212 39092
rect 27160 39049 27169 39083
rect 27169 39049 27203 39083
rect 27203 39049 27212 39083
rect 27160 39040 27212 39049
rect 6736 38904 6788 38913
rect 2872 38768 2924 38820
rect 5264 38768 5316 38820
rect 5448 38768 5500 38820
rect 7656 38836 7708 38888
rect 12532 38904 12584 38956
rect 15568 38904 15620 38956
rect 23020 38972 23072 39024
rect 24952 38972 25004 39024
rect 27896 39040 27948 39092
rect 30840 39040 30892 39092
rect 22652 38947 22704 38956
rect 22652 38913 22661 38947
rect 22661 38913 22695 38947
rect 22695 38913 22704 38947
rect 22652 38904 22704 38913
rect 23296 38904 23348 38956
rect 24584 38904 24636 38956
rect 25412 38947 25464 38956
rect 25412 38913 25421 38947
rect 25421 38913 25455 38947
rect 25455 38913 25464 38947
rect 25412 38904 25464 38913
rect 25596 38947 25648 38956
rect 25596 38913 25605 38947
rect 25605 38913 25639 38947
rect 25639 38913 25648 38947
rect 25596 38904 25648 38913
rect 27620 38947 27672 38956
rect 27620 38913 27629 38947
rect 27629 38913 27663 38947
rect 27663 38913 27672 38947
rect 27620 38904 27672 38913
rect 28080 38904 28132 38956
rect 29000 38904 29052 38956
rect 30380 38904 30432 38956
rect 27712 38836 27764 38888
rect 31024 38904 31076 38956
rect 31576 38904 31628 38956
rect 31760 38904 31812 38956
rect 32772 38904 32824 38956
rect 2688 38743 2740 38752
rect 2688 38709 2697 38743
rect 2697 38709 2731 38743
rect 2731 38709 2740 38743
rect 2688 38700 2740 38709
rect 3332 38700 3384 38752
rect 4804 38700 4856 38752
rect 5816 38700 5868 38752
rect 10324 38743 10376 38752
rect 10324 38709 10333 38743
rect 10333 38709 10367 38743
rect 10367 38709 10376 38743
rect 10324 38700 10376 38709
rect 10968 38700 11020 38752
rect 16304 38768 16356 38820
rect 20628 38768 20680 38820
rect 30840 38768 30892 38820
rect 58164 38811 58216 38820
rect 58164 38777 58173 38811
rect 58173 38777 58207 38811
rect 58207 38777 58216 38811
rect 58164 38768 58216 38777
rect 13820 38700 13872 38752
rect 19432 38700 19484 38752
rect 21640 38700 21692 38752
rect 24768 38743 24820 38752
rect 24768 38709 24777 38743
rect 24777 38709 24811 38743
rect 24811 38709 24820 38743
rect 24768 38700 24820 38709
rect 25228 38700 25280 38752
rect 25596 38700 25648 38752
rect 25964 38700 26016 38752
rect 29092 38700 29144 38752
rect 30472 38743 30524 38752
rect 30472 38709 30481 38743
rect 30481 38709 30515 38743
rect 30515 38709 30524 38743
rect 30472 38700 30524 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 6092 38496 6144 38548
rect 6736 38496 6788 38548
rect 9404 38496 9456 38548
rect 27528 38539 27580 38548
rect 27528 38505 27537 38539
rect 27537 38505 27571 38539
rect 27571 38505 27580 38539
rect 27528 38496 27580 38505
rect 19248 38428 19300 38480
rect 21088 38428 21140 38480
rect 1860 38335 1912 38344
rect 1860 38301 1869 38335
rect 1869 38301 1903 38335
rect 1903 38301 1912 38335
rect 1860 38292 1912 38301
rect 2688 38292 2740 38344
rect 12532 38360 12584 38412
rect 8576 38292 8628 38344
rect 9312 38335 9364 38344
rect 9312 38301 9321 38335
rect 9321 38301 9355 38335
rect 9355 38301 9364 38335
rect 9312 38292 9364 38301
rect 10324 38292 10376 38344
rect 6736 38224 6788 38276
rect 9680 38224 9732 38276
rect 10876 38224 10928 38276
rect 13636 38224 13688 38276
rect 17592 38335 17644 38344
rect 17592 38301 17601 38335
rect 17601 38301 17635 38335
rect 17635 38301 17644 38335
rect 17592 38292 17644 38301
rect 17684 38335 17736 38344
rect 17684 38301 17694 38335
rect 17694 38301 17728 38335
rect 17728 38301 17736 38335
rect 17960 38335 18012 38344
rect 17684 38292 17736 38301
rect 17960 38301 17969 38335
rect 17969 38301 18003 38335
rect 18003 38301 18012 38335
rect 17960 38292 18012 38301
rect 19156 38360 19208 38412
rect 19248 38335 19300 38344
rect 19248 38301 19257 38335
rect 19257 38301 19291 38335
rect 19291 38301 19300 38335
rect 19248 38292 19300 38301
rect 19340 38335 19392 38344
rect 19340 38301 19350 38335
rect 19350 38301 19384 38335
rect 19384 38301 19392 38335
rect 19340 38292 19392 38301
rect 20352 38292 20404 38344
rect 24584 38335 24636 38344
rect 5080 38156 5132 38208
rect 13728 38156 13780 38208
rect 15476 38224 15528 38276
rect 20076 38224 20128 38276
rect 20536 38267 20588 38276
rect 20536 38233 20545 38267
rect 20545 38233 20579 38267
rect 20579 38233 20588 38267
rect 20536 38224 20588 38233
rect 20720 38267 20772 38276
rect 20720 38233 20729 38267
rect 20729 38233 20763 38267
rect 20763 38233 20772 38267
rect 20720 38224 20772 38233
rect 18604 38156 18656 38208
rect 19248 38156 19300 38208
rect 20168 38156 20220 38208
rect 24584 38301 24593 38335
rect 24593 38301 24627 38335
rect 24627 38301 24636 38335
rect 24584 38292 24636 38301
rect 24768 38335 24820 38344
rect 24768 38301 24777 38335
rect 24777 38301 24811 38335
rect 24811 38301 24820 38335
rect 24768 38292 24820 38301
rect 24952 38428 25004 38480
rect 27896 38428 27948 38480
rect 25688 38335 25740 38344
rect 25688 38301 25697 38335
rect 25697 38301 25731 38335
rect 25731 38301 25740 38335
rect 25688 38292 25740 38301
rect 25964 38335 26016 38344
rect 25964 38301 25998 38335
rect 25998 38301 26016 38335
rect 25964 38292 26016 38301
rect 27344 38292 27396 38344
rect 29092 38360 29144 38412
rect 28080 38292 28132 38344
rect 28816 38267 28868 38276
rect 28816 38233 28825 38267
rect 28825 38233 28859 38267
rect 28859 38233 28868 38267
rect 28816 38224 28868 38233
rect 29184 38292 29236 38344
rect 30472 38335 30524 38344
rect 30472 38301 30506 38335
rect 30506 38301 30524 38335
rect 30472 38292 30524 38301
rect 32680 38335 32732 38344
rect 32680 38301 32689 38335
rect 32689 38301 32723 38335
rect 32723 38301 32732 38335
rect 32680 38292 32732 38301
rect 30564 38224 30616 38276
rect 33048 38224 33100 38276
rect 33140 38224 33192 38276
rect 24676 38156 24728 38208
rect 25320 38156 25372 38208
rect 26332 38156 26384 38208
rect 31760 38156 31812 38208
rect 33508 38156 33560 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 3056 37952 3108 38004
rect 3148 37952 3200 38004
rect 11704 37952 11756 38004
rect 4712 37884 4764 37936
rect 17592 37952 17644 38004
rect 17776 37952 17828 38004
rect 20352 37952 20404 38004
rect 25412 37952 25464 38004
rect 29184 37952 29236 38004
rect 31116 37995 31168 38004
rect 31116 37961 31125 37995
rect 31125 37961 31159 37995
rect 31159 37961 31168 37995
rect 31116 37952 31168 37961
rect 13360 37884 13412 37936
rect 13728 37884 13780 37936
rect 16764 37884 16816 37936
rect 19432 37884 19484 37936
rect 2780 37816 2832 37868
rect 3332 37859 3384 37868
rect 3332 37825 3341 37859
rect 3341 37825 3375 37859
rect 3375 37825 3384 37859
rect 3332 37816 3384 37825
rect 3424 37816 3476 37868
rect 5080 37816 5132 37868
rect 9312 37816 9364 37868
rect 11704 37859 11756 37868
rect 11704 37825 11713 37859
rect 11713 37825 11747 37859
rect 11747 37825 11756 37859
rect 11704 37816 11756 37825
rect 12256 37816 12308 37868
rect 10508 37748 10560 37800
rect 18144 37859 18196 37868
rect 12256 37680 12308 37732
rect 13636 37680 13688 37732
rect 18144 37825 18153 37859
rect 18153 37825 18187 37859
rect 18187 37825 18196 37859
rect 18144 37816 18196 37825
rect 18236 37816 18288 37868
rect 19156 37816 19208 37868
rect 19708 37816 19760 37868
rect 20168 37859 20220 37868
rect 20168 37825 20177 37859
rect 20177 37825 20211 37859
rect 20211 37825 20220 37859
rect 20168 37816 20220 37825
rect 23664 37884 23716 37936
rect 25044 37884 25096 37936
rect 25320 37859 25372 37868
rect 25688 37884 25740 37936
rect 26148 37884 26200 37936
rect 32772 37952 32824 38004
rect 33048 37995 33100 38004
rect 33048 37961 33057 37995
rect 33057 37961 33091 37995
rect 33091 37961 33100 37995
rect 33048 37952 33100 37961
rect 25320 37825 25338 37859
rect 25338 37825 25372 37859
rect 25320 37816 25372 37825
rect 26332 37816 26384 37868
rect 29184 37816 29236 37868
rect 31300 37859 31352 37868
rect 31300 37825 31309 37859
rect 31309 37825 31343 37859
rect 31343 37825 31352 37859
rect 31300 37816 31352 37825
rect 31576 37816 31628 37868
rect 32588 37859 32640 37868
rect 32588 37825 32597 37859
rect 32597 37825 32631 37859
rect 32631 37825 32640 37859
rect 32588 37816 32640 37825
rect 20628 37748 20680 37800
rect 22192 37748 22244 37800
rect 27436 37748 27488 37800
rect 29092 37791 29144 37800
rect 29092 37757 29101 37791
rect 29101 37757 29135 37791
rect 29135 37757 29144 37791
rect 29092 37748 29144 37757
rect 33048 37816 33100 37868
rect 33784 37748 33836 37800
rect 20168 37680 20220 37732
rect 2688 37655 2740 37664
rect 2688 37621 2697 37655
rect 2697 37621 2731 37655
rect 2731 37621 2740 37655
rect 2688 37612 2740 37621
rect 6736 37612 6788 37664
rect 11336 37612 11388 37664
rect 13728 37612 13780 37664
rect 17776 37612 17828 37664
rect 19340 37612 19392 37664
rect 20076 37612 20128 37664
rect 20444 37612 20496 37664
rect 20996 37612 21048 37664
rect 24216 37655 24268 37664
rect 24216 37621 24225 37655
rect 24225 37621 24259 37655
rect 24259 37621 24268 37655
rect 24216 37612 24268 37621
rect 27344 37655 27396 37664
rect 27344 37621 27353 37655
rect 27353 37621 27387 37655
rect 27387 37621 27396 37655
rect 27344 37612 27396 37621
rect 30380 37612 30432 37664
rect 33048 37612 33100 37664
rect 34336 37612 34388 37664
rect 58164 37655 58216 37664
rect 58164 37621 58173 37655
rect 58173 37621 58207 37655
rect 58207 37621 58216 37655
rect 58164 37612 58216 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 2780 37408 2832 37460
rect 4068 37408 4120 37460
rect 12348 37408 12400 37460
rect 17408 37408 17460 37460
rect 18236 37408 18288 37460
rect 18512 37451 18564 37460
rect 18512 37417 18521 37451
rect 18521 37417 18555 37451
rect 18555 37417 18564 37451
rect 18512 37408 18564 37417
rect 16856 37340 16908 37392
rect 17684 37340 17736 37392
rect 1860 37315 1912 37324
rect 1860 37281 1869 37315
rect 1869 37281 1903 37315
rect 1903 37281 1912 37315
rect 1860 37272 1912 37281
rect 14648 37272 14700 37324
rect 20536 37408 20588 37460
rect 24768 37408 24820 37460
rect 31484 37408 31536 37460
rect 32588 37408 32640 37460
rect 2688 37204 2740 37256
rect 6092 37204 6144 37256
rect 7104 37136 7156 37188
rect 3332 37068 3384 37120
rect 8116 37247 8168 37256
rect 8116 37213 8125 37247
rect 8125 37213 8159 37247
rect 8159 37213 8168 37247
rect 8116 37204 8168 37213
rect 8208 37247 8260 37256
rect 8208 37213 8217 37247
rect 8217 37213 8251 37247
rect 8251 37213 8260 37247
rect 8208 37204 8260 37213
rect 8024 37179 8076 37188
rect 8024 37145 8033 37179
rect 8033 37145 8067 37179
rect 8067 37145 8076 37179
rect 11704 37204 11756 37256
rect 8024 37136 8076 37145
rect 11336 37179 11388 37188
rect 11336 37145 11345 37179
rect 11345 37145 11379 37179
rect 11379 37145 11388 37179
rect 11336 37136 11388 37145
rect 12348 37136 12400 37188
rect 14372 37179 14424 37188
rect 14372 37145 14381 37179
rect 14381 37145 14415 37179
rect 14415 37145 14424 37179
rect 14372 37136 14424 37145
rect 14556 37179 14608 37188
rect 14556 37145 14565 37179
rect 14565 37145 14599 37179
rect 14599 37145 14608 37179
rect 14556 37136 14608 37145
rect 7564 37068 7616 37120
rect 8944 37068 8996 37120
rect 13268 37111 13320 37120
rect 13268 37077 13277 37111
rect 13277 37077 13311 37111
rect 13311 37077 13320 37111
rect 13268 37068 13320 37077
rect 13728 37068 13780 37120
rect 15200 37136 15252 37188
rect 17408 37247 17460 37256
rect 17408 37213 17417 37247
rect 17417 37213 17451 37247
rect 17451 37213 17460 37247
rect 17592 37247 17644 37256
rect 17408 37204 17460 37213
rect 17592 37213 17601 37247
rect 17601 37213 17635 37247
rect 17635 37213 17644 37247
rect 17592 37204 17644 37213
rect 18512 37204 18564 37256
rect 15568 37179 15620 37188
rect 15568 37145 15602 37179
rect 15602 37145 15620 37179
rect 19340 37247 19392 37256
rect 19340 37213 19350 37247
rect 19350 37213 19384 37247
rect 19384 37213 19392 37247
rect 31576 37272 31628 37324
rect 33324 37272 33376 37324
rect 19340 37204 19392 37213
rect 19708 37247 19760 37256
rect 19708 37213 19722 37247
rect 19722 37213 19756 37247
rect 19756 37213 19760 37247
rect 19708 37204 19760 37213
rect 20996 37204 21048 37256
rect 21824 37247 21876 37256
rect 21824 37213 21833 37247
rect 21833 37213 21867 37247
rect 21867 37213 21876 37247
rect 21824 37204 21876 37213
rect 33416 37204 33468 37256
rect 34244 37272 34296 37324
rect 33692 37247 33744 37256
rect 33692 37213 33701 37247
rect 33701 37213 33735 37247
rect 33735 37213 33744 37247
rect 33692 37204 33744 37213
rect 33784 37247 33836 37256
rect 33784 37213 33793 37247
rect 33793 37213 33827 37247
rect 33827 37213 33836 37247
rect 33784 37204 33836 37213
rect 34336 37204 34388 37256
rect 36728 37204 36780 37256
rect 15568 37136 15620 37145
rect 19432 37136 19484 37188
rect 24216 37136 24268 37188
rect 24952 37136 25004 37188
rect 26148 37136 26200 37188
rect 16120 37068 16172 37120
rect 17408 37068 17460 37120
rect 19156 37068 19208 37120
rect 19708 37068 19760 37120
rect 20904 37068 20956 37120
rect 22836 37068 22888 37120
rect 33508 37068 33560 37120
rect 34520 37068 34572 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 6644 36839 6696 36848
rect 6644 36805 6653 36839
rect 6653 36805 6687 36839
rect 6687 36805 6696 36839
rect 6644 36796 6696 36805
rect 5172 36728 5224 36780
rect 8208 36864 8260 36916
rect 12256 36864 12308 36916
rect 14372 36864 14424 36916
rect 7564 36839 7616 36848
rect 7564 36805 7573 36839
rect 7573 36805 7607 36839
rect 7607 36805 7616 36839
rect 7564 36796 7616 36805
rect 11704 36796 11756 36848
rect 12716 36796 12768 36848
rect 13360 36796 13412 36848
rect 15568 36864 15620 36916
rect 17592 36864 17644 36916
rect 19248 36864 19300 36916
rect 20076 36864 20128 36916
rect 16856 36839 16908 36848
rect 7288 36728 7340 36780
rect 10232 36728 10284 36780
rect 12808 36728 12860 36780
rect 14096 36728 14148 36780
rect 15752 36771 15804 36780
rect 15752 36737 15761 36771
rect 15761 36737 15795 36771
rect 15795 36737 15804 36771
rect 15752 36728 15804 36737
rect 16120 36771 16172 36780
rect 8024 36660 8076 36712
rect 9772 36660 9824 36712
rect 10416 36660 10468 36712
rect 13268 36660 13320 36712
rect 15200 36660 15252 36712
rect 16120 36737 16129 36771
rect 16129 36737 16163 36771
rect 16163 36737 16172 36771
rect 16120 36728 16172 36737
rect 16856 36805 16865 36839
rect 16865 36805 16899 36839
rect 16899 36805 16908 36839
rect 16856 36796 16908 36805
rect 17776 36796 17828 36848
rect 24216 36796 24268 36848
rect 17684 36771 17736 36780
rect 17684 36737 17693 36771
rect 17693 36737 17727 36771
rect 17727 36737 17736 36771
rect 17684 36728 17736 36737
rect 22836 36728 22888 36780
rect 23296 36771 23348 36780
rect 23296 36737 23305 36771
rect 23305 36737 23339 36771
rect 23339 36737 23348 36771
rect 23296 36728 23348 36737
rect 29000 36728 29052 36780
rect 34428 36728 34480 36780
rect 35348 36728 35400 36780
rect 36728 36703 36780 36712
rect 14556 36592 14608 36644
rect 19340 36592 19392 36644
rect 36728 36669 36737 36703
rect 36737 36669 36771 36703
rect 36771 36669 36780 36703
rect 36728 36660 36780 36669
rect 6920 36567 6972 36576
rect 6920 36533 6929 36567
rect 6929 36533 6963 36567
rect 6963 36533 6972 36567
rect 6920 36524 6972 36533
rect 7656 36524 7708 36576
rect 12624 36524 12676 36576
rect 22376 36524 22428 36576
rect 22928 36524 22980 36576
rect 25044 36567 25096 36576
rect 25044 36533 25053 36567
rect 25053 36533 25087 36567
rect 25087 36533 25096 36567
rect 25044 36524 25096 36533
rect 27528 36524 27580 36576
rect 33140 36524 33192 36576
rect 34796 36567 34848 36576
rect 34796 36533 34805 36567
rect 34805 36533 34839 36567
rect 34839 36533 34848 36567
rect 34796 36524 34848 36533
rect 35440 36524 35492 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 5172 36363 5224 36372
rect 5172 36329 5181 36363
rect 5181 36329 5215 36363
rect 5215 36329 5224 36363
rect 5172 36320 5224 36329
rect 7104 36363 7156 36372
rect 7104 36329 7113 36363
rect 7113 36329 7147 36363
rect 7147 36329 7156 36363
rect 7104 36320 7156 36329
rect 14096 36363 14148 36372
rect 14096 36329 14105 36363
rect 14105 36329 14139 36363
rect 14139 36329 14148 36363
rect 14096 36320 14148 36329
rect 15752 36320 15804 36372
rect 16304 36363 16356 36372
rect 16304 36329 16313 36363
rect 16313 36329 16347 36363
rect 16347 36329 16356 36363
rect 16304 36320 16356 36329
rect 29000 36320 29052 36372
rect 29736 36320 29788 36372
rect 1860 36184 1912 36236
rect 7380 36159 7432 36168
rect 7380 36125 7389 36159
rect 7389 36125 7423 36159
rect 7423 36125 7432 36159
rect 7380 36116 7432 36125
rect 8116 36252 8168 36304
rect 27896 36295 27948 36304
rect 27896 36261 27905 36295
rect 27905 36261 27939 36295
rect 27939 36261 27948 36295
rect 27896 36252 27948 36261
rect 28724 36252 28776 36304
rect 7656 36116 7708 36168
rect 9772 36184 9824 36236
rect 12716 36227 12768 36236
rect 12716 36193 12725 36227
rect 12725 36193 12759 36227
rect 12759 36193 12768 36227
rect 12716 36184 12768 36193
rect 8208 36116 8260 36168
rect 4712 36048 4764 36100
rect 10324 36091 10376 36100
rect 10324 36057 10358 36091
rect 10358 36057 10376 36091
rect 10324 36048 10376 36057
rect 10416 36048 10468 36100
rect 12440 36159 12492 36168
rect 12440 36125 12449 36159
rect 12449 36125 12483 36159
rect 12483 36125 12492 36159
rect 12440 36116 12492 36125
rect 14280 36116 14332 36168
rect 21640 36184 21692 36236
rect 22100 36184 22152 36236
rect 13268 36048 13320 36100
rect 14648 36116 14700 36168
rect 14740 36159 14792 36168
rect 14740 36125 14749 36159
rect 14749 36125 14783 36159
rect 14783 36125 14792 36159
rect 22192 36159 22244 36168
rect 14740 36116 14792 36125
rect 22192 36125 22201 36159
rect 22201 36125 22235 36159
rect 22235 36125 22244 36159
rect 22192 36116 22244 36125
rect 24768 36184 24820 36236
rect 28448 36184 28500 36236
rect 22560 36159 22612 36168
rect 22560 36125 22569 36159
rect 22569 36125 22603 36159
rect 22603 36125 22612 36159
rect 22560 36116 22612 36125
rect 22836 36116 22888 36168
rect 15200 36048 15252 36100
rect 22376 36091 22428 36100
rect 22376 36057 22385 36091
rect 22385 36057 22419 36091
rect 22419 36057 22428 36091
rect 22376 36048 22428 36057
rect 27528 36116 27580 36168
rect 29184 36184 29236 36236
rect 28724 36159 28776 36168
rect 28724 36125 28733 36159
rect 28733 36125 28767 36159
rect 28767 36125 28776 36159
rect 28724 36116 28776 36125
rect 30380 36116 30432 36168
rect 33692 36320 33744 36372
rect 35348 36363 35400 36372
rect 35348 36329 35357 36363
rect 35357 36329 35391 36363
rect 35391 36329 35400 36363
rect 35348 36320 35400 36329
rect 33324 36184 33376 36236
rect 34428 36116 34480 36168
rect 34796 36184 34848 36236
rect 34888 36159 34940 36168
rect 34888 36125 34897 36159
rect 34897 36125 34931 36159
rect 34931 36125 34940 36159
rect 34888 36116 34940 36125
rect 33416 36091 33468 36100
rect 33416 36057 33425 36091
rect 33425 36057 33459 36091
rect 33459 36057 33468 36091
rect 33416 36048 33468 36057
rect 34520 36048 34572 36100
rect 9680 35980 9732 36032
rect 11428 36023 11480 36032
rect 11428 35989 11437 36023
rect 11437 35989 11471 36023
rect 11471 35989 11480 36023
rect 11428 35980 11480 35989
rect 21732 35980 21784 36032
rect 22192 35980 22244 36032
rect 22836 35980 22888 36032
rect 23296 35980 23348 36032
rect 27068 36023 27120 36032
rect 27068 35989 27077 36023
rect 27077 35989 27111 36023
rect 27111 35989 27120 36023
rect 27068 35980 27120 35989
rect 29644 35980 29696 36032
rect 34244 35980 34296 36032
rect 36636 36116 36688 36168
rect 58164 36159 58216 36168
rect 58164 36125 58173 36159
rect 58173 36125 58207 36159
rect 58207 36125 58216 36159
rect 58164 36116 58216 36125
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 11428 35776 11480 35828
rect 12256 35776 12308 35828
rect 5172 35708 5224 35760
rect 9680 35708 9732 35760
rect 13728 35776 13780 35828
rect 27068 35776 27120 35828
rect 34888 35776 34940 35828
rect 16120 35708 16172 35760
rect 3608 35640 3660 35692
rect 7288 35640 7340 35692
rect 9864 35683 9916 35692
rect 9864 35649 9873 35683
rect 9873 35649 9907 35683
rect 9907 35649 9916 35683
rect 9864 35640 9916 35649
rect 11796 35640 11848 35692
rect 13176 35640 13228 35692
rect 8208 35572 8260 35624
rect 9220 35572 9272 35624
rect 10968 35615 11020 35624
rect 10968 35581 10977 35615
rect 10977 35581 11011 35615
rect 11011 35581 11020 35615
rect 17132 35640 17184 35692
rect 17408 35683 17460 35692
rect 17408 35649 17417 35683
rect 17417 35649 17451 35683
rect 17451 35649 17460 35683
rect 21824 35708 21876 35760
rect 25044 35708 25096 35760
rect 27804 35708 27856 35760
rect 28448 35708 28500 35760
rect 17408 35640 17460 35649
rect 22192 35640 22244 35692
rect 10968 35572 11020 35581
rect 9496 35504 9548 35556
rect 12624 35504 12676 35556
rect 14740 35504 14792 35556
rect 15200 35504 15252 35556
rect 17132 35504 17184 35556
rect 21180 35504 21232 35556
rect 22836 35683 22888 35692
rect 22836 35649 22845 35683
rect 22845 35649 22879 35683
rect 22879 35649 22888 35683
rect 22836 35640 22888 35649
rect 23388 35640 23440 35692
rect 24216 35683 24268 35692
rect 24216 35649 24225 35683
rect 24225 35649 24259 35683
rect 24259 35649 24268 35683
rect 24216 35640 24268 35649
rect 24308 35640 24360 35692
rect 27436 35640 27488 35692
rect 27620 35683 27672 35692
rect 27620 35649 27654 35683
rect 27654 35649 27672 35683
rect 27620 35640 27672 35649
rect 30288 35683 30340 35692
rect 23296 35572 23348 35624
rect 30288 35649 30297 35683
rect 30297 35649 30331 35683
rect 30331 35649 30340 35683
rect 30288 35640 30340 35649
rect 30656 35708 30708 35760
rect 30472 35683 30524 35692
rect 30472 35649 30481 35683
rect 30481 35649 30515 35683
rect 30515 35649 30524 35683
rect 30472 35640 30524 35649
rect 33416 35640 33468 35692
rect 35348 35640 35400 35692
rect 30932 35572 30984 35624
rect 5172 35479 5224 35488
rect 5172 35445 5181 35479
rect 5181 35445 5215 35479
rect 5215 35445 5224 35479
rect 5172 35436 5224 35445
rect 10784 35436 10836 35488
rect 17224 35436 17276 35488
rect 22468 35479 22520 35488
rect 22468 35445 22477 35479
rect 22477 35445 22511 35479
rect 22511 35445 22520 35479
rect 22468 35436 22520 35445
rect 26424 35436 26476 35488
rect 27528 35436 27580 35488
rect 30472 35504 30524 35556
rect 28448 35436 28500 35488
rect 30748 35479 30800 35488
rect 30748 35445 30757 35479
rect 30757 35445 30791 35479
rect 30791 35445 30800 35479
rect 30748 35436 30800 35445
rect 31484 35479 31536 35488
rect 31484 35445 31493 35479
rect 31493 35445 31527 35479
rect 31527 35445 31536 35479
rect 33324 35572 33376 35624
rect 31484 35436 31536 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4712 35275 4764 35284
rect 4712 35241 4721 35275
rect 4721 35241 4755 35275
rect 4755 35241 4764 35275
rect 4712 35232 4764 35241
rect 11796 35275 11848 35284
rect 2688 35096 2740 35148
rect 11796 35241 11805 35275
rect 11805 35241 11839 35275
rect 11839 35241 11848 35275
rect 11796 35232 11848 35241
rect 17316 35232 17368 35284
rect 8116 35207 8168 35216
rect 8116 35173 8125 35207
rect 8125 35173 8159 35207
rect 8159 35173 8168 35207
rect 8116 35164 8168 35173
rect 5172 35071 5224 35080
rect 5172 35037 5181 35071
rect 5181 35037 5215 35071
rect 5215 35037 5224 35071
rect 5172 35028 5224 35037
rect 5264 34960 5316 35012
rect 2964 34892 3016 34944
rect 6828 35028 6880 35080
rect 9220 35028 9272 35080
rect 9772 35096 9824 35148
rect 10416 35139 10468 35148
rect 10416 35105 10425 35139
rect 10425 35105 10459 35139
rect 10459 35105 10468 35139
rect 10416 35096 10468 35105
rect 9496 35071 9548 35080
rect 9496 35037 9505 35071
rect 9505 35037 9539 35071
rect 9539 35037 9548 35071
rect 9496 35028 9548 35037
rect 7012 34960 7064 35012
rect 10968 35028 11020 35080
rect 13544 35096 13596 35148
rect 17132 35071 17184 35080
rect 9864 34960 9916 35012
rect 12440 34960 12492 35012
rect 7564 34892 7616 34944
rect 12808 34892 12860 34944
rect 17132 35037 17141 35071
rect 17141 35037 17175 35071
rect 17175 35037 17184 35071
rect 17132 35028 17184 35037
rect 17224 35028 17276 35080
rect 20076 35028 20128 35080
rect 24768 35232 24820 35284
rect 25780 35275 25832 35284
rect 25780 35241 25789 35275
rect 25789 35241 25823 35275
rect 25823 35241 25832 35275
rect 25780 35232 25832 35241
rect 27620 35232 27672 35284
rect 20812 35164 20864 35216
rect 18696 34960 18748 35012
rect 20720 34960 20772 35012
rect 22284 35071 22336 35080
rect 22284 35037 22293 35071
rect 22293 35037 22327 35071
rect 22327 35037 22336 35071
rect 22284 35028 22336 35037
rect 22560 35028 22612 35080
rect 27068 35164 27120 35216
rect 24216 35096 24268 35148
rect 27528 35096 27580 35148
rect 27620 35096 27672 35148
rect 26424 35071 26476 35080
rect 26424 35037 26433 35071
rect 26433 35037 26467 35071
rect 26467 35037 26476 35071
rect 26424 35028 26476 35037
rect 27712 35071 27764 35080
rect 27712 35037 27721 35071
rect 27721 35037 27755 35071
rect 27755 35037 27764 35071
rect 27712 35028 27764 35037
rect 33140 35096 33192 35148
rect 22744 34960 22796 35012
rect 23020 34960 23072 35012
rect 24492 34960 24544 35012
rect 28448 35028 28500 35080
rect 30748 35028 30800 35080
rect 32128 35028 32180 35080
rect 32772 35071 32824 35080
rect 32772 35037 32781 35071
rect 32781 35037 32815 35071
rect 32815 35037 32824 35071
rect 32772 35028 32824 35037
rect 58164 35071 58216 35080
rect 58164 35037 58173 35071
rect 58173 35037 58207 35071
rect 58207 35037 58216 35071
rect 58164 35028 58216 35037
rect 29552 34960 29604 35012
rect 18328 34892 18380 34944
rect 18512 34935 18564 34944
rect 18512 34901 18521 34935
rect 18521 34901 18555 34935
rect 18555 34901 18564 34935
rect 18512 34892 18564 34901
rect 19984 34892 20036 34944
rect 21640 34935 21692 34944
rect 21640 34901 21649 34935
rect 21649 34901 21683 34935
rect 21683 34901 21692 34935
rect 21640 34892 21692 34901
rect 21916 34892 21968 34944
rect 23848 34935 23900 34944
rect 23848 34901 23857 34935
rect 23857 34901 23891 34935
rect 23891 34901 23900 34935
rect 23848 34892 23900 34901
rect 24216 34892 24268 34944
rect 24952 34892 25004 34944
rect 25964 34892 26016 34944
rect 26240 34935 26292 34944
rect 26240 34901 26249 34935
rect 26249 34901 26283 34935
rect 26283 34901 26292 34935
rect 26240 34892 26292 34901
rect 29644 34892 29696 34944
rect 30196 34892 30248 34944
rect 31116 34892 31168 34944
rect 34060 34892 34112 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 7012 34731 7064 34740
rect 7012 34697 7021 34731
rect 7021 34697 7055 34731
rect 7055 34697 7064 34731
rect 7012 34688 7064 34697
rect 10324 34731 10376 34740
rect 10324 34697 10333 34731
rect 10333 34697 10367 34731
rect 10367 34697 10376 34731
rect 10324 34688 10376 34697
rect 10416 34688 10468 34740
rect 12624 34688 12676 34740
rect 16672 34688 16724 34740
rect 17408 34688 17460 34740
rect 5448 34620 5500 34672
rect 7196 34620 7248 34672
rect 2780 34595 2832 34604
rect 2780 34561 2814 34595
rect 2814 34561 2832 34595
rect 4712 34595 4764 34604
rect 2780 34552 2832 34561
rect 4712 34561 4721 34595
rect 4721 34561 4755 34595
rect 4755 34561 4764 34595
rect 4712 34552 4764 34561
rect 2412 34484 2464 34536
rect 5540 34527 5592 34536
rect 5540 34493 5549 34527
rect 5549 34493 5583 34527
rect 5583 34493 5592 34527
rect 5540 34484 5592 34493
rect 5724 34484 5776 34536
rect 7196 34484 7248 34536
rect 7472 34595 7524 34604
rect 7472 34561 7481 34595
rect 7481 34561 7515 34595
rect 7515 34561 7524 34595
rect 7472 34552 7524 34561
rect 10508 34620 10560 34672
rect 12900 34620 12952 34672
rect 18512 34620 18564 34672
rect 10600 34595 10652 34604
rect 10600 34561 10609 34595
rect 10609 34561 10643 34595
rect 10643 34561 10652 34595
rect 10600 34552 10652 34561
rect 9864 34484 9916 34536
rect 10784 34595 10836 34604
rect 10784 34561 10793 34595
rect 10793 34561 10827 34595
rect 10827 34561 10836 34595
rect 10784 34552 10836 34561
rect 11152 34552 11204 34604
rect 12256 34595 12308 34604
rect 12256 34561 12265 34595
rect 12265 34561 12299 34595
rect 12299 34561 12308 34595
rect 12256 34552 12308 34561
rect 12440 34595 12492 34604
rect 12440 34561 12449 34595
rect 12449 34561 12483 34595
rect 12483 34561 12492 34595
rect 12440 34552 12492 34561
rect 12808 34552 12860 34604
rect 17684 34595 17736 34604
rect 17684 34561 17693 34595
rect 17693 34561 17727 34595
rect 17727 34561 17736 34595
rect 17684 34552 17736 34561
rect 18328 34552 18380 34604
rect 18972 34620 19024 34672
rect 20076 34688 20128 34740
rect 21640 34620 21692 34672
rect 22744 34688 22796 34740
rect 24492 34731 24544 34740
rect 24492 34697 24501 34731
rect 24501 34697 24535 34731
rect 24535 34697 24544 34731
rect 24492 34688 24544 34697
rect 27068 34731 27120 34740
rect 23112 34620 23164 34672
rect 23664 34620 23716 34672
rect 25780 34663 25832 34672
rect 19156 34484 19208 34536
rect 20720 34552 20772 34604
rect 21824 34595 21876 34604
rect 21824 34561 21833 34595
rect 21833 34561 21867 34595
rect 21867 34561 21876 34595
rect 21824 34552 21876 34561
rect 25780 34629 25789 34663
rect 25789 34629 25823 34663
rect 25823 34629 25832 34663
rect 25780 34620 25832 34629
rect 25964 34663 26016 34672
rect 25964 34629 25973 34663
rect 25973 34629 26007 34663
rect 26007 34629 26016 34663
rect 25964 34620 26016 34629
rect 27068 34697 27077 34731
rect 27077 34697 27111 34731
rect 27111 34697 27120 34731
rect 27068 34688 27120 34697
rect 27712 34688 27764 34740
rect 30288 34688 30340 34740
rect 24860 34595 24912 34604
rect 24860 34561 24869 34595
rect 24869 34561 24903 34595
rect 24903 34561 24912 34595
rect 24860 34552 24912 34561
rect 25136 34595 25188 34604
rect 25136 34561 25145 34595
rect 25145 34561 25179 34595
rect 25179 34561 25188 34595
rect 25136 34552 25188 34561
rect 29552 34595 29604 34604
rect 29552 34561 29561 34595
rect 29561 34561 29595 34595
rect 29595 34561 29604 34595
rect 29552 34552 29604 34561
rect 30196 34620 30248 34672
rect 33048 34620 33100 34672
rect 30932 34595 30984 34604
rect 30932 34561 30941 34595
rect 30941 34561 30975 34595
rect 30975 34561 30984 34595
rect 30932 34552 30984 34561
rect 32128 34595 32180 34604
rect 32128 34561 32137 34595
rect 32137 34561 32171 34595
rect 32171 34561 32180 34595
rect 32128 34552 32180 34561
rect 34796 34688 34848 34740
rect 33416 34552 33468 34604
rect 29644 34484 29696 34536
rect 31484 34484 31536 34536
rect 33324 34484 33376 34536
rect 34244 34416 34296 34468
rect 3148 34348 3200 34400
rect 10600 34348 10652 34400
rect 15936 34348 15988 34400
rect 17224 34348 17276 34400
rect 34060 34348 34112 34400
rect 35900 34484 35952 34536
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2780 34144 2832 34196
rect 4068 34144 4120 34196
rect 5540 34144 5592 34196
rect 7472 34144 7524 34196
rect 10508 34144 10560 34196
rect 19248 34144 19300 34196
rect 20720 34144 20772 34196
rect 24308 34144 24360 34196
rect 24492 34144 24544 34196
rect 2872 33983 2924 33992
rect 2872 33949 2881 33983
rect 2881 33949 2915 33983
rect 2915 33949 2924 33983
rect 2872 33940 2924 33949
rect 3148 33940 3200 33992
rect 4068 33983 4120 33992
rect 4068 33949 4077 33983
rect 4077 33949 4111 33983
rect 4111 33949 4120 33983
rect 4068 33940 4120 33949
rect 4344 33940 4396 33992
rect 7288 34076 7340 34128
rect 7932 34076 7984 34128
rect 5172 33940 5224 33992
rect 5540 33983 5592 33992
rect 5540 33949 5549 33983
rect 5549 33949 5583 33983
rect 5583 33949 5592 33983
rect 5540 33940 5592 33949
rect 7564 34008 7616 34060
rect 8944 33983 8996 33992
rect 8944 33949 8953 33983
rect 8953 33949 8987 33983
rect 8987 33949 8996 33983
rect 8944 33940 8996 33949
rect 9036 33983 9088 33992
rect 9036 33949 9046 33983
rect 9046 33949 9080 33983
rect 9080 33949 9088 33983
rect 15200 34008 15252 34060
rect 9036 33940 9088 33949
rect 13636 33940 13688 33992
rect 13820 33940 13872 33992
rect 15936 33983 15988 33992
rect 15936 33949 15945 33983
rect 15945 33949 15979 33983
rect 15979 33949 15988 33983
rect 15936 33940 15988 33949
rect 5264 33872 5316 33924
rect 7564 33872 7616 33924
rect 9220 33915 9272 33924
rect 9220 33881 9229 33915
rect 9229 33881 9263 33915
rect 9263 33881 9272 33915
rect 9220 33872 9272 33881
rect 15476 33872 15528 33924
rect 16580 33940 16632 33992
rect 17684 33940 17736 33992
rect 19248 33940 19300 33992
rect 19892 33983 19944 33992
rect 19892 33949 19901 33983
rect 19901 33949 19935 33983
rect 19935 33949 19944 33983
rect 19892 33940 19944 33949
rect 19984 33983 20036 33992
rect 19984 33949 19993 33983
rect 19993 33949 20027 33983
rect 20027 33949 20036 33983
rect 19984 33940 20036 33949
rect 20352 33940 20404 33992
rect 24124 33940 24176 33992
rect 24400 33940 24452 33992
rect 24768 33983 24820 33992
rect 24768 33949 24777 33983
rect 24777 33949 24811 33983
rect 24811 33949 24820 33983
rect 24768 33940 24820 33949
rect 26240 34008 26292 34060
rect 27068 34008 27120 34060
rect 16856 33872 16908 33924
rect 18512 33915 18564 33924
rect 18512 33881 18521 33915
rect 18521 33881 18555 33915
rect 18555 33881 18564 33915
rect 18512 33872 18564 33881
rect 23848 33872 23900 33924
rect 25136 33940 25188 33992
rect 26700 33983 26752 33992
rect 26700 33949 26709 33983
rect 26709 33949 26743 33983
rect 26743 33949 26752 33983
rect 26700 33940 26752 33949
rect 27344 33940 27396 33992
rect 27712 33983 27764 33992
rect 27712 33949 27726 33983
rect 27726 33949 27760 33983
rect 27760 33949 27764 33983
rect 27712 33940 27764 33949
rect 30012 33940 30064 33992
rect 30656 33983 30708 33992
rect 30656 33949 30665 33983
rect 30665 33949 30699 33983
rect 30699 33949 30708 33983
rect 30656 33940 30708 33949
rect 30932 33983 30984 33992
rect 30932 33949 30941 33983
rect 30941 33949 30975 33983
rect 30975 33949 30984 33983
rect 30932 33940 30984 33949
rect 33324 33940 33376 33992
rect 33692 33983 33744 33992
rect 33692 33949 33701 33983
rect 33701 33949 33735 33983
rect 33735 33949 33744 33983
rect 33692 33940 33744 33949
rect 36268 34144 36320 34196
rect 29552 33872 29604 33924
rect 31576 33915 31628 33924
rect 31576 33881 31585 33915
rect 31585 33881 31619 33915
rect 31619 33881 31628 33915
rect 31576 33872 31628 33881
rect 33232 33872 33284 33924
rect 34244 33940 34296 33992
rect 34428 33940 34480 33992
rect 36176 33940 36228 33992
rect 36728 33940 36780 33992
rect 37280 33872 37332 33924
rect 3240 33804 3292 33856
rect 3792 33847 3844 33856
rect 3792 33813 3801 33847
rect 3801 33813 3835 33847
rect 3835 33813 3844 33847
rect 3792 33804 3844 33813
rect 5172 33804 5224 33856
rect 8852 33804 8904 33856
rect 11152 33847 11204 33856
rect 11152 33813 11161 33847
rect 11161 33813 11195 33847
rect 11195 33813 11204 33847
rect 11152 33804 11204 33813
rect 15660 33847 15712 33856
rect 15660 33813 15669 33847
rect 15669 33813 15703 33847
rect 15703 33813 15712 33847
rect 15660 33804 15712 33813
rect 16120 33804 16172 33856
rect 27252 33847 27304 33856
rect 27252 33813 27261 33847
rect 27261 33813 27295 33847
rect 27295 33813 27304 33847
rect 27252 33804 27304 33813
rect 27620 33804 27672 33856
rect 30288 33847 30340 33856
rect 30288 33813 30297 33847
rect 30297 33813 30331 33847
rect 30331 33813 30340 33847
rect 30288 33804 30340 33813
rect 33968 33804 34020 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4344 33643 4396 33652
rect 4344 33609 4353 33643
rect 4353 33609 4387 33643
rect 4387 33609 4396 33643
rect 4344 33600 4396 33609
rect 6736 33643 6788 33652
rect 6736 33609 6745 33643
rect 6745 33609 6779 33643
rect 6779 33609 6788 33643
rect 6736 33600 6788 33609
rect 9220 33600 9272 33652
rect 12624 33643 12676 33652
rect 12624 33609 12633 33643
rect 12633 33609 12667 33643
rect 12667 33609 12676 33643
rect 12624 33600 12676 33609
rect 13636 33600 13688 33652
rect 19156 33600 19208 33652
rect 19248 33600 19300 33652
rect 3792 33532 3844 33584
rect 5172 33532 5224 33584
rect 6460 33532 6512 33584
rect 14464 33532 14516 33584
rect 2412 33396 2464 33448
rect 4620 33464 4672 33516
rect 4712 33507 4764 33516
rect 4712 33473 4721 33507
rect 4721 33473 4755 33507
rect 4755 33473 4764 33507
rect 4712 33464 4764 33473
rect 7564 33464 7616 33516
rect 13268 33507 13320 33516
rect 8116 33260 8168 33312
rect 13268 33473 13277 33507
rect 13277 33473 13311 33507
rect 13311 33473 13320 33507
rect 13268 33464 13320 33473
rect 13544 33507 13596 33516
rect 13544 33473 13578 33507
rect 13578 33473 13596 33507
rect 13544 33464 13596 33473
rect 15200 33464 15252 33516
rect 16672 33507 16724 33516
rect 16672 33473 16681 33507
rect 16681 33473 16715 33507
rect 16715 33473 16724 33507
rect 16672 33464 16724 33473
rect 16856 33507 16908 33516
rect 16856 33473 16863 33507
rect 16863 33473 16908 33507
rect 16856 33464 16908 33473
rect 17408 33532 17460 33584
rect 29828 33600 29880 33652
rect 33692 33600 33744 33652
rect 34796 33643 34848 33652
rect 34796 33609 34805 33643
rect 34805 33609 34839 33643
rect 34839 33609 34848 33643
rect 34796 33600 34848 33609
rect 24768 33532 24820 33584
rect 18696 33507 18748 33516
rect 15200 33328 15252 33380
rect 18696 33473 18705 33507
rect 18705 33473 18739 33507
rect 18739 33473 18748 33507
rect 18696 33464 18748 33473
rect 24584 33464 24636 33516
rect 24860 33507 24912 33516
rect 24860 33473 24869 33507
rect 24869 33473 24903 33507
rect 24903 33473 24912 33507
rect 24860 33464 24912 33473
rect 27252 33532 27304 33584
rect 35900 33575 35952 33584
rect 35900 33541 35918 33575
rect 35918 33541 35952 33575
rect 35900 33532 35952 33541
rect 20628 33396 20680 33448
rect 25504 33464 25556 33516
rect 29644 33464 29696 33516
rect 33416 33464 33468 33516
rect 33968 33464 34020 33516
rect 27160 33439 27212 33448
rect 20352 33328 20404 33380
rect 27160 33405 27169 33439
rect 27169 33405 27203 33439
rect 27203 33405 27212 33439
rect 27160 33396 27212 33405
rect 30564 33396 30616 33448
rect 33232 33396 33284 33448
rect 36176 33439 36228 33448
rect 36176 33405 36185 33439
rect 36185 33405 36219 33439
rect 36219 33405 36228 33439
rect 36176 33396 36228 33405
rect 32956 33328 33008 33380
rect 58164 33371 58216 33380
rect 58164 33337 58173 33371
rect 58173 33337 58207 33371
rect 58207 33337 58216 33371
rect 58164 33328 58216 33337
rect 14372 33260 14424 33312
rect 14648 33303 14700 33312
rect 14648 33269 14657 33303
rect 14657 33269 14691 33303
rect 14691 33269 14700 33303
rect 14648 33260 14700 33269
rect 17316 33303 17368 33312
rect 17316 33269 17325 33303
rect 17325 33269 17359 33303
rect 17359 33269 17368 33303
rect 17316 33260 17368 33269
rect 18236 33260 18288 33312
rect 19248 33303 19300 33312
rect 19248 33269 19257 33303
rect 19257 33269 19291 33303
rect 19291 33269 19300 33303
rect 19248 33260 19300 33269
rect 23848 33260 23900 33312
rect 25320 33303 25372 33312
rect 25320 33269 25329 33303
rect 25329 33269 25363 33303
rect 25363 33269 25372 33303
rect 25320 33260 25372 33269
rect 25504 33260 25556 33312
rect 28540 33303 28592 33312
rect 28540 33269 28549 33303
rect 28549 33269 28583 33303
rect 28583 33269 28592 33303
rect 28540 33260 28592 33269
rect 29644 33260 29696 33312
rect 30932 33260 30984 33312
rect 35992 33260 36044 33312
rect 37280 33303 37332 33312
rect 37280 33269 37289 33303
rect 37289 33269 37323 33303
rect 37323 33269 37332 33303
rect 37280 33260 37332 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 5172 33056 5224 33108
rect 5264 33056 5316 33108
rect 7196 33056 7248 33108
rect 6736 32852 6788 32904
rect 8116 32920 8168 32972
rect 7380 32895 7432 32904
rect 7380 32861 7389 32895
rect 7389 32861 7423 32895
rect 7423 32861 7432 32895
rect 7380 32852 7432 32861
rect 6828 32784 6880 32836
rect 7656 32852 7708 32904
rect 9956 33056 10008 33108
rect 10416 33056 10468 33108
rect 13544 33099 13596 33108
rect 13544 33065 13553 33099
rect 13553 33065 13587 33099
rect 13587 33065 13596 33099
rect 13544 33056 13596 33065
rect 12716 32988 12768 33040
rect 10416 32920 10468 32972
rect 10232 32895 10284 32904
rect 10232 32861 10241 32895
rect 10241 32861 10275 32895
rect 10275 32861 10284 32895
rect 10232 32852 10284 32861
rect 10876 32852 10928 32904
rect 12716 32852 12768 32904
rect 13084 32895 13136 32904
rect 13084 32861 13093 32895
rect 13093 32861 13127 32895
rect 13127 32861 13136 32895
rect 13084 32852 13136 32861
rect 13820 32920 13872 32972
rect 14096 32895 14148 32904
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 16580 33056 16632 33108
rect 16856 33056 16908 33108
rect 19248 33056 19300 33108
rect 25228 33056 25280 33108
rect 25780 33056 25832 33108
rect 27712 33056 27764 33108
rect 31024 33056 31076 33108
rect 31576 33056 31628 33108
rect 15476 32920 15528 32972
rect 16672 32920 16724 32972
rect 14740 32852 14792 32904
rect 17132 32852 17184 32904
rect 17960 32852 18012 32904
rect 18144 32920 18196 32972
rect 20628 33031 20680 33040
rect 20628 32997 20637 33031
rect 20637 32997 20671 33031
rect 20671 32997 20680 33031
rect 20628 32988 20680 32997
rect 18236 32895 18288 32904
rect 18236 32861 18245 32895
rect 18245 32861 18279 32895
rect 18279 32861 18288 32895
rect 18236 32852 18288 32861
rect 24584 32920 24636 32972
rect 19248 32895 19300 32904
rect 15660 32784 15712 32836
rect 7196 32716 7248 32768
rect 7472 32716 7524 32768
rect 10140 32716 10192 32768
rect 12900 32716 12952 32768
rect 17040 32716 17092 32768
rect 19248 32861 19257 32895
rect 19257 32861 19291 32895
rect 19291 32861 19300 32895
rect 19248 32852 19300 32861
rect 28540 32852 28592 32904
rect 33140 32852 33192 32904
rect 29552 32784 29604 32836
rect 29920 32784 29972 32836
rect 30288 32784 30340 32836
rect 32128 32827 32180 32836
rect 32128 32793 32137 32827
rect 32137 32793 32171 32827
rect 32171 32793 32180 32827
rect 32128 32784 32180 32793
rect 33232 32784 33284 32836
rect 19984 32716 20036 32768
rect 21916 32716 21968 32768
rect 24032 32716 24084 32768
rect 32404 32716 32456 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 4896 32512 4948 32564
rect 5356 32512 5408 32564
rect 6460 32555 6512 32564
rect 6460 32521 6469 32555
rect 6469 32521 6503 32555
rect 6503 32521 6512 32555
rect 6460 32512 6512 32521
rect 6736 32512 6788 32564
rect 7656 32512 7708 32564
rect 6000 32444 6052 32496
rect 9128 32512 9180 32564
rect 7196 32419 7248 32428
rect 7196 32385 7230 32419
rect 7230 32385 7248 32419
rect 7196 32376 7248 32385
rect 6828 32308 6880 32360
rect 9036 32444 9088 32496
rect 11888 32444 11940 32496
rect 13084 32512 13136 32564
rect 14648 32444 14700 32496
rect 17040 32487 17092 32496
rect 17040 32453 17049 32487
rect 17049 32453 17083 32487
rect 17083 32453 17092 32487
rect 17040 32444 17092 32453
rect 9680 32376 9732 32428
rect 12532 32376 12584 32428
rect 13268 32376 13320 32428
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 16856 32419 16908 32428
rect 16856 32385 16865 32419
rect 16865 32385 16899 32419
rect 16899 32385 16908 32419
rect 16856 32376 16908 32385
rect 7564 32172 7616 32224
rect 13452 32308 13504 32360
rect 12072 32240 12124 32292
rect 17132 32308 17184 32360
rect 18144 32512 18196 32564
rect 21180 32555 21232 32564
rect 21180 32521 21189 32555
rect 21189 32521 21223 32555
rect 21223 32521 21232 32555
rect 21180 32512 21232 32521
rect 21640 32512 21692 32564
rect 22100 32555 22152 32564
rect 22100 32521 22109 32555
rect 22109 32521 22143 32555
rect 22143 32521 22152 32555
rect 22100 32512 22152 32521
rect 24860 32512 24912 32564
rect 18512 32444 18564 32496
rect 18696 32376 18748 32428
rect 21916 32419 21968 32428
rect 21916 32385 21925 32419
rect 21925 32385 21959 32419
rect 21959 32385 21968 32419
rect 21916 32376 21968 32385
rect 22836 32376 22888 32428
rect 23756 32444 23808 32496
rect 25412 32512 25464 32564
rect 28816 32512 28868 32564
rect 29736 32555 29788 32564
rect 25320 32444 25372 32496
rect 28448 32444 28500 32496
rect 28540 32444 28592 32496
rect 24032 32376 24084 32428
rect 24216 32376 24268 32428
rect 20812 32308 20864 32360
rect 27160 32308 27212 32360
rect 21364 32240 21416 32292
rect 23848 32240 23900 32292
rect 13636 32172 13688 32224
rect 25044 32172 25096 32224
rect 28172 32376 28224 32428
rect 29736 32521 29745 32555
rect 29745 32521 29779 32555
rect 29779 32521 29788 32555
rect 29736 32512 29788 32521
rect 30564 32487 30616 32496
rect 30564 32453 30573 32487
rect 30573 32453 30607 32487
rect 30607 32453 30616 32487
rect 30564 32444 30616 32453
rect 30748 32444 30800 32496
rect 33048 32444 33100 32496
rect 29000 32308 29052 32360
rect 32864 32376 32916 32428
rect 36176 32376 36228 32428
rect 37464 32419 37516 32428
rect 37464 32385 37473 32419
rect 37473 32385 37507 32419
rect 37507 32385 37516 32419
rect 37464 32376 37516 32385
rect 37556 32376 37608 32428
rect 30564 32240 30616 32292
rect 29000 32172 29052 32224
rect 30104 32172 30156 32224
rect 30472 32215 30524 32224
rect 30472 32181 30481 32215
rect 30481 32181 30515 32215
rect 30515 32181 30524 32215
rect 30472 32172 30524 32181
rect 30840 32172 30892 32224
rect 33232 32172 33284 32224
rect 33784 32172 33836 32224
rect 35900 32215 35952 32224
rect 35900 32181 35909 32215
rect 35909 32181 35943 32215
rect 35943 32181 35952 32215
rect 35900 32172 35952 32181
rect 38660 32172 38712 32224
rect 58164 32215 58216 32224
rect 58164 32181 58173 32215
rect 58173 32181 58207 32215
rect 58207 32181 58216 32215
rect 58164 32172 58216 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2412 31764 2464 31816
rect 6736 31968 6788 32020
rect 13452 31968 13504 32020
rect 16028 31968 16080 32020
rect 17132 31968 17184 32020
rect 22836 31968 22888 32020
rect 23664 32011 23716 32020
rect 5264 31900 5316 31952
rect 6184 31900 6236 31952
rect 6828 31900 6880 31952
rect 11888 31943 11940 31952
rect 5172 31807 5224 31816
rect 5172 31773 5181 31807
rect 5181 31773 5215 31807
rect 5215 31773 5224 31807
rect 5172 31764 5224 31773
rect 5356 31807 5408 31816
rect 5356 31773 5365 31807
rect 5365 31773 5399 31807
rect 5399 31773 5408 31807
rect 5356 31764 5408 31773
rect 6000 31764 6052 31816
rect 7196 31832 7248 31884
rect 7288 31832 7340 31884
rect 11888 31909 11897 31943
rect 11897 31909 11931 31943
rect 11931 31909 11940 31943
rect 11888 31900 11940 31909
rect 22560 31900 22612 31952
rect 6736 31764 6788 31816
rect 8484 31764 8536 31816
rect 9864 31807 9916 31816
rect 9864 31773 9898 31807
rect 9898 31773 9916 31807
rect 9864 31764 9916 31773
rect 11520 31764 11572 31816
rect 14740 31764 14792 31816
rect 18788 31764 18840 31816
rect 22652 31832 22704 31884
rect 22836 31832 22888 31884
rect 23664 31977 23673 32011
rect 23673 31977 23707 32011
rect 23707 31977 23716 32011
rect 23664 31968 23716 31977
rect 23848 31968 23900 32020
rect 24124 31968 24176 32020
rect 29920 31968 29972 32020
rect 32864 32011 32916 32020
rect 32864 31977 32873 32011
rect 32873 31977 32907 32011
rect 32907 31977 32916 32011
rect 32864 31968 32916 31977
rect 37556 31968 37608 32020
rect 31668 31900 31720 31952
rect 27160 31875 27212 31884
rect 27160 31841 27169 31875
rect 27169 31841 27203 31875
rect 27203 31841 27212 31875
rect 27160 31832 27212 31841
rect 30288 31832 30340 31884
rect 2136 31739 2188 31748
rect 2136 31705 2170 31739
rect 2170 31705 2188 31739
rect 2136 31696 2188 31705
rect 12348 31696 12400 31748
rect 12992 31739 13044 31748
rect 12992 31705 13010 31739
rect 13010 31705 13044 31739
rect 12992 31696 13044 31705
rect 29736 31764 29788 31816
rect 30748 31764 30800 31816
rect 30932 31807 30984 31816
rect 30932 31773 30941 31807
rect 30941 31773 30975 31807
rect 30975 31773 30984 31807
rect 30932 31764 30984 31773
rect 31024 31807 31076 31816
rect 31024 31773 31033 31807
rect 31033 31773 31067 31807
rect 31067 31773 31076 31807
rect 31300 31807 31352 31816
rect 31024 31764 31076 31773
rect 31300 31773 31309 31807
rect 31309 31773 31343 31807
rect 31343 31773 31352 31807
rect 31300 31764 31352 31773
rect 33324 31900 33376 31952
rect 35900 31900 35952 31952
rect 32404 31807 32456 31816
rect 32404 31773 32413 31807
rect 32413 31773 32447 31807
rect 32447 31773 32456 31807
rect 32404 31764 32456 31773
rect 32956 31832 33008 31884
rect 36084 31832 36136 31884
rect 32864 31764 32916 31816
rect 35440 31764 35492 31816
rect 35992 31807 36044 31816
rect 35992 31773 36001 31807
rect 36001 31773 36035 31807
rect 36035 31773 36044 31807
rect 35992 31764 36044 31773
rect 36176 31807 36228 31816
rect 36176 31773 36185 31807
rect 36185 31773 36219 31807
rect 36219 31773 36228 31807
rect 36176 31764 36228 31773
rect 28080 31696 28132 31748
rect 31208 31696 31260 31748
rect 35164 31739 35216 31748
rect 35164 31705 35173 31739
rect 35173 31705 35207 31739
rect 35207 31705 35216 31739
rect 35164 31696 35216 31705
rect 3424 31628 3476 31680
rect 5632 31671 5684 31680
rect 5632 31637 5641 31671
rect 5641 31637 5675 31671
rect 5675 31637 5684 31671
rect 5632 31628 5684 31637
rect 6184 31671 6236 31680
rect 6184 31637 6193 31671
rect 6193 31637 6227 31671
rect 6227 31637 6236 31671
rect 6184 31628 6236 31637
rect 10968 31671 11020 31680
rect 10968 31637 10977 31671
rect 10977 31637 11011 31671
rect 11011 31637 11020 31671
rect 10968 31628 11020 31637
rect 13360 31628 13412 31680
rect 15016 31628 15068 31680
rect 17960 31628 18012 31680
rect 24676 31628 24728 31680
rect 34060 31628 34112 31680
rect 36360 31628 36412 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 2136 31467 2188 31476
rect 2136 31433 2145 31467
rect 2145 31433 2179 31467
rect 2179 31433 2188 31467
rect 2136 31424 2188 31433
rect 5172 31424 5224 31476
rect 2688 31356 2740 31408
rect 6736 31424 6788 31476
rect 12992 31424 13044 31476
rect 6184 31356 6236 31408
rect 11888 31356 11940 31408
rect 12900 31356 12952 31408
rect 18328 31424 18380 31476
rect 24216 31467 24268 31476
rect 24216 31433 24225 31467
rect 24225 31433 24259 31467
rect 24259 31433 24268 31467
rect 24216 31424 24268 31433
rect 15844 31399 15896 31408
rect 15844 31365 15853 31399
rect 15853 31365 15887 31399
rect 15887 31365 15896 31399
rect 15844 31356 15896 31365
rect 16028 31399 16080 31408
rect 16028 31365 16037 31399
rect 16037 31365 16071 31399
rect 16071 31365 16080 31399
rect 16028 31356 16080 31365
rect 23020 31399 23072 31408
rect 23020 31365 23029 31399
rect 23029 31365 23063 31399
rect 23063 31365 23072 31399
rect 23020 31356 23072 31365
rect 32772 31424 32824 31476
rect 36176 31424 36228 31476
rect 2872 31288 2924 31340
rect 3424 31331 3476 31340
rect 3424 31297 3433 31331
rect 3433 31297 3467 31331
rect 3467 31297 3476 31331
rect 3424 31288 3476 31297
rect 3608 31331 3660 31340
rect 3608 31297 3617 31331
rect 3617 31297 3651 31331
rect 3651 31297 3660 31331
rect 3608 31288 3660 31297
rect 7564 31288 7616 31340
rect 8208 31288 8260 31340
rect 10968 31288 11020 31340
rect 6368 31263 6420 31272
rect 6368 31229 6377 31263
rect 6377 31229 6411 31263
rect 6411 31229 6420 31263
rect 6368 31220 6420 31229
rect 9680 31263 9732 31272
rect 9680 31229 9689 31263
rect 9689 31229 9723 31263
rect 9723 31229 9732 31263
rect 9680 31220 9732 31229
rect 11980 31220 12032 31272
rect 2780 31152 2832 31204
rect 7288 31084 7340 31136
rect 8392 31084 8444 31136
rect 9128 31084 9180 31136
rect 10324 31084 10376 31136
rect 12624 31288 12676 31340
rect 13360 31331 13412 31340
rect 13360 31297 13369 31331
rect 13369 31297 13403 31331
rect 13403 31297 13412 31331
rect 13360 31288 13412 31297
rect 12992 31220 13044 31272
rect 13636 31288 13688 31340
rect 13728 31331 13780 31340
rect 13728 31297 13737 31331
rect 13737 31297 13771 31331
rect 13771 31297 13780 31331
rect 13728 31288 13780 31297
rect 12440 31084 12492 31136
rect 14648 31331 14700 31340
rect 14648 31297 14658 31331
rect 14658 31297 14692 31331
rect 14692 31297 14700 31331
rect 14648 31288 14700 31297
rect 14832 31331 14884 31340
rect 14832 31297 14841 31331
rect 14841 31297 14875 31331
rect 14875 31297 14884 31331
rect 14832 31288 14884 31297
rect 15200 31288 15252 31340
rect 19984 31288 20036 31340
rect 21640 31288 21692 31340
rect 22560 31331 22612 31340
rect 14372 31220 14424 31272
rect 15476 31152 15528 31204
rect 21180 31220 21232 31272
rect 21824 31220 21876 31272
rect 22560 31297 22569 31331
rect 22569 31297 22603 31331
rect 22603 31297 22612 31331
rect 22560 31288 22612 31297
rect 23204 31331 23256 31340
rect 23204 31297 23213 31331
rect 23213 31297 23247 31331
rect 23247 31297 23256 31331
rect 23204 31288 23256 31297
rect 23664 31288 23716 31340
rect 29460 31356 29512 31408
rect 30288 31399 30340 31408
rect 30288 31365 30297 31399
rect 30297 31365 30331 31399
rect 30331 31365 30340 31399
rect 30288 31356 30340 31365
rect 31116 31399 31168 31408
rect 31116 31365 31125 31399
rect 31125 31365 31159 31399
rect 31159 31365 31168 31399
rect 31116 31356 31168 31365
rect 31208 31399 31260 31408
rect 31208 31365 31217 31399
rect 31217 31365 31251 31399
rect 31251 31365 31260 31399
rect 31208 31356 31260 31365
rect 35164 31356 35216 31408
rect 35532 31356 35584 31408
rect 30932 31288 30984 31340
rect 31760 31288 31812 31340
rect 35992 31356 36044 31408
rect 36084 31331 36136 31340
rect 15292 31084 15344 31136
rect 19156 31127 19208 31136
rect 19156 31093 19165 31127
rect 19165 31093 19199 31127
rect 19199 31093 19208 31127
rect 19156 31084 19208 31093
rect 19984 31084 20036 31136
rect 21916 31127 21968 31136
rect 21916 31093 21925 31127
rect 21925 31093 21959 31127
rect 21959 31093 21968 31127
rect 21916 31084 21968 31093
rect 22284 31152 22336 31204
rect 33140 31220 33192 31272
rect 33232 31220 33284 31272
rect 36084 31297 36093 31331
rect 36093 31297 36127 31331
rect 36127 31297 36136 31331
rect 36084 31288 36136 31297
rect 36360 31356 36412 31408
rect 36268 31331 36320 31340
rect 36268 31297 36277 31331
rect 36277 31297 36311 31331
rect 36311 31297 36320 31331
rect 36268 31288 36320 31297
rect 37464 31288 37516 31340
rect 37924 31288 37976 31340
rect 38660 31288 38712 31340
rect 23020 31084 23072 31136
rect 24860 31084 24912 31136
rect 25688 31084 25740 31136
rect 28724 31084 28776 31136
rect 31024 31084 31076 31136
rect 32864 31084 32916 31136
rect 35440 31084 35492 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2412 30744 2464 30796
rect 6368 30880 6420 30932
rect 7196 30923 7248 30932
rect 7196 30889 7205 30923
rect 7205 30889 7239 30923
rect 7239 30889 7248 30923
rect 7196 30880 7248 30889
rect 11520 30880 11572 30932
rect 5632 30719 5684 30728
rect 5632 30685 5666 30719
rect 5666 30685 5684 30719
rect 5632 30676 5684 30685
rect 7564 30719 7616 30728
rect 7564 30685 7573 30719
rect 7573 30685 7607 30719
rect 7607 30685 7616 30719
rect 7564 30676 7616 30685
rect 13728 30812 13780 30864
rect 15844 30812 15896 30864
rect 14740 30787 14792 30796
rect 14740 30753 14749 30787
rect 14749 30753 14783 30787
rect 14783 30753 14792 30787
rect 14740 30744 14792 30753
rect 17960 30744 18012 30796
rect 19248 30787 19300 30796
rect 19248 30753 19257 30787
rect 19257 30753 19291 30787
rect 19291 30753 19300 30787
rect 19248 30744 19300 30753
rect 23204 30880 23256 30932
rect 23848 30880 23900 30932
rect 27896 30880 27948 30932
rect 34060 30880 34112 30932
rect 30564 30812 30616 30864
rect 18328 30719 18380 30728
rect 18328 30685 18337 30719
rect 18337 30685 18371 30719
rect 18371 30685 18380 30719
rect 18328 30676 18380 30685
rect 7288 30608 7340 30660
rect 14740 30608 14792 30660
rect 18512 30719 18564 30728
rect 18512 30685 18521 30719
rect 18521 30685 18555 30719
rect 18555 30685 18564 30719
rect 18512 30676 18564 30685
rect 18880 30676 18932 30728
rect 21548 30719 21600 30728
rect 21548 30685 21557 30719
rect 21557 30685 21591 30719
rect 21591 30685 21600 30719
rect 21548 30676 21600 30685
rect 24768 30744 24820 30796
rect 22284 30676 22336 30728
rect 24400 30719 24452 30728
rect 2780 30540 2832 30592
rect 6736 30583 6788 30592
rect 6736 30549 6745 30583
rect 6745 30549 6779 30583
rect 6779 30549 6788 30583
rect 6736 30540 6788 30549
rect 16948 30540 17000 30592
rect 18052 30583 18104 30592
rect 18052 30549 18061 30583
rect 18061 30549 18095 30583
rect 18095 30549 18104 30583
rect 18052 30540 18104 30549
rect 19432 30540 19484 30592
rect 21916 30608 21968 30660
rect 24400 30685 24409 30719
rect 24409 30685 24443 30719
rect 24443 30685 24452 30719
rect 24400 30676 24452 30685
rect 27068 30719 27120 30728
rect 27068 30685 27077 30719
rect 27077 30685 27111 30719
rect 27111 30685 27120 30719
rect 27068 30676 27120 30685
rect 27896 30676 27948 30728
rect 30472 30744 30524 30796
rect 30656 30787 30708 30796
rect 30656 30753 30665 30787
rect 30665 30753 30699 30787
rect 30699 30753 30708 30787
rect 30656 30744 30708 30753
rect 28724 30719 28776 30728
rect 28724 30685 28733 30719
rect 28733 30685 28767 30719
rect 28767 30685 28776 30719
rect 28724 30676 28776 30685
rect 29000 30676 29052 30728
rect 31392 30719 31444 30728
rect 24860 30608 24912 30660
rect 26240 30608 26292 30660
rect 31392 30685 31401 30719
rect 31401 30685 31435 30719
rect 31435 30685 31444 30719
rect 31392 30676 31444 30685
rect 33140 30719 33192 30728
rect 33140 30685 33149 30719
rect 33149 30685 33183 30719
rect 33183 30685 33192 30719
rect 33140 30676 33192 30685
rect 33232 30719 33284 30728
rect 33232 30685 33241 30719
rect 33241 30685 33275 30719
rect 33275 30685 33284 30719
rect 33508 30719 33560 30728
rect 33232 30676 33284 30685
rect 33508 30685 33517 30719
rect 33517 30685 33551 30719
rect 33551 30685 33560 30719
rect 33508 30676 33560 30685
rect 31852 30608 31904 30660
rect 32588 30608 32640 30660
rect 33416 30608 33468 30660
rect 33876 30608 33928 30660
rect 35992 30812 36044 30864
rect 35992 30719 36044 30728
rect 35992 30685 36001 30719
rect 36001 30685 36035 30719
rect 36035 30685 36044 30719
rect 35992 30676 36044 30685
rect 36360 30744 36412 30796
rect 37924 30787 37976 30796
rect 37924 30753 37933 30787
rect 37933 30753 37967 30787
rect 37967 30753 37976 30787
rect 37924 30744 37976 30753
rect 58164 30719 58216 30728
rect 58164 30685 58173 30719
rect 58173 30685 58207 30719
rect 58207 30685 58216 30719
rect 58164 30676 58216 30685
rect 20076 30540 20128 30592
rect 22100 30540 22152 30592
rect 23848 30540 23900 30592
rect 25136 30540 25188 30592
rect 28356 30540 28408 30592
rect 32128 30540 32180 30592
rect 32312 30540 32364 30592
rect 32956 30583 33008 30592
rect 32956 30549 32965 30583
rect 32965 30549 32999 30583
rect 32999 30549 33008 30583
rect 32956 30540 33008 30549
rect 37372 30540 37424 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 8484 30336 8536 30388
rect 14740 30379 14792 30388
rect 9864 30311 9916 30320
rect 9864 30277 9873 30311
rect 9873 30277 9907 30311
rect 9907 30277 9916 30311
rect 9864 30268 9916 30277
rect 2412 30243 2464 30252
rect 2412 30209 2421 30243
rect 2421 30209 2455 30243
rect 2455 30209 2464 30243
rect 2412 30200 2464 30209
rect 2504 30200 2556 30252
rect 11704 30268 11756 30320
rect 11980 30268 12032 30320
rect 14740 30345 14749 30379
rect 14749 30345 14783 30379
rect 14783 30345 14792 30379
rect 14740 30336 14792 30345
rect 15200 30336 15252 30388
rect 14648 30268 14700 30320
rect 9312 30132 9364 30184
rect 10324 30243 10376 30252
rect 10324 30209 10333 30243
rect 10333 30209 10367 30243
rect 10367 30209 10376 30243
rect 10324 30200 10376 30209
rect 10968 30200 11020 30252
rect 14832 30200 14884 30252
rect 15016 30243 15068 30252
rect 15016 30209 15025 30243
rect 15025 30209 15059 30243
rect 15059 30209 15068 30243
rect 15016 30200 15068 30209
rect 16856 30268 16908 30320
rect 15292 30200 15344 30252
rect 15384 30243 15436 30252
rect 15384 30209 15393 30243
rect 15393 30209 15427 30243
rect 15427 30209 15436 30243
rect 15384 30200 15436 30209
rect 16672 30200 16724 30252
rect 19432 30336 19484 30388
rect 29460 30379 29512 30388
rect 29460 30345 29469 30379
rect 29469 30345 29503 30379
rect 29503 30345 29512 30379
rect 29460 30336 29512 30345
rect 18052 30268 18104 30320
rect 18880 30268 18932 30320
rect 21180 30311 21232 30320
rect 19248 30200 19300 30252
rect 11060 30132 11112 30184
rect 15844 30132 15896 30184
rect 16580 30132 16632 30184
rect 17960 30175 18012 30184
rect 17960 30141 17969 30175
rect 17969 30141 18003 30175
rect 18003 30141 18012 30175
rect 17960 30132 18012 30141
rect 20260 30243 20312 30252
rect 20260 30209 20269 30243
rect 20269 30209 20303 30243
rect 20303 30209 20312 30243
rect 21180 30277 21189 30311
rect 21189 30277 21223 30311
rect 21223 30277 21232 30311
rect 21180 30268 21232 30277
rect 23756 30268 23808 30320
rect 20260 30200 20312 30209
rect 20352 30132 20404 30184
rect 22192 30200 22244 30252
rect 22560 30243 22612 30252
rect 22560 30209 22569 30243
rect 22569 30209 22603 30243
rect 22603 30209 22612 30243
rect 22560 30200 22612 30209
rect 23204 30200 23256 30252
rect 23664 30243 23716 30252
rect 23664 30209 23673 30243
rect 23673 30209 23707 30243
rect 23707 30209 23716 30243
rect 23664 30200 23716 30209
rect 23480 30132 23532 30184
rect 25136 30268 25188 30320
rect 26240 30268 26292 30320
rect 24216 30200 24268 30252
rect 24584 30243 24636 30252
rect 24584 30209 24593 30243
rect 24593 30209 24627 30243
rect 24627 30209 24636 30243
rect 24584 30200 24636 30209
rect 25688 30243 25740 30252
rect 3700 29996 3752 30048
rect 9312 29996 9364 30048
rect 24400 30064 24452 30116
rect 25688 30209 25697 30243
rect 25697 30209 25731 30243
rect 25731 30209 25740 30243
rect 29920 30268 29972 30320
rect 30380 30268 30432 30320
rect 25688 30200 25740 30209
rect 27068 30200 27120 30252
rect 28356 30243 28408 30252
rect 28356 30209 28390 30243
rect 28390 30209 28408 30243
rect 28356 30200 28408 30209
rect 30104 30243 30156 30252
rect 30104 30209 30113 30243
rect 30113 30209 30147 30243
rect 30147 30209 30156 30243
rect 30104 30200 30156 30209
rect 31208 30268 31260 30320
rect 32588 30311 32640 30320
rect 32588 30277 32597 30311
rect 32597 30277 32631 30311
rect 32631 30277 32640 30311
rect 32588 30268 32640 30277
rect 33692 30311 33744 30320
rect 33692 30277 33701 30311
rect 33701 30277 33735 30311
rect 33735 30277 33744 30311
rect 33692 30268 33744 30277
rect 35992 30336 36044 30388
rect 37372 30268 37424 30320
rect 24952 30064 25004 30116
rect 11704 29996 11756 30048
rect 12900 29996 12952 30048
rect 13176 29996 13228 30048
rect 15016 29996 15068 30048
rect 15936 30039 15988 30048
rect 15936 30005 15945 30039
rect 15945 30005 15979 30039
rect 15979 30005 15988 30039
rect 15936 29996 15988 30005
rect 17132 30039 17184 30048
rect 17132 30005 17141 30039
rect 17141 30005 17175 30039
rect 17175 30005 17184 30039
rect 17132 29996 17184 30005
rect 19340 30039 19392 30048
rect 19340 30005 19349 30039
rect 19349 30005 19383 30039
rect 19383 30005 19392 30039
rect 19340 29996 19392 30005
rect 22376 29996 22428 30048
rect 25872 30039 25924 30048
rect 25872 30005 25881 30039
rect 25881 30005 25915 30039
rect 25915 30005 25924 30039
rect 25872 29996 25924 30005
rect 30564 30132 30616 30184
rect 33140 30200 33192 30252
rect 33508 30200 33560 30252
rect 33876 30200 33928 30252
rect 34060 30200 34112 30252
rect 35532 30243 35584 30252
rect 35532 30209 35541 30243
rect 35541 30209 35575 30243
rect 35575 30209 35584 30243
rect 35532 30200 35584 30209
rect 34796 30132 34848 30184
rect 32864 30064 32916 30116
rect 33692 30064 33744 30116
rect 35440 30064 35492 30116
rect 29276 29996 29328 30048
rect 30656 29996 30708 30048
rect 31392 29996 31444 30048
rect 33324 29996 33376 30048
rect 33876 29996 33928 30048
rect 36636 30039 36688 30048
rect 36636 30005 36645 30039
rect 36645 30005 36679 30039
rect 36679 30005 36688 30039
rect 36636 29996 36688 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2504 29792 2556 29844
rect 8208 29792 8260 29844
rect 2964 29724 3016 29776
rect 7472 29724 7524 29776
rect 7748 29724 7800 29776
rect 12992 29792 13044 29844
rect 18512 29792 18564 29844
rect 20260 29835 20312 29844
rect 20260 29801 20269 29835
rect 20269 29801 20303 29835
rect 20303 29801 20312 29835
rect 20260 29792 20312 29801
rect 15936 29724 15988 29776
rect 24952 29792 25004 29844
rect 24676 29724 24728 29776
rect 3332 29656 3384 29708
rect 9312 29699 9364 29708
rect 2596 29631 2648 29640
rect 2596 29597 2605 29631
rect 2605 29597 2639 29631
rect 2639 29597 2648 29631
rect 2596 29588 2648 29597
rect 2872 29631 2924 29640
rect 2872 29597 2881 29631
rect 2881 29597 2915 29631
rect 2915 29597 2924 29631
rect 2872 29588 2924 29597
rect 3424 29588 3476 29640
rect 9312 29665 9321 29699
rect 9321 29665 9355 29699
rect 9355 29665 9364 29699
rect 9312 29656 9364 29665
rect 16580 29656 16632 29708
rect 24124 29656 24176 29708
rect 26332 29792 26384 29844
rect 29828 29835 29880 29844
rect 29828 29801 29837 29835
rect 29837 29801 29871 29835
rect 29871 29801 29880 29835
rect 29828 29792 29880 29801
rect 31484 29792 31536 29844
rect 36636 29792 36688 29844
rect 30840 29724 30892 29776
rect 5172 29588 5224 29640
rect 9496 29588 9548 29640
rect 10508 29631 10560 29640
rect 10508 29597 10517 29631
rect 10517 29597 10551 29631
rect 10551 29597 10560 29631
rect 10508 29588 10560 29597
rect 19340 29588 19392 29640
rect 10784 29563 10836 29572
rect 10784 29529 10818 29563
rect 10818 29529 10836 29563
rect 2688 29452 2740 29504
rect 10784 29520 10836 29529
rect 15752 29520 15804 29572
rect 19984 29588 20036 29640
rect 22192 29588 22244 29640
rect 22560 29631 22612 29640
rect 22560 29597 22569 29631
rect 22569 29597 22603 29631
rect 22603 29597 22612 29631
rect 22560 29588 22612 29597
rect 22744 29631 22796 29640
rect 22744 29597 22753 29631
rect 22753 29597 22787 29631
rect 22787 29597 22796 29631
rect 22744 29588 22796 29597
rect 20076 29563 20128 29572
rect 20076 29529 20085 29563
rect 20085 29529 20119 29563
rect 20119 29529 20128 29563
rect 20076 29520 20128 29529
rect 27068 29656 27120 29708
rect 4712 29452 4764 29504
rect 4804 29452 4856 29504
rect 7748 29452 7800 29504
rect 9772 29452 9824 29504
rect 11060 29452 11112 29504
rect 11704 29452 11756 29504
rect 16580 29495 16632 29504
rect 16580 29461 16589 29495
rect 16589 29461 16623 29495
rect 16623 29461 16632 29495
rect 16580 29452 16632 29461
rect 16948 29452 17000 29504
rect 20352 29452 20404 29504
rect 23020 29452 23072 29504
rect 24584 29452 24636 29504
rect 29828 29588 29880 29640
rect 25596 29520 25648 29572
rect 31208 29631 31260 29640
rect 31208 29597 31217 29631
rect 31217 29597 31251 29631
rect 31251 29597 31260 29631
rect 31944 29631 31996 29640
rect 31208 29588 31260 29597
rect 31944 29597 31953 29631
rect 31953 29597 31987 29631
rect 31987 29597 31996 29631
rect 31944 29588 31996 29597
rect 36360 29656 36412 29708
rect 34612 29588 34664 29640
rect 35624 29588 35676 29640
rect 36084 29588 36136 29640
rect 37004 29631 37056 29640
rect 37004 29597 37013 29631
rect 37013 29597 37047 29631
rect 37047 29597 37056 29631
rect 37004 29588 37056 29597
rect 58164 29631 58216 29640
rect 58164 29597 58173 29631
rect 58173 29597 58207 29631
rect 58207 29597 58216 29631
rect 58164 29588 58216 29597
rect 32312 29520 32364 29572
rect 26424 29452 26476 29504
rect 30012 29452 30064 29504
rect 31208 29452 31260 29504
rect 33232 29452 33284 29504
rect 35532 29452 35584 29504
rect 37464 29495 37516 29504
rect 37464 29461 37473 29495
rect 37473 29461 37507 29495
rect 37507 29461 37516 29495
rect 37464 29452 37516 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 2872 29248 2924 29300
rect 2596 29180 2648 29232
rect 2872 28908 2924 28960
rect 10140 29248 10192 29300
rect 10416 29248 10468 29300
rect 10784 29291 10836 29300
rect 10784 29257 10793 29291
rect 10793 29257 10827 29291
rect 10827 29257 10836 29291
rect 10784 29248 10836 29257
rect 13728 29248 13780 29300
rect 5080 29180 5132 29232
rect 8208 29223 8260 29232
rect 8208 29189 8217 29223
rect 8217 29189 8251 29223
rect 8251 29189 8260 29223
rect 8208 29180 8260 29189
rect 8576 29223 8628 29232
rect 8576 29189 8585 29223
rect 8585 29189 8619 29223
rect 8619 29189 8628 29223
rect 8576 29180 8628 29189
rect 3700 29112 3752 29164
rect 4712 29155 4764 29164
rect 4712 29121 4721 29155
rect 4721 29121 4755 29155
rect 4755 29121 4764 29155
rect 4712 29112 4764 29121
rect 5172 29112 5224 29164
rect 3792 29044 3844 29096
rect 4896 28976 4948 29028
rect 7472 29019 7524 29028
rect 7472 28985 7481 29019
rect 7481 28985 7515 29019
rect 7515 28985 7524 29019
rect 7472 28976 7524 28985
rect 7748 29112 7800 29164
rect 9128 29112 9180 29164
rect 9220 29112 9272 29164
rect 9588 29112 9640 29164
rect 9772 29112 9824 29164
rect 10140 29155 10192 29164
rect 10140 29121 10149 29155
rect 10149 29121 10183 29155
rect 10183 29121 10192 29155
rect 10140 29112 10192 29121
rect 11704 29223 11756 29232
rect 11704 29189 11713 29223
rect 11713 29189 11747 29223
rect 11747 29189 11756 29223
rect 11704 29180 11756 29189
rect 14188 29180 14240 29232
rect 17132 29180 17184 29232
rect 10784 29112 10836 29164
rect 11980 29112 12032 29164
rect 15660 29155 15712 29164
rect 15660 29121 15669 29155
rect 15669 29121 15703 29155
rect 15703 29121 15712 29155
rect 15660 29112 15712 29121
rect 18512 29180 18564 29232
rect 19248 29180 19300 29232
rect 19432 29180 19484 29232
rect 23480 29248 23532 29300
rect 22560 29223 22612 29232
rect 18144 29112 18196 29164
rect 18788 29112 18840 29164
rect 19340 29112 19392 29164
rect 17408 29044 17460 29096
rect 9220 28976 9272 29028
rect 9404 28976 9456 29028
rect 17316 28976 17368 29028
rect 18052 28976 18104 29028
rect 18880 28976 18932 29028
rect 19984 29044 20036 29096
rect 21456 29112 21508 29164
rect 22560 29189 22569 29223
rect 22569 29189 22603 29223
rect 22603 29189 22612 29223
rect 22560 29180 22612 29189
rect 23296 29180 23348 29232
rect 24584 29248 24636 29300
rect 25504 29248 25556 29300
rect 30748 29248 30800 29300
rect 30840 29291 30892 29300
rect 30840 29257 30849 29291
rect 30849 29257 30883 29291
rect 30883 29257 30892 29291
rect 30840 29248 30892 29257
rect 23664 29112 23716 29164
rect 24216 29155 24268 29164
rect 24216 29121 24225 29155
rect 24225 29121 24259 29155
rect 24259 29121 24268 29155
rect 24216 29112 24268 29121
rect 24676 29180 24728 29232
rect 30012 29180 30064 29232
rect 30564 29180 30616 29232
rect 23756 29044 23808 29096
rect 24952 29112 25004 29164
rect 26148 29112 26200 29164
rect 30104 29112 30156 29164
rect 30840 29155 30892 29164
rect 30840 29121 30849 29155
rect 30849 29121 30883 29155
rect 30883 29121 30892 29155
rect 30840 29112 30892 29121
rect 20352 28976 20404 29028
rect 22836 28976 22888 29028
rect 23204 28976 23256 29028
rect 24124 28976 24176 29028
rect 30656 29044 30708 29096
rect 30748 29044 30800 29096
rect 34612 29248 34664 29300
rect 36268 29248 36320 29300
rect 35532 29180 35584 29232
rect 33416 29155 33468 29164
rect 33416 29121 33425 29155
rect 33425 29121 33459 29155
rect 33459 29121 33468 29155
rect 33416 29112 33468 29121
rect 35440 29155 35492 29164
rect 35440 29121 35449 29155
rect 35449 29121 35483 29155
rect 35483 29121 35492 29155
rect 35440 29112 35492 29121
rect 36084 29155 36136 29164
rect 36084 29121 36093 29155
rect 36093 29121 36127 29155
rect 36127 29121 36136 29155
rect 36084 29112 36136 29121
rect 37464 29180 37516 29232
rect 33600 29044 33652 29096
rect 34244 29044 34296 29096
rect 36544 29112 36596 29164
rect 39488 29087 39540 29096
rect 39488 29053 39497 29087
rect 39497 29053 39531 29087
rect 39531 29053 39540 29087
rect 39488 29044 39540 29053
rect 25596 28976 25648 29028
rect 26148 29019 26200 29028
rect 26148 28985 26157 29019
rect 26157 28985 26191 29019
rect 26191 28985 26200 29019
rect 26148 28976 26200 28985
rect 36452 28976 36504 29028
rect 38384 28976 38436 29028
rect 7380 28908 7432 28960
rect 9036 28951 9088 28960
rect 9036 28917 9045 28951
rect 9045 28917 9079 28951
rect 9079 28917 9088 28951
rect 9036 28908 9088 28917
rect 9312 28908 9364 28960
rect 10784 28908 10836 28960
rect 13636 28908 13688 28960
rect 15568 28908 15620 28960
rect 17132 28908 17184 28960
rect 20536 28908 20588 28960
rect 25872 28908 25924 28960
rect 30840 28908 30892 28960
rect 31392 28908 31444 28960
rect 36360 28908 36412 28960
rect 36544 28908 36596 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2688 28704 2740 28756
rect 3792 28747 3844 28756
rect 3792 28713 3801 28747
rect 3801 28713 3835 28747
rect 3835 28713 3844 28747
rect 3792 28704 3844 28713
rect 7564 28747 7616 28756
rect 7564 28713 7573 28747
rect 7573 28713 7607 28747
rect 7607 28713 7616 28747
rect 7564 28704 7616 28713
rect 9128 28704 9180 28756
rect 10784 28747 10836 28756
rect 10784 28713 10793 28747
rect 10793 28713 10827 28747
rect 10827 28713 10836 28747
rect 10784 28704 10836 28713
rect 13084 28704 13136 28756
rect 12532 28636 12584 28688
rect 12992 28636 13044 28688
rect 3700 28500 3752 28552
rect 3976 28543 4028 28552
rect 3976 28509 3985 28543
rect 3985 28509 4019 28543
rect 4019 28509 4028 28543
rect 3976 28500 4028 28509
rect 4988 28543 5040 28552
rect 4988 28509 4997 28543
rect 4997 28509 5031 28543
rect 5031 28509 5040 28543
rect 4988 28500 5040 28509
rect 5172 28500 5224 28552
rect 3608 28432 3660 28484
rect 7656 28475 7708 28484
rect 4712 28364 4764 28416
rect 7656 28441 7665 28475
rect 7665 28441 7699 28475
rect 7699 28441 7708 28475
rect 7656 28432 7708 28441
rect 6368 28364 6420 28416
rect 9772 28500 9824 28552
rect 10508 28500 10560 28552
rect 9036 28432 9088 28484
rect 9496 28364 9548 28416
rect 11888 28364 11940 28416
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 13360 28543 13412 28552
rect 13360 28509 13369 28543
rect 13369 28509 13403 28543
rect 13403 28509 13412 28543
rect 13360 28500 13412 28509
rect 13728 28500 13780 28552
rect 15660 28704 15712 28756
rect 17224 28704 17276 28756
rect 24952 28704 25004 28756
rect 25780 28704 25832 28756
rect 34336 28704 34388 28756
rect 36360 28704 36412 28756
rect 37004 28704 37056 28756
rect 19432 28636 19484 28688
rect 21456 28636 21508 28688
rect 14188 28543 14240 28552
rect 14188 28509 14198 28543
rect 14198 28509 14232 28543
rect 14232 28509 14240 28543
rect 17960 28568 18012 28620
rect 20076 28568 20128 28620
rect 14188 28500 14240 28509
rect 14556 28543 14608 28552
rect 14556 28509 14570 28543
rect 14570 28509 14604 28543
rect 14604 28509 14608 28543
rect 14556 28500 14608 28509
rect 15200 28500 15252 28552
rect 17132 28500 17184 28552
rect 19984 28500 20036 28552
rect 22100 28568 22152 28620
rect 22744 28568 22796 28620
rect 30564 28568 30616 28620
rect 33508 28611 33560 28620
rect 33508 28577 33517 28611
rect 33517 28577 33551 28611
rect 33551 28577 33560 28611
rect 33508 28568 33560 28577
rect 14832 28432 14884 28484
rect 16028 28432 16080 28484
rect 13636 28364 13688 28416
rect 15200 28364 15252 28416
rect 17316 28364 17368 28416
rect 17500 28364 17552 28416
rect 21088 28407 21140 28416
rect 21088 28373 21097 28407
rect 21097 28373 21131 28407
rect 21131 28373 21140 28407
rect 21088 28364 21140 28373
rect 21456 28475 21508 28484
rect 21456 28441 21465 28475
rect 21465 28441 21499 28475
rect 21499 28441 21508 28475
rect 21456 28432 21508 28441
rect 23296 28500 23348 28552
rect 24124 28500 24176 28552
rect 30748 28543 30800 28552
rect 30748 28509 30757 28543
rect 30757 28509 30791 28543
rect 30791 28509 30800 28543
rect 30748 28500 30800 28509
rect 31392 28543 31444 28552
rect 25136 28475 25188 28484
rect 22192 28364 22244 28416
rect 25136 28441 25145 28475
rect 25145 28441 25179 28475
rect 25179 28441 25188 28475
rect 25136 28432 25188 28441
rect 30104 28432 30156 28484
rect 31392 28509 31401 28543
rect 31401 28509 31435 28543
rect 31435 28509 31444 28543
rect 31392 28500 31444 28509
rect 33416 28500 33468 28552
rect 35348 28500 35400 28552
rect 35532 28500 35584 28552
rect 36268 28543 36320 28552
rect 36268 28509 36277 28543
rect 36277 28509 36311 28543
rect 36311 28509 36320 28543
rect 36268 28500 36320 28509
rect 38384 28543 38436 28552
rect 38384 28509 38402 28543
rect 38402 28509 38436 28543
rect 38384 28500 38436 28509
rect 39488 28500 39540 28552
rect 39948 28500 40000 28552
rect 33600 28432 33652 28484
rect 22744 28407 22796 28416
rect 22744 28373 22753 28407
rect 22753 28373 22787 28407
rect 22787 28373 22796 28407
rect 23756 28407 23808 28416
rect 22744 28364 22796 28373
rect 23756 28373 23765 28407
rect 23765 28373 23799 28407
rect 23799 28373 23808 28407
rect 23756 28364 23808 28373
rect 24584 28364 24636 28416
rect 31852 28364 31904 28416
rect 34796 28364 34848 28416
rect 35440 28364 35492 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 3976 28203 4028 28212
rect 3976 28169 3985 28203
rect 3985 28169 4019 28203
rect 4019 28169 4028 28203
rect 3976 28160 4028 28169
rect 9404 28203 9456 28212
rect 9404 28169 9413 28203
rect 9413 28169 9447 28203
rect 9447 28169 9456 28203
rect 9404 28160 9456 28169
rect 10048 28203 10100 28212
rect 10048 28169 10057 28203
rect 10057 28169 10091 28203
rect 10091 28169 10100 28203
rect 10048 28160 10100 28169
rect 10784 28160 10836 28212
rect 12440 28160 12492 28212
rect 13084 28203 13136 28212
rect 6736 28135 6788 28144
rect 6736 28101 6745 28135
rect 6745 28101 6779 28135
rect 6779 28101 6788 28135
rect 6736 28092 6788 28101
rect 9220 28092 9272 28144
rect 13084 28169 13093 28203
rect 13093 28169 13127 28203
rect 13127 28169 13136 28203
rect 13084 28160 13136 28169
rect 13360 28160 13412 28212
rect 16028 28203 16080 28212
rect 16028 28169 16037 28203
rect 16037 28169 16071 28203
rect 16071 28169 16080 28203
rect 16028 28160 16080 28169
rect 17132 28160 17184 28212
rect 13452 28092 13504 28144
rect 14648 28092 14700 28144
rect 2872 28067 2924 28076
rect 2872 28033 2906 28067
rect 2906 28033 2924 28067
rect 2872 28024 2924 28033
rect 6368 28067 6420 28076
rect 6368 28033 6377 28067
rect 6377 28033 6411 28067
rect 6411 28033 6420 28067
rect 6368 28024 6420 28033
rect 6460 28067 6512 28076
rect 6460 28033 6470 28067
rect 6470 28033 6504 28067
rect 6504 28033 6512 28067
rect 6460 28024 6512 28033
rect 6644 28067 6696 28076
rect 6644 28033 6653 28067
rect 6653 28033 6687 28067
rect 6687 28033 6696 28067
rect 6644 28024 6696 28033
rect 6828 28067 6880 28076
rect 6828 28033 6842 28067
rect 6842 28033 6876 28067
rect 6876 28033 6880 28067
rect 6828 28024 6880 28033
rect 8944 28024 8996 28076
rect 9496 28067 9548 28076
rect 9496 28033 9505 28067
rect 9505 28033 9539 28067
rect 9539 28033 9548 28067
rect 9496 28024 9548 28033
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 11888 28067 11940 28076
rect 11888 28033 11897 28067
rect 11897 28033 11931 28067
rect 11931 28033 11940 28067
rect 11888 28024 11940 28033
rect 12532 28067 12584 28076
rect 12532 28033 12541 28067
rect 12541 28033 12575 28067
rect 12575 28033 12584 28067
rect 12532 28024 12584 28033
rect 12624 28024 12676 28076
rect 13268 28024 13320 28076
rect 15384 28067 15436 28076
rect 15384 28033 15393 28067
rect 15393 28033 15427 28067
rect 15427 28033 15436 28067
rect 15384 28024 15436 28033
rect 15568 28067 15620 28076
rect 15568 28033 15577 28067
rect 15577 28033 15611 28067
rect 15611 28033 15620 28067
rect 15568 28024 15620 28033
rect 2596 27999 2648 28008
rect 2596 27965 2605 27999
rect 2605 27965 2639 27999
rect 2639 27965 2648 27999
rect 2596 27956 2648 27965
rect 13636 27956 13688 28008
rect 17224 28024 17276 28076
rect 23756 28092 23808 28144
rect 19432 28024 19484 28076
rect 19984 28067 20036 28076
rect 19984 28033 19993 28067
rect 19993 28033 20027 28067
rect 20027 28033 20036 28067
rect 19984 28024 20036 28033
rect 17684 27956 17736 28008
rect 19340 27956 19392 28008
rect 17960 27888 18012 27940
rect 7012 27863 7064 27872
rect 7012 27829 7021 27863
rect 7021 27829 7055 27863
rect 7055 27829 7064 27863
rect 7012 27820 7064 27829
rect 8944 27820 8996 27872
rect 11060 27820 11112 27872
rect 13268 27820 13320 27872
rect 21180 27888 21232 27940
rect 21640 27888 21692 27940
rect 35440 28092 35492 28144
rect 26424 28067 26476 28076
rect 26424 28033 26433 28067
rect 26433 28033 26467 28067
rect 26467 28033 26476 28067
rect 26424 28024 26476 28033
rect 29368 28024 29420 28076
rect 30104 28024 30156 28076
rect 30748 28024 30800 28076
rect 33416 28024 33468 28076
rect 34520 28067 34572 28076
rect 25136 27888 25188 27940
rect 26608 27888 26660 27940
rect 19156 27863 19208 27872
rect 19156 27829 19165 27863
rect 19165 27829 19199 27863
rect 19199 27829 19208 27863
rect 19156 27820 19208 27829
rect 26700 27820 26752 27872
rect 27068 27863 27120 27872
rect 27068 27829 27077 27863
rect 27077 27829 27111 27863
rect 27111 27829 27120 27863
rect 27068 27820 27120 27829
rect 28724 27820 28776 27872
rect 30472 27956 30524 28008
rect 33140 27956 33192 28008
rect 33600 27956 33652 28008
rect 34520 28033 34529 28067
rect 34529 28033 34563 28067
rect 34563 28033 34572 28067
rect 34520 28024 34572 28033
rect 39856 28024 39908 28076
rect 39948 27999 40000 28008
rect 39948 27965 39957 27999
rect 39957 27965 39991 27999
rect 39991 27965 40000 27999
rect 39948 27956 40000 27965
rect 58164 27931 58216 27940
rect 58164 27897 58173 27931
rect 58173 27897 58207 27931
rect 58207 27897 58216 27931
rect 58164 27888 58216 27897
rect 33968 27863 34020 27872
rect 33968 27829 33977 27863
rect 33977 27829 34011 27863
rect 34011 27829 34020 27863
rect 33968 27820 34020 27829
rect 39028 27820 39080 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 7656 27616 7708 27668
rect 10416 27616 10468 27668
rect 13452 27616 13504 27668
rect 17224 27616 17276 27668
rect 4896 27455 4948 27464
rect 4896 27421 4905 27455
rect 4905 27421 4939 27455
rect 4939 27421 4948 27455
rect 4896 27412 4948 27421
rect 5448 27548 5500 27600
rect 6828 27548 6880 27600
rect 9312 27548 9364 27600
rect 4068 27344 4120 27396
rect 5540 27412 5592 27464
rect 7104 27480 7156 27532
rect 9680 27548 9732 27600
rect 29000 27591 29052 27600
rect 29000 27557 29009 27591
rect 29009 27557 29043 27591
rect 29043 27557 29052 27591
rect 29000 27548 29052 27557
rect 30472 27591 30524 27600
rect 30472 27557 30481 27591
rect 30481 27557 30515 27591
rect 30515 27557 30524 27591
rect 30472 27548 30524 27557
rect 6460 27412 6512 27464
rect 8944 27455 8996 27464
rect 8944 27421 8953 27455
rect 8953 27421 8987 27455
rect 8987 27421 8996 27455
rect 8944 27412 8996 27421
rect 5080 27344 5132 27396
rect 6644 27344 6696 27396
rect 7104 27387 7156 27396
rect 6828 27276 6880 27328
rect 7104 27353 7113 27387
rect 7113 27353 7147 27387
rect 7147 27353 7156 27387
rect 7104 27344 7156 27353
rect 9404 27412 9456 27464
rect 9496 27412 9548 27464
rect 10600 27480 10652 27532
rect 16028 27480 16080 27532
rect 24400 27480 24452 27532
rect 10692 27412 10744 27464
rect 7656 27276 7708 27328
rect 12900 27412 12952 27464
rect 17960 27412 18012 27464
rect 19156 27412 19208 27464
rect 20628 27344 20680 27396
rect 21548 27344 21600 27396
rect 26148 27387 26200 27396
rect 12440 27276 12492 27328
rect 16212 27276 16264 27328
rect 16580 27276 16632 27328
rect 18420 27319 18472 27328
rect 18420 27285 18429 27319
rect 18429 27285 18463 27319
rect 18463 27285 18472 27319
rect 18420 27276 18472 27285
rect 19984 27276 20036 27328
rect 24676 27319 24728 27328
rect 24676 27285 24685 27319
rect 24685 27285 24719 27319
rect 24719 27285 24728 27319
rect 24676 27276 24728 27285
rect 24860 27276 24912 27328
rect 26148 27353 26157 27387
rect 26157 27353 26191 27387
rect 26191 27353 26200 27387
rect 26148 27344 26200 27353
rect 26700 27412 26752 27464
rect 29000 27412 29052 27464
rect 32772 27412 32824 27464
rect 33232 27412 33284 27464
rect 33416 27412 33468 27464
rect 34704 27480 34756 27532
rect 33784 27412 33836 27464
rect 26884 27387 26936 27396
rect 26884 27353 26918 27387
rect 26918 27353 26936 27387
rect 26884 27344 26936 27353
rect 27160 27344 27212 27396
rect 28724 27344 28776 27396
rect 27620 27276 27672 27328
rect 27988 27319 28040 27328
rect 27988 27285 27997 27319
rect 27997 27285 28031 27319
rect 28031 27285 28040 27319
rect 27988 27276 28040 27285
rect 28632 27276 28684 27328
rect 33140 27344 33192 27396
rect 34612 27344 34664 27396
rect 29644 27276 29696 27328
rect 32312 27319 32364 27328
rect 32312 27285 32321 27319
rect 32321 27285 32355 27319
rect 32355 27285 32364 27319
rect 32312 27276 32364 27285
rect 33508 27276 33560 27328
rect 34428 27276 34480 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 2780 27072 2832 27124
rect 4620 27072 4672 27124
rect 3976 27004 4028 27056
rect 5080 27047 5132 27056
rect 4804 26979 4856 26988
rect 4804 26945 4813 26979
rect 4813 26945 4847 26979
rect 4847 26945 4856 26979
rect 4804 26936 4856 26945
rect 5080 27013 5089 27047
rect 5089 27013 5123 27047
rect 5123 27013 5132 27047
rect 5080 27004 5132 27013
rect 6460 27072 6512 27124
rect 11520 27115 11572 27124
rect 5448 27004 5500 27056
rect 7104 27004 7156 27056
rect 7748 27004 7800 27056
rect 10968 27047 11020 27056
rect 5540 26936 5592 26988
rect 7472 26979 7524 26988
rect 7472 26945 7490 26979
rect 7490 26945 7524 26979
rect 7472 26936 7524 26945
rect 9312 26979 9364 26988
rect 9312 26945 9321 26979
rect 9321 26945 9355 26979
rect 9355 26945 9364 26979
rect 9312 26936 9364 26945
rect 10968 27013 10977 27047
rect 10977 27013 11011 27047
rect 11011 27013 11020 27047
rect 10968 27004 11020 27013
rect 11520 27081 11529 27115
rect 11529 27081 11563 27115
rect 11563 27081 11572 27115
rect 11520 27072 11572 27081
rect 16028 27115 16080 27124
rect 16028 27081 16037 27115
rect 16037 27081 16071 27115
rect 16071 27081 16080 27115
rect 16028 27072 16080 27081
rect 16856 27072 16908 27124
rect 17408 27072 17460 27124
rect 18420 27072 18472 27124
rect 25596 27072 25648 27124
rect 26884 27072 26936 27124
rect 9864 26936 9916 26988
rect 12624 26936 12676 26988
rect 19616 27004 19668 27056
rect 20536 27004 20588 27056
rect 21180 27047 21232 27056
rect 21180 27013 21189 27047
rect 21189 27013 21223 27047
rect 21223 27013 21232 27047
rect 21180 27004 21232 27013
rect 21916 27004 21968 27056
rect 5448 26868 5500 26920
rect 7748 26911 7800 26920
rect 7748 26877 7757 26911
rect 7757 26877 7791 26911
rect 7791 26877 7800 26911
rect 7748 26868 7800 26877
rect 9772 26868 9824 26920
rect 10600 26868 10652 26920
rect 11980 26868 12032 26920
rect 13360 26868 13412 26920
rect 16212 26868 16264 26920
rect 17592 26936 17644 26988
rect 18144 26936 18196 26988
rect 19892 26936 19944 26988
rect 22468 26979 22520 26988
rect 22468 26945 22502 26979
rect 22502 26945 22520 26979
rect 22468 26936 22520 26945
rect 18236 26868 18288 26920
rect 20536 26868 20588 26920
rect 3240 26800 3292 26852
rect 8484 26800 8536 26852
rect 18328 26800 18380 26852
rect 3056 26732 3108 26784
rect 5448 26775 5500 26784
rect 5448 26741 5457 26775
rect 5457 26741 5491 26775
rect 5491 26741 5500 26775
rect 5448 26732 5500 26741
rect 6092 26732 6144 26784
rect 9956 26732 10008 26784
rect 18696 26732 18748 26784
rect 22560 26732 22612 26784
rect 25780 27004 25832 27056
rect 31392 27072 31444 27124
rect 32404 27072 32456 27124
rect 34244 27072 34296 27124
rect 29092 27004 29144 27056
rect 24676 26936 24728 26988
rect 24768 26868 24820 26920
rect 25136 26800 25188 26852
rect 27712 26936 27764 26988
rect 31208 27004 31260 27056
rect 32404 26979 32456 26988
rect 32404 26945 32413 26979
rect 32413 26945 32447 26979
rect 32447 26945 32456 26979
rect 32404 26936 32456 26945
rect 32588 26979 32640 26988
rect 32588 26945 32597 26979
rect 32597 26945 32631 26979
rect 32631 26945 32640 26979
rect 32588 26936 32640 26945
rect 34244 26979 34296 26988
rect 31944 26868 31996 26920
rect 34244 26945 34253 26979
rect 34253 26945 34287 26979
rect 34287 26945 34296 26979
rect 34244 26936 34296 26945
rect 34428 26979 34480 26988
rect 34428 26945 34437 26979
rect 34437 26945 34471 26979
rect 34471 26945 34480 26979
rect 34428 26936 34480 26945
rect 35624 27004 35676 27056
rect 31852 26800 31904 26852
rect 32864 26800 32916 26852
rect 40500 26936 40552 26988
rect 39948 26911 40000 26920
rect 39948 26877 39957 26911
rect 39957 26877 39991 26911
rect 39991 26877 40000 26911
rect 39948 26868 40000 26877
rect 25596 26732 25648 26784
rect 25872 26732 25924 26784
rect 28172 26775 28224 26784
rect 28172 26741 28181 26775
rect 28181 26741 28215 26775
rect 28215 26741 28224 26775
rect 28172 26732 28224 26741
rect 33600 26732 33652 26784
rect 35808 26732 35860 26784
rect 37096 26732 37148 26784
rect 40040 26732 40092 26784
rect 58164 26775 58216 26784
rect 58164 26741 58173 26775
rect 58173 26741 58207 26775
rect 58207 26741 58216 26775
rect 58164 26732 58216 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5724 26528 5776 26580
rect 7472 26528 7524 26580
rect 11704 26571 11756 26580
rect 11704 26537 11713 26571
rect 11713 26537 11747 26571
rect 11747 26537 11756 26571
rect 11704 26528 11756 26537
rect 18328 26528 18380 26580
rect 19892 26571 19944 26580
rect 6092 26460 6144 26512
rect 7564 26460 7616 26512
rect 7656 26460 7708 26512
rect 2780 26324 2832 26376
rect 3148 26392 3200 26444
rect 3056 26367 3108 26376
rect 3056 26333 3065 26367
rect 3065 26333 3099 26367
rect 3099 26333 3108 26367
rect 3056 26324 3108 26333
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 4068 26324 4120 26376
rect 6092 26367 6144 26376
rect 6092 26333 6101 26367
rect 6101 26333 6135 26367
rect 6135 26333 6144 26367
rect 6092 26324 6144 26333
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 5356 26256 5408 26308
rect 5724 26256 5776 26308
rect 7472 26324 7524 26376
rect 14556 26460 14608 26512
rect 19340 26460 19392 26512
rect 19892 26537 19901 26571
rect 19901 26537 19935 26571
rect 19935 26537 19944 26571
rect 19892 26528 19944 26537
rect 22468 26528 22520 26580
rect 24308 26528 24360 26580
rect 28632 26528 28684 26580
rect 29000 26528 29052 26580
rect 30288 26528 30340 26580
rect 34704 26571 34756 26580
rect 17776 26392 17828 26444
rect 8208 26324 8260 26376
rect 6552 26256 6604 26308
rect 11520 26324 11572 26376
rect 17408 26324 17460 26376
rect 17960 26324 18012 26376
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 20076 26324 20128 26376
rect 20444 26367 20496 26376
rect 20444 26333 20453 26367
rect 20453 26333 20487 26367
rect 20487 26333 20496 26367
rect 20444 26324 20496 26333
rect 20628 26367 20680 26376
rect 20628 26333 20637 26367
rect 20637 26333 20671 26367
rect 20671 26333 20680 26367
rect 20628 26324 20680 26333
rect 20812 26367 20864 26376
rect 20812 26333 20821 26367
rect 20821 26333 20855 26367
rect 20855 26333 20864 26367
rect 20812 26324 20864 26333
rect 11980 26256 12032 26308
rect 12440 26299 12492 26308
rect 12440 26265 12449 26299
rect 12449 26265 12483 26299
rect 12483 26265 12492 26299
rect 12440 26256 12492 26265
rect 17316 26256 17368 26308
rect 21732 26367 21784 26376
rect 21732 26333 21741 26367
rect 21741 26333 21775 26367
rect 21775 26333 21784 26367
rect 21732 26324 21784 26333
rect 22468 26392 22520 26444
rect 21916 26367 21968 26376
rect 21916 26333 21925 26367
rect 21925 26333 21959 26367
rect 21959 26333 21968 26367
rect 21916 26324 21968 26333
rect 22560 26324 22612 26376
rect 24584 26367 24636 26376
rect 24584 26333 24593 26367
rect 24593 26333 24627 26367
rect 24627 26333 24636 26367
rect 24584 26324 24636 26333
rect 24860 26460 24912 26512
rect 25136 26392 25188 26444
rect 27620 26392 27672 26444
rect 28724 26392 28776 26444
rect 25596 26324 25648 26376
rect 26792 26324 26844 26376
rect 34704 26537 34713 26571
rect 34713 26537 34747 26571
rect 34747 26537 34756 26571
rect 34704 26528 34756 26537
rect 31944 26392 31996 26444
rect 35808 26367 35860 26376
rect 35808 26333 35826 26367
rect 35826 26333 35860 26367
rect 35808 26324 35860 26333
rect 37188 26324 37240 26376
rect 37372 26324 37424 26376
rect 21640 26256 21692 26308
rect 2872 26188 2924 26240
rect 3056 26188 3108 26240
rect 6736 26231 6788 26240
rect 6736 26197 6745 26231
rect 6745 26197 6779 26231
rect 6779 26197 6788 26231
rect 6736 26188 6788 26197
rect 10600 26231 10652 26240
rect 10600 26197 10609 26231
rect 10609 26197 10643 26231
rect 10643 26197 10652 26231
rect 10600 26188 10652 26197
rect 12348 26188 12400 26240
rect 20260 26188 20312 26240
rect 21456 26188 21508 26240
rect 26148 26256 26200 26308
rect 28172 26256 28224 26308
rect 29736 26256 29788 26308
rect 39120 26299 39172 26308
rect 39120 26265 39129 26299
rect 39129 26265 39163 26299
rect 39163 26265 39172 26299
rect 39120 26256 39172 26265
rect 40316 26324 40368 26376
rect 40040 26299 40092 26308
rect 40040 26265 40049 26299
rect 40049 26265 40083 26299
rect 40083 26265 40092 26299
rect 40040 26256 40092 26265
rect 25780 26188 25832 26240
rect 41144 26188 41196 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 3976 26027 4028 26036
rect 3976 25993 3985 26027
rect 3985 25993 4019 26027
rect 4019 25993 4028 26027
rect 3976 25984 4028 25993
rect 6276 25984 6328 26036
rect 9496 25984 9548 26036
rect 12440 25984 12492 26036
rect 13636 25984 13688 26036
rect 17316 26027 17368 26036
rect 17316 25993 17325 26027
rect 17325 25993 17359 26027
rect 17359 25993 17368 26027
rect 17316 25984 17368 25993
rect 17776 25984 17828 26036
rect 19432 25984 19484 26036
rect 20628 25984 20680 26036
rect 2872 25959 2924 25968
rect 2872 25925 2906 25959
rect 2906 25925 2924 25959
rect 2872 25916 2924 25925
rect 5356 25916 5408 25968
rect 7288 25959 7340 25968
rect 2596 25891 2648 25900
rect 2596 25857 2605 25891
rect 2605 25857 2639 25891
rect 2639 25857 2648 25891
rect 2596 25848 2648 25857
rect 6920 25891 6972 25900
rect 6920 25857 6929 25891
rect 6929 25857 6963 25891
rect 6963 25857 6972 25891
rect 6920 25848 6972 25857
rect 7288 25925 7297 25959
rect 7297 25925 7331 25959
rect 7331 25925 7340 25959
rect 7288 25916 7340 25925
rect 9312 25959 9364 25968
rect 9312 25925 9321 25959
rect 9321 25925 9355 25959
rect 9355 25925 9364 25959
rect 9312 25916 9364 25925
rect 9404 25916 9456 25968
rect 7104 25848 7156 25900
rect 9496 25891 9548 25900
rect 9496 25857 9505 25891
rect 9505 25857 9539 25891
rect 9539 25857 9548 25891
rect 9496 25848 9548 25857
rect 12348 25848 12400 25900
rect 13268 25848 13320 25900
rect 16028 25848 16080 25900
rect 16856 25891 16908 25900
rect 16856 25857 16865 25891
rect 16865 25857 16899 25891
rect 16899 25857 16908 25891
rect 16856 25848 16908 25857
rect 17132 25848 17184 25900
rect 17500 25848 17552 25900
rect 18788 25916 18840 25968
rect 20260 25916 20312 25968
rect 20812 25916 20864 25968
rect 21456 25916 21508 25968
rect 21640 25916 21692 25968
rect 25136 25916 25188 25968
rect 27712 25984 27764 26036
rect 32772 26027 32824 26036
rect 32772 25993 32781 26027
rect 32781 25993 32815 26027
rect 32815 25993 32824 26027
rect 32772 25984 32824 25993
rect 37280 25984 37332 26036
rect 9864 25780 9916 25832
rect 10876 25780 10928 25832
rect 13728 25780 13780 25832
rect 18144 25848 18196 25900
rect 18696 25891 18748 25900
rect 18696 25857 18705 25891
rect 18705 25857 18739 25891
rect 18739 25857 18748 25891
rect 18696 25848 18748 25857
rect 19432 25848 19484 25900
rect 20536 25780 20588 25832
rect 8300 25712 8352 25764
rect 17316 25712 17368 25764
rect 19064 25712 19116 25764
rect 24584 25848 24636 25900
rect 24952 25848 25004 25900
rect 25780 25891 25832 25900
rect 25780 25857 25802 25891
rect 25802 25857 25832 25891
rect 25780 25848 25832 25857
rect 25872 25891 25924 25900
rect 25872 25857 25881 25891
rect 25881 25857 25915 25891
rect 25915 25857 25924 25891
rect 25872 25848 25924 25857
rect 27068 25916 27120 25968
rect 28632 25959 28684 25968
rect 28632 25925 28641 25959
rect 28641 25925 28675 25959
rect 28675 25925 28684 25959
rect 28632 25916 28684 25925
rect 33600 25916 33652 25968
rect 28908 25848 28960 25900
rect 30012 25891 30064 25900
rect 30012 25857 30021 25891
rect 30021 25857 30055 25891
rect 30055 25857 30064 25891
rect 30012 25848 30064 25857
rect 34152 25823 34204 25832
rect 34152 25789 34161 25823
rect 34161 25789 34195 25823
rect 34195 25789 34204 25823
rect 34152 25780 34204 25789
rect 37188 25712 37240 25764
rect 39948 25712 40000 25764
rect 6184 25644 6236 25696
rect 7472 25644 7524 25696
rect 8208 25644 8260 25696
rect 15016 25644 15068 25696
rect 17224 25644 17276 25696
rect 18144 25644 18196 25696
rect 20444 25644 20496 25696
rect 22836 25644 22888 25696
rect 29552 25644 29604 25696
rect 30472 25644 30524 25696
rect 31300 25644 31352 25696
rect 37832 25644 37884 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 7104 25440 7156 25492
rect 16304 25440 16356 25492
rect 22192 25440 22244 25492
rect 24676 25440 24728 25492
rect 24768 25440 24820 25492
rect 31300 25440 31352 25492
rect 39856 25483 39908 25492
rect 9956 25372 10008 25424
rect 20076 25415 20128 25424
rect 20076 25381 20085 25415
rect 20085 25381 20119 25415
rect 20119 25381 20128 25415
rect 20076 25372 20128 25381
rect 21548 25372 21600 25424
rect 27804 25372 27856 25424
rect 2596 25236 2648 25288
rect 2872 25279 2924 25288
rect 2872 25245 2881 25279
rect 2881 25245 2915 25279
rect 2915 25245 2924 25279
rect 2872 25236 2924 25245
rect 3148 25304 3200 25356
rect 11796 25304 11848 25356
rect 17592 25304 17644 25356
rect 18236 25304 18288 25356
rect 18420 25304 18472 25356
rect 19248 25304 19300 25356
rect 30012 25372 30064 25424
rect 39856 25449 39865 25483
rect 39865 25449 39899 25483
rect 39899 25449 39908 25483
rect 39856 25440 39908 25449
rect 40500 25440 40552 25492
rect 40132 25372 40184 25424
rect 3056 25279 3108 25288
rect 3056 25245 3065 25279
rect 3065 25245 3099 25279
rect 3099 25245 3108 25279
rect 3056 25236 3108 25245
rect 3240 25279 3292 25288
rect 3240 25245 3249 25279
rect 3249 25245 3283 25279
rect 3283 25245 3292 25279
rect 3240 25236 3292 25245
rect 7748 25236 7800 25288
rect 10876 25236 10928 25288
rect 12348 25236 12400 25288
rect 18696 25236 18748 25288
rect 6460 25168 6512 25220
rect 6736 25168 6788 25220
rect 2872 25100 2924 25152
rect 11428 25143 11480 25152
rect 11428 25109 11437 25143
rect 11437 25109 11471 25143
rect 11471 25109 11480 25143
rect 11428 25100 11480 25109
rect 13268 25143 13320 25152
rect 13268 25109 13277 25143
rect 13277 25109 13311 25143
rect 13311 25109 13320 25143
rect 13268 25100 13320 25109
rect 14648 25100 14700 25152
rect 15016 25168 15068 25220
rect 21364 25236 21416 25288
rect 21916 25211 21968 25220
rect 15568 25100 15620 25152
rect 17132 25100 17184 25152
rect 19340 25143 19392 25152
rect 19340 25109 19349 25143
rect 19349 25109 19383 25143
rect 19383 25109 19392 25143
rect 19340 25100 19392 25109
rect 20812 25100 20864 25152
rect 21916 25177 21925 25211
rect 21925 25177 21959 25211
rect 21959 25177 21968 25211
rect 21916 25168 21968 25177
rect 22652 25236 22704 25288
rect 25228 25236 25280 25288
rect 26148 25279 26200 25288
rect 26148 25245 26157 25279
rect 26157 25245 26191 25279
rect 26191 25245 26200 25279
rect 26148 25236 26200 25245
rect 29000 25236 29052 25288
rect 26792 25211 26844 25220
rect 26792 25177 26801 25211
rect 26801 25177 26835 25211
rect 26835 25177 26844 25211
rect 26792 25168 26844 25177
rect 30472 25279 30524 25288
rect 30472 25245 30481 25279
rect 30481 25245 30515 25279
rect 30515 25245 30524 25279
rect 30472 25236 30524 25245
rect 30564 25279 30616 25288
rect 30564 25245 30573 25279
rect 30573 25245 30607 25279
rect 30607 25245 30616 25279
rect 30564 25236 30616 25245
rect 31300 25236 31352 25288
rect 31944 25236 31996 25288
rect 34152 25236 34204 25288
rect 37188 25236 37240 25288
rect 37832 25279 37884 25288
rect 37832 25245 37841 25279
rect 37841 25245 37875 25279
rect 37875 25245 37884 25279
rect 37832 25236 37884 25245
rect 38016 25279 38068 25288
rect 38016 25245 38025 25279
rect 38025 25245 38059 25279
rect 38059 25245 38068 25279
rect 38016 25236 38068 25245
rect 40132 25279 40184 25288
rect 40132 25245 40141 25279
rect 40141 25245 40175 25279
rect 40175 25245 40184 25279
rect 40132 25236 40184 25245
rect 40868 25304 40920 25356
rect 40316 25279 40368 25288
rect 40316 25245 40325 25279
rect 40325 25245 40359 25279
rect 40359 25245 40368 25279
rect 40316 25236 40368 25245
rect 41144 25279 41196 25288
rect 39764 25168 39816 25220
rect 41144 25245 41153 25279
rect 41153 25245 41187 25279
rect 41187 25245 41196 25279
rect 41144 25236 41196 25245
rect 58164 25279 58216 25288
rect 27988 25100 28040 25152
rect 29000 25100 29052 25152
rect 29828 25143 29880 25152
rect 29828 25109 29837 25143
rect 29837 25109 29871 25143
rect 29871 25109 29880 25143
rect 29828 25100 29880 25109
rect 36176 25100 36228 25152
rect 41236 25100 41288 25152
rect 58164 25245 58173 25279
rect 58173 25245 58207 25279
rect 58207 25245 58216 25279
rect 58164 25236 58216 25245
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 6552 24896 6604 24948
rect 8208 24896 8260 24948
rect 11428 24896 11480 24948
rect 16304 24896 16356 24948
rect 2872 24871 2924 24880
rect 2872 24837 2906 24871
rect 2906 24837 2924 24871
rect 2872 24828 2924 24837
rect 9680 24828 9732 24880
rect 2596 24803 2648 24812
rect 2596 24769 2605 24803
rect 2605 24769 2639 24803
rect 2639 24769 2648 24803
rect 2596 24760 2648 24769
rect 3332 24760 3384 24812
rect 6276 24760 6328 24812
rect 7012 24760 7064 24812
rect 7932 24692 7984 24744
rect 8208 24692 8260 24744
rect 9036 24692 9088 24744
rect 9937 24803 9989 24812
rect 9937 24769 9962 24803
rect 9962 24769 9989 24803
rect 9937 24760 9989 24769
rect 10324 24760 10376 24812
rect 15384 24828 15436 24880
rect 14096 24760 14148 24812
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 18144 24803 18196 24812
rect 18144 24769 18153 24803
rect 18153 24769 18187 24803
rect 18187 24769 18196 24803
rect 18144 24760 18196 24769
rect 19340 24896 19392 24948
rect 23664 24896 23716 24948
rect 20536 24828 20588 24880
rect 21916 24828 21968 24880
rect 19340 24803 19392 24812
rect 19340 24769 19374 24803
rect 19374 24769 19392 24803
rect 10784 24692 10836 24744
rect 4068 24624 4120 24676
rect 13636 24667 13688 24676
rect 13636 24633 13645 24667
rect 13645 24633 13679 24667
rect 13679 24633 13688 24667
rect 13636 24624 13688 24633
rect 17776 24692 17828 24744
rect 19340 24760 19392 24769
rect 21364 24760 21416 24812
rect 6276 24556 6328 24608
rect 9036 24599 9088 24608
rect 9036 24565 9045 24599
rect 9045 24565 9079 24599
rect 9079 24565 9088 24599
rect 9036 24556 9088 24565
rect 9588 24599 9640 24608
rect 9588 24565 9597 24599
rect 9597 24565 9631 24599
rect 9631 24565 9640 24599
rect 9588 24556 9640 24565
rect 11612 24599 11664 24608
rect 11612 24565 11621 24599
rect 11621 24565 11655 24599
rect 11655 24565 11664 24599
rect 11612 24556 11664 24565
rect 12900 24556 12952 24608
rect 14188 24556 14240 24608
rect 17408 24624 17460 24676
rect 22652 24803 22704 24812
rect 22652 24769 22661 24803
rect 22661 24769 22695 24803
rect 22695 24769 22704 24803
rect 22836 24803 22888 24812
rect 22652 24760 22704 24769
rect 22836 24769 22844 24803
rect 22844 24769 22878 24803
rect 22878 24769 22888 24803
rect 22836 24760 22888 24769
rect 22928 24803 22980 24812
rect 22928 24769 22937 24803
rect 22937 24769 22971 24803
rect 22971 24769 22980 24803
rect 22928 24760 22980 24769
rect 38016 24896 38068 24948
rect 24676 24828 24728 24880
rect 24952 24803 25004 24812
rect 24952 24769 24961 24803
rect 24961 24769 24995 24803
rect 24995 24769 25004 24803
rect 24952 24760 25004 24769
rect 25136 24803 25188 24812
rect 25136 24769 25145 24803
rect 25145 24769 25179 24803
rect 25179 24769 25188 24803
rect 25136 24760 25188 24769
rect 25872 24828 25924 24880
rect 30472 24828 30524 24880
rect 32772 24828 32824 24880
rect 26792 24760 26844 24812
rect 29092 24760 29144 24812
rect 30564 24760 30616 24812
rect 25596 24735 25648 24744
rect 25596 24701 25605 24735
rect 25605 24701 25639 24735
rect 25639 24701 25648 24735
rect 25596 24692 25648 24701
rect 29644 24692 29696 24744
rect 28540 24624 28592 24676
rect 29828 24624 29880 24676
rect 32588 24760 32640 24812
rect 37372 24760 37424 24812
rect 34612 24692 34664 24744
rect 36176 24692 36228 24744
rect 40040 24760 40092 24812
rect 40224 24760 40276 24812
rect 15568 24599 15620 24608
rect 15568 24565 15577 24599
rect 15577 24565 15611 24599
rect 15611 24565 15620 24599
rect 15568 24556 15620 24565
rect 19340 24556 19392 24608
rect 21732 24556 21784 24608
rect 22100 24556 22152 24608
rect 28908 24556 28960 24608
rect 30380 24599 30432 24608
rect 30380 24565 30389 24599
rect 30389 24565 30423 24599
rect 30423 24565 30432 24599
rect 30380 24556 30432 24565
rect 30564 24556 30616 24608
rect 31484 24599 31536 24608
rect 31484 24565 31493 24599
rect 31493 24565 31527 24599
rect 31527 24565 31536 24599
rect 31484 24556 31536 24565
rect 38752 24599 38804 24608
rect 38752 24565 38761 24599
rect 38761 24565 38795 24599
rect 38795 24565 38804 24599
rect 38752 24556 38804 24565
rect 41236 24556 41288 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3240 24352 3292 24404
rect 5448 24352 5500 24404
rect 7932 24352 7984 24404
rect 10784 24395 10836 24404
rect 10784 24361 10793 24395
rect 10793 24361 10827 24395
rect 10827 24361 10836 24395
rect 10784 24352 10836 24361
rect 12992 24352 13044 24404
rect 14096 24395 14148 24404
rect 14096 24361 14105 24395
rect 14105 24361 14139 24395
rect 14139 24361 14148 24395
rect 14096 24352 14148 24361
rect 14924 24352 14976 24404
rect 18144 24352 18196 24404
rect 25136 24352 25188 24404
rect 9680 24148 9732 24200
rect 10600 24148 10652 24200
rect 11612 24148 11664 24200
rect 9588 24080 9640 24132
rect 11152 24123 11204 24132
rect 10232 24012 10284 24064
rect 11152 24089 11161 24123
rect 11161 24089 11195 24123
rect 11195 24089 11204 24123
rect 11152 24080 11204 24089
rect 11336 24080 11388 24132
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 12900 24191 12952 24200
rect 12900 24157 12909 24191
rect 12909 24157 12943 24191
rect 12943 24157 12952 24191
rect 12900 24148 12952 24157
rect 15016 24284 15068 24336
rect 13544 24148 13596 24200
rect 13636 24148 13688 24200
rect 14648 24148 14700 24200
rect 14832 24148 14884 24200
rect 17132 24284 17184 24336
rect 16856 24216 16908 24268
rect 18788 24284 18840 24336
rect 24952 24284 25004 24336
rect 28908 24352 28960 24404
rect 29644 24352 29696 24404
rect 29920 24352 29972 24404
rect 31116 24352 31168 24404
rect 16304 24191 16356 24200
rect 16304 24157 16313 24191
rect 16313 24157 16347 24191
rect 16347 24157 16356 24191
rect 16304 24148 16356 24157
rect 17776 24191 17828 24200
rect 17776 24157 17785 24191
rect 17785 24157 17819 24191
rect 17819 24157 17828 24191
rect 17776 24148 17828 24157
rect 18144 24148 18196 24200
rect 13728 24080 13780 24132
rect 11244 24012 11296 24064
rect 13452 24012 13504 24064
rect 14924 24080 14976 24132
rect 17132 24080 17184 24132
rect 17500 24080 17552 24132
rect 21364 24148 21416 24200
rect 21732 24191 21784 24200
rect 21732 24157 21777 24191
rect 21777 24157 21784 24191
rect 21916 24191 21968 24200
rect 21732 24148 21784 24157
rect 21916 24157 21925 24191
rect 21925 24157 21959 24191
rect 21959 24157 21968 24191
rect 21916 24148 21968 24157
rect 18788 24080 18840 24132
rect 17224 24012 17276 24064
rect 17776 24012 17828 24064
rect 18236 24012 18288 24064
rect 18512 24012 18564 24064
rect 21180 24012 21232 24064
rect 21640 24123 21692 24132
rect 21640 24089 21649 24123
rect 21649 24089 21683 24123
rect 21683 24089 21692 24123
rect 21640 24080 21692 24089
rect 25504 24191 25556 24200
rect 25504 24157 25513 24191
rect 25513 24157 25547 24191
rect 25547 24157 25556 24191
rect 25504 24148 25556 24157
rect 26792 24148 26844 24200
rect 28540 24148 28592 24200
rect 31944 24216 31996 24268
rect 30380 24148 30432 24200
rect 38752 24148 38804 24200
rect 58164 24191 58216 24200
rect 58164 24157 58173 24191
rect 58173 24157 58207 24191
rect 58207 24157 58216 24191
rect 58164 24148 58216 24157
rect 25228 24080 25280 24132
rect 25596 24080 25648 24132
rect 28632 24123 28684 24132
rect 28632 24089 28641 24123
rect 28641 24089 28675 24123
rect 28675 24089 28684 24123
rect 28632 24080 28684 24089
rect 40132 24080 40184 24132
rect 40408 24123 40460 24132
rect 26884 24055 26936 24064
rect 26884 24021 26893 24055
rect 26893 24021 26927 24055
rect 26927 24021 26936 24055
rect 26884 24012 26936 24021
rect 27252 24012 27304 24064
rect 32312 24012 32364 24064
rect 40408 24089 40417 24123
rect 40417 24089 40451 24123
rect 40451 24089 40460 24123
rect 40408 24080 40460 24089
rect 40960 24012 41012 24064
rect 41420 24055 41472 24064
rect 41420 24021 41429 24055
rect 41429 24021 41463 24055
rect 41463 24021 41472 24055
rect 41420 24012 41472 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 5264 23808 5316 23860
rect 8576 23808 8628 23860
rect 2228 23715 2280 23724
rect 2228 23681 2237 23715
rect 2237 23681 2271 23715
rect 2271 23681 2280 23715
rect 2228 23672 2280 23681
rect 3240 23672 3292 23724
rect 9588 23672 9640 23724
rect 9956 23808 10008 23860
rect 11336 23808 11388 23860
rect 12256 23808 12308 23860
rect 12440 23808 12492 23860
rect 11152 23740 11204 23792
rect 12992 23740 13044 23792
rect 6092 23604 6144 23656
rect 10324 23672 10376 23724
rect 10784 23715 10836 23724
rect 10784 23681 10793 23715
rect 10793 23681 10827 23715
rect 10827 23681 10836 23715
rect 10784 23672 10836 23681
rect 14188 23740 14240 23792
rect 21548 23808 21600 23860
rect 22192 23808 22244 23860
rect 24768 23808 24820 23860
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 29092 23851 29144 23860
rect 24952 23808 25004 23817
rect 17132 23740 17184 23792
rect 22652 23783 22704 23792
rect 13452 23715 13504 23724
rect 13452 23681 13486 23715
rect 13486 23681 13504 23715
rect 13452 23672 13504 23681
rect 17224 23715 17276 23724
rect 17224 23681 17233 23715
rect 17233 23681 17267 23715
rect 17267 23681 17276 23715
rect 17224 23672 17276 23681
rect 17776 23672 17828 23724
rect 22652 23749 22661 23783
rect 22661 23749 22695 23783
rect 22695 23749 22704 23783
rect 22652 23740 22704 23749
rect 25320 23740 25372 23792
rect 11704 23604 11756 23656
rect 14832 23604 14884 23656
rect 11796 23536 11848 23588
rect 14464 23536 14516 23588
rect 14924 23536 14976 23588
rect 18236 23715 18288 23724
rect 18236 23681 18265 23715
rect 18265 23681 18288 23715
rect 22376 23715 22428 23724
rect 18236 23672 18288 23681
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 22560 23715 22612 23724
rect 22560 23681 22567 23715
rect 22567 23681 22612 23715
rect 22560 23672 22612 23681
rect 18512 23604 18564 23656
rect 19340 23604 19392 23656
rect 21364 23604 21416 23656
rect 24952 23672 25004 23724
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 29092 23817 29101 23851
rect 29101 23817 29135 23851
rect 29135 23817 29144 23851
rect 29092 23808 29144 23817
rect 30840 23808 30892 23860
rect 33968 23808 34020 23860
rect 31576 23740 31628 23792
rect 32956 23783 33008 23792
rect 24676 23604 24728 23656
rect 28816 23672 28868 23724
rect 28264 23604 28316 23656
rect 29552 23715 29604 23724
rect 32956 23749 32965 23783
rect 32965 23749 32999 23783
rect 32999 23749 33008 23783
rect 32956 23740 33008 23749
rect 33324 23740 33376 23792
rect 36084 23740 36136 23792
rect 41236 23808 41288 23860
rect 29552 23681 29566 23715
rect 29566 23681 29600 23715
rect 29600 23681 29604 23715
rect 29552 23672 29604 23681
rect 2504 23468 2556 23520
rect 9496 23511 9548 23520
rect 9496 23477 9505 23511
rect 9505 23477 9539 23511
rect 9539 23477 9548 23511
rect 9496 23468 9548 23477
rect 9588 23468 9640 23520
rect 12440 23468 12492 23520
rect 12532 23468 12584 23520
rect 13544 23468 13596 23520
rect 15384 23468 15436 23520
rect 16304 23468 16356 23520
rect 18144 23536 18196 23588
rect 21456 23536 21508 23588
rect 18512 23511 18564 23520
rect 18512 23477 18521 23511
rect 18521 23477 18555 23511
rect 18555 23477 18564 23511
rect 18512 23468 18564 23477
rect 23204 23468 23256 23520
rect 26148 23511 26200 23520
rect 26148 23477 26157 23511
rect 26157 23477 26191 23511
rect 26191 23477 26200 23511
rect 26148 23468 26200 23477
rect 28816 23468 28868 23520
rect 29460 23536 29512 23588
rect 29828 23604 29880 23656
rect 35624 23672 35676 23724
rect 35808 23715 35860 23724
rect 35808 23681 35817 23715
rect 35817 23681 35851 23715
rect 35851 23681 35860 23715
rect 35808 23672 35860 23681
rect 35992 23715 36044 23724
rect 35992 23681 36001 23715
rect 36001 23681 36035 23715
rect 36035 23681 36044 23715
rect 35992 23672 36044 23681
rect 36176 23715 36228 23724
rect 36176 23681 36185 23715
rect 36185 23681 36219 23715
rect 36219 23681 36228 23715
rect 36176 23672 36228 23681
rect 40040 23672 40092 23724
rect 34244 23604 34296 23656
rect 37924 23647 37976 23656
rect 37924 23613 37933 23647
rect 37933 23613 37967 23647
rect 37967 23613 37976 23647
rect 37924 23604 37976 23613
rect 41052 23715 41104 23724
rect 41052 23681 41066 23715
rect 41066 23681 41100 23715
rect 41100 23681 41104 23715
rect 41052 23672 41104 23681
rect 38384 23536 38436 23588
rect 40960 23536 41012 23588
rect 41052 23536 41104 23588
rect 30472 23468 30524 23520
rect 32496 23511 32548 23520
rect 32496 23477 32505 23511
rect 32505 23477 32539 23511
rect 32539 23477 32548 23511
rect 32496 23468 32548 23477
rect 32680 23511 32732 23520
rect 32680 23477 32689 23511
rect 32689 23477 32723 23511
rect 32723 23477 32732 23511
rect 32680 23468 32732 23477
rect 32772 23468 32824 23520
rect 33508 23468 33560 23520
rect 35900 23468 35952 23520
rect 40408 23468 40460 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2964 23264 3016 23316
rect 3976 23264 4028 23316
rect 18236 23307 18288 23316
rect 18236 23273 18245 23307
rect 18245 23273 18279 23307
rect 18279 23273 18288 23307
rect 18236 23264 18288 23273
rect 23112 23264 23164 23316
rect 2688 23103 2740 23112
rect 2688 23069 2697 23103
rect 2697 23069 2731 23103
rect 2731 23069 2740 23103
rect 2688 23060 2740 23069
rect 2780 23103 2832 23112
rect 2780 23069 2789 23103
rect 2789 23069 2823 23103
rect 2823 23069 2832 23103
rect 2780 23060 2832 23069
rect 2964 23103 3016 23112
rect 2964 23069 2973 23103
rect 2973 23069 3007 23103
rect 3007 23069 3016 23103
rect 7380 23103 7432 23112
rect 2964 23060 3016 23069
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 2228 22992 2280 23044
rect 4620 22992 4672 23044
rect 2688 22924 2740 22976
rect 7656 22924 7708 22976
rect 9680 23060 9732 23112
rect 11244 23103 11296 23112
rect 11244 23069 11278 23103
rect 11278 23069 11296 23103
rect 11244 23060 11296 23069
rect 11520 23060 11572 23112
rect 14832 23103 14884 23112
rect 14832 23069 14841 23103
rect 14841 23069 14875 23103
rect 14875 23069 14884 23103
rect 14832 23060 14884 23069
rect 9496 22992 9548 23044
rect 11888 22992 11940 23044
rect 14372 23035 14424 23044
rect 14372 23001 14381 23035
rect 14381 23001 14415 23035
rect 14415 23001 14424 23035
rect 14372 22992 14424 23001
rect 10140 22924 10192 22976
rect 10784 22924 10836 22976
rect 11704 22924 11756 22976
rect 14924 22924 14976 22976
rect 15568 22992 15620 23044
rect 15936 23060 15988 23112
rect 17592 23128 17644 23180
rect 23112 23128 23164 23180
rect 22744 23060 22796 23112
rect 23204 23103 23256 23112
rect 23204 23069 23213 23103
rect 23213 23069 23247 23103
rect 23247 23069 23256 23103
rect 23204 23060 23256 23069
rect 29552 23264 29604 23316
rect 36084 23196 36136 23248
rect 25504 23128 25556 23180
rect 34152 23171 34204 23180
rect 34152 23137 34161 23171
rect 34161 23137 34195 23171
rect 34195 23137 34204 23171
rect 34152 23128 34204 23137
rect 23388 23060 23440 23112
rect 24676 23103 24728 23112
rect 24676 23069 24685 23103
rect 24685 23069 24719 23103
rect 24719 23069 24728 23103
rect 24676 23060 24728 23069
rect 26148 23103 26200 23112
rect 26148 23069 26182 23103
rect 26182 23069 26200 23103
rect 26148 23060 26200 23069
rect 35808 23128 35860 23180
rect 39120 23264 39172 23316
rect 40224 23264 40276 23316
rect 37188 23060 37240 23112
rect 37924 23060 37976 23112
rect 38200 23103 38252 23112
rect 38200 23069 38209 23103
rect 38209 23069 38243 23103
rect 38243 23069 38252 23103
rect 38200 23060 38252 23069
rect 38384 23103 38436 23112
rect 38384 23069 38393 23103
rect 38393 23069 38427 23103
rect 38427 23069 38436 23103
rect 40408 23103 40460 23112
rect 38384 23060 38436 23069
rect 40408 23069 40431 23103
rect 40431 23069 40460 23103
rect 40408 23060 40460 23069
rect 41420 23128 41472 23180
rect 20444 23035 20496 23044
rect 20444 23001 20453 23035
rect 20453 23001 20487 23035
rect 20487 23001 20496 23035
rect 20444 22992 20496 23001
rect 15292 22924 15344 22976
rect 17408 22924 17460 22976
rect 20536 22924 20588 22976
rect 22284 22967 22336 22976
rect 22284 22933 22293 22967
rect 22293 22933 22327 22967
rect 22327 22933 22336 22967
rect 22284 22924 22336 22933
rect 25320 22992 25372 23044
rect 28448 22992 28500 23044
rect 33416 22992 33468 23044
rect 27620 22924 27672 22976
rect 29368 22924 29420 22976
rect 32312 22924 32364 22976
rect 32864 22924 32916 22976
rect 34152 22924 34204 22976
rect 35992 22992 36044 23044
rect 41052 23060 41104 23112
rect 40960 22992 41012 23044
rect 38752 22924 38804 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 2780 22720 2832 22772
rect 3792 22763 3844 22772
rect 3792 22729 3801 22763
rect 3801 22729 3835 22763
rect 3835 22729 3844 22763
rect 3792 22720 3844 22729
rect 9220 22720 9272 22772
rect 11060 22720 11112 22772
rect 15936 22763 15988 22772
rect 2228 22652 2280 22704
rect 2596 22652 2648 22704
rect 2688 22627 2740 22636
rect 2688 22593 2722 22627
rect 2722 22593 2740 22627
rect 2688 22584 2740 22593
rect 4620 22627 4672 22636
rect 4620 22593 4629 22627
rect 4629 22593 4663 22627
rect 4663 22593 4672 22627
rect 8668 22652 8720 22704
rect 13268 22652 13320 22704
rect 14464 22695 14516 22704
rect 14464 22661 14473 22695
rect 14473 22661 14507 22695
rect 14507 22661 14516 22695
rect 14464 22652 14516 22661
rect 4620 22584 4672 22593
rect 4712 22516 4764 22568
rect 3792 22380 3844 22432
rect 4620 22380 4672 22432
rect 6368 22380 6420 22432
rect 6828 22627 6880 22636
rect 6828 22593 6862 22627
rect 6862 22593 6880 22627
rect 6828 22584 6880 22593
rect 9036 22584 9088 22636
rect 10048 22584 10100 22636
rect 7656 22516 7708 22568
rect 8024 22516 8076 22568
rect 8944 22516 8996 22568
rect 12164 22584 12216 22636
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 15936 22729 15945 22763
rect 15945 22729 15979 22763
rect 15979 22729 15988 22763
rect 15936 22720 15988 22729
rect 14188 22516 14240 22568
rect 14924 22516 14976 22568
rect 18512 22652 18564 22704
rect 19340 22763 19392 22772
rect 19340 22729 19349 22763
rect 19349 22729 19383 22763
rect 19383 22729 19392 22763
rect 19340 22720 19392 22729
rect 20628 22720 20680 22772
rect 23112 22720 23164 22772
rect 25228 22763 25280 22772
rect 23296 22652 23348 22704
rect 25228 22729 25237 22763
rect 25237 22729 25271 22763
rect 25271 22729 25280 22763
rect 25228 22720 25280 22729
rect 26700 22652 26752 22704
rect 17408 22584 17460 22636
rect 18604 22584 18656 22636
rect 14832 22448 14884 22500
rect 8024 22380 8076 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 14556 22380 14608 22432
rect 15752 22380 15804 22432
rect 19340 22380 19392 22432
rect 20812 22584 20864 22636
rect 21180 22627 21232 22636
rect 21180 22593 21189 22627
rect 21189 22593 21223 22627
rect 21223 22593 21232 22627
rect 21180 22584 21232 22593
rect 25044 22627 25096 22636
rect 25044 22593 25053 22627
rect 25053 22593 25087 22627
rect 25087 22593 25096 22627
rect 25044 22584 25096 22593
rect 32772 22720 32824 22772
rect 33416 22763 33468 22772
rect 33416 22729 33425 22763
rect 33425 22729 33459 22763
rect 33459 22729 33468 22763
rect 33416 22720 33468 22729
rect 35624 22763 35676 22772
rect 35624 22729 35633 22763
rect 35633 22729 35667 22763
rect 35667 22729 35676 22763
rect 35624 22720 35676 22729
rect 38200 22720 38252 22772
rect 40316 22720 40368 22772
rect 27620 22652 27672 22704
rect 28448 22695 28500 22704
rect 28448 22661 28457 22695
rect 28457 22661 28491 22695
rect 28491 22661 28500 22695
rect 28448 22652 28500 22661
rect 29920 22652 29972 22704
rect 31208 22695 31260 22704
rect 31208 22661 31217 22695
rect 31217 22661 31251 22695
rect 31251 22661 31260 22695
rect 31208 22652 31260 22661
rect 32312 22652 32364 22704
rect 33876 22695 33928 22704
rect 33876 22661 33885 22695
rect 33885 22661 33919 22695
rect 33919 22661 33928 22695
rect 33876 22652 33928 22661
rect 35900 22695 35952 22704
rect 35900 22661 35909 22695
rect 35909 22661 35943 22695
rect 35943 22661 35952 22695
rect 35900 22652 35952 22661
rect 36084 22652 36136 22704
rect 40132 22652 40184 22704
rect 40592 22652 40644 22704
rect 28632 22627 28684 22636
rect 28632 22593 28641 22627
rect 28641 22593 28675 22627
rect 28675 22593 28684 22627
rect 28632 22584 28684 22593
rect 29736 22584 29788 22636
rect 31392 22627 31444 22636
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 32588 22584 32640 22636
rect 32496 22516 32548 22568
rect 31760 22448 31812 22500
rect 34152 22627 34204 22636
rect 32956 22448 33008 22500
rect 33048 22448 33100 22500
rect 34152 22593 34161 22627
rect 34161 22593 34195 22627
rect 34195 22593 34204 22627
rect 34152 22584 34204 22593
rect 35808 22627 35860 22636
rect 35808 22593 35817 22627
rect 35817 22593 35851 22627
rect 35851 22593 35860 22627
rect 35808 22584 35860 22593
rect 35992 22627 36044 22636
rect 35992 22593 36001 22627
rect 36001 22593 36035 22627
rect 36035 22593 36044 22627
rect 35992 22584 36044 22593
rect 37096 22584 37148 22636
rect 37372 22584 37424 22636
rect 38108 22584 38160 22636
rect 38292 22584 38344 22636
rect 33784 22516 33836 22568
rect 36268 22516 36320 22568
rect 34336 22491 34388 22500
rect 20904 22380 20956 22432
rect 20996 22423 21048 22432
rect 20996 22389 21005 22423
rect 21005 22389 21039 22423
rect 21039 22389 21048 22423
rect 20996 22380 21048 22389
rect 25688 22380 25740 22432
rect 28356 22380 28408 22432
rect 30932 22380 30984 22432
rect 31484 22380 31536 22432
rect 33876 22423 33928 22432
rect 33876 22389 33885 22423
rect 33885 22389 33919 22423
rect 33919 22389 33928 22423
rect 33876 22380 33928 22389
rect 34336 22457 34345 22491
rect 34345 22457 34379 22491
rect 34379 22457 34388 22491
rect 34336 22448 34388 22457
rect 41236 22448 41288 22500
rect 58164 22491 58216 22500
rect 58164 22457 58173 22491
rect 58173 22457 58207 22491
rect 58207 22457 58216 22491
rect 58164 22448 58216 22457
rect 38936 22380 38988 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 6828 22219 6880 22228
rect 3240 22176 3292 22185
rect 6828 22185 6837 22219
rect 6837 22185 6871 22219
rect 6871 22185 6880 22219
rect 6828 22176 6880 22185
rect 8116 22219 8168 22228
rect 8116 22185 8125 22219
rect 8125 22185 8159 22219
rect 8159 22185 8168 22219
rect 8116 22176 8168 22185
rect 14924 22219 14976 22228
rect 14924 22185 14933 22219
rect 14933 22185 14967 22219
rect 14967 22185 14976 22219
rect 14924 22176 14976 22185
rect 21272 22176 21324 22228
rect 31116 22176 31168 22228
rect 31484 22176 31536 22228
rect 33876 22176 33928 22228
rect 37832 22176 37884 22228
rect 38292 22176 38344 22228
rect 11888 22108 11940 22160
rect 16948 22108 17000 22160
rect 18236 22108 18288 22160
rect 22468 22108 22520 22160
rect 15752 22083 15804 22092
rect 2688 21972 2740 22024
rect 5172 21972 5224 22024
rect 6092 21972 6144 22024
rect 6363 22015 6415 22024
rect 6363 21981 6372 22015
rect 6372 21981 6406 22015
rect 6406 21981 6415 22015
rect 6363 21972 6415 21981
rect 7656 22015 7708 22024
rect 2136 21947 2188 21956
rect 2136 21913 2170 21947
rect 2170 21913 2188 21947
rect 2136 21904 2188 21913
rect 3608 21904 3660 21956
rect 6000 21904 6052 21956
rect 7656 21981 7665 22015
rect 7665 21981 7699 22015
rect 7699 21981 7708 22015
rect 7656 21972 7708 21981
rect 9220 21972 9272 22024
rect 10324 21972 10376 22024
rect 15752 22049 15761 22083
rect 15761 22049 15795 22083
rect 15795 22049 15804 22083
rect 15752 22040 15804 22049
rect 11704 22015 11756 22024
rect 11704 21981 11713 22015
rect 11713 21981 11747 22015
rect 11747 21981 11756 22015
rect 11704 21972 11756 21981
rect 12440 21972 12492 22024
rect 13360 21972 13412 22024
rect 14832 21972 14884 22024
rect 15384 21972 15436 22024
rect 4712 21836 4764 21888
rect 5264 21836 5316 21888
rect 5908 21836 5960 21888
rect 7748 21904 7800 21956
rect 10048 21947 10100 21956
rect 10048 21913 10057 21947
rect 10057 21913 10091 21947
rect 10091 21913 10100 21947
rect 10048 21904 10100 21913
rect 11612 21947 11664 21956
rect 11612 21913 11621 21947
rect 11621 21913 11655 21947
rect 11655 21913 11664 21947
rect 11612 21904 11664 21913
rect 12164 21904 12216 21956
rect 17132 21972 17184 22024
rect 17684 21972 17736 22024
rect 21088 22015 21140 22024
rect 21088 21981 21097 22015
rect 21097 21981 21131 22015
rect 21131 21981 21140 22015
rect 21088 21972 21140 21981
rect 22100 21972 22152 22024
rect 22192 21972 22244 22024
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 22928 22108 22980 22160
rect 23388 22108 23440 22160
rect 31392 22108 31444 22160
rect 26884 22040 26936 22092
rect 22468 21904 22520 21956
rect 27436 21972 27488 22024
rect 31852 21972 31904 22024
rect 33140 22108 33192 22160
rect 32772 22015 32824 22024
rect 32772 21981 32781 22015
rect 32781 21981 32815 22015
rect 32815 21981 32824 22015
rect 32772 21972 32824 21981
rect 33692 22040 33744 22092
rect 33140 22015 33192 22024
rect 33140 21981 33149 22015
rect 33149 21981 33183 22015
rect 33183 21981 33192 22015
rect 33140 21972 33192 21981
rect 38844 21972 38896 22024
rect 27896 21947 27948 21956
rect 27896 21913 27930 21947
rect 27930 21913 27948 21947
rect 27896 21904 27948 21913
rect 28724 21904 28776 21956
rect 30840 21904 30892 21956
rect 31208 21904 31260 21956
rect 38476 21904 38528 21956
rect 8116 21836 8168 21888
rect 9036 21879 9088 21888
rect 9036 21845 9045 21879
rect 9045 21845 9079 21879
rect 9079 21845 9088 21879
rect 9036 21836 9088 21845
rect 10232 21836 10284 21888
rect 10968 21836 11020 21888
rect 12072 21836 12124 21888
rect 13544 21836 13596 21888
rect 15384 21879 15436 21888
rect 15384 21845 15393 21879
rect 15393 21845 15427 21879
rect 15427 21845 15436 21879
rect 15384 21836 15436 21845
rect 15844 21836 15896 21888
rect 21180 21836 21232 21888
rect 22652 21836 22704 21888
rect 23112 21836 23164 21888
rect 23296 21836 23348 21888
rect 28448 21836 28500 21888
rect 32680 21836 32732 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2136 21675 2188 21684
rect 2136 21641 2145 21675
rect 2145 21641 2179 21675
rect 2179 21641 2188 21675
rect 2136 21632 2188 21641
rect 3608 21675 3660 21684
rect 3608 21641 3617 21675
rect 3617 21641 3651 21675
rect 3651 21641 3660 21675
rect 3608 21632 3660 21641
rect 3056 21564 3108 21616
rect 2596 21539 2648 21548
rect 2596 21505 2605 21539
rect 2605 21505 2639 21539
rect 2639 21505 2648 21539
rect 2596 21496 2648 21505
rect 3884 21539 3936 21548
rect 3884 21505 3893 21539
rect 3893 21505 3927 21539
rect 3927 21505 3936 21539
rect 3884 21496 3936 21505
rect 4620 21564 4672 21616
rect 6000 21632 6052 21684
rect 7380 21632 7432 21684
rect 10048 21632 10100 21684
rect 11612 21632 11664 21684
rect 14372 21632 14424 21684
rect 15568 21632 15620 21684
rect 5172 21539 5224 21548
rect 2964 21428 3016 21480
rect 5172 21505 5181 21539
rect 5181 21505 5215 21539
rect 5215 21505 5224 21539
rect 5172 21496 5224 21505
rect 10140 21607 10192 21616
rect 10140 21573 10149 21607
rect 10149 21573 10183 21607
rect 10183 21573 10192 21607
rect 10140 21564 10192 21573
rect 14464 21564 14516 21616
rect 21088 21632 21140 21684
rect 33508 21632 33560 21684
rect 38476 21675 38528 21684
rect 38476 21641 38485 21675
rect 38485 21641 38519 21675
rect 38519 21641 38528 21675
rect 38476 21632 38528 21641
rect 21640 21564 21692 21616
rect 23112 21564 23164 21616
rect 25044 21564 25096 21616
rect 27896 21607 27948 21616
rect 27896 21573 27905 21607
rect 27905 21573 27939 21607
rect 27939 21573 27948 21607
rect 27896 21564 27948 21573
rect 28448 21564 28500 21616
rect 32864 21564 32916 21616
rect 5724 21496 5776 21548
rect 5908 21428 5960 21480
rect 2780 21360 2832 21412
rect 5264 21360 5316 21412
rect 10048 21539 10100 21548
rect 10048 21505 10057 21539
rect 10057 21505 10091 21539
rect 10091 21505 10100 21539
rect 10048 21496 10100 21505
rect 10324 21496 10376 21548
rect 12440 21496 12492 21548
rect 15752 21539 15804 21548
rect 15752 21505 15761 21539
rect 15761 21505 15795 21539
rect 15795 21505 15804 21539
rect 15752 21496 15804 21505
rect 6368 21471 6420 21480
rect 6368 21437 6377 21471
rect 6377 21437 6411 21471
rect 6411 21437 6420 21471
rect 6368 21428 6420 21437
rect 9036 21428 9088 21480
rect 7748 21403 7800 21412
rect 7748 21369 7757 21403
rect 7757 21369 7791 21403
rect 7791 21369 7800 21403
rect 7748 21360 7800 21369
rect 11060 21360 11112 21412
rect 13544 21428 13596 21480
rect 15384 21360 15436 21412
rect 16948 21428 17000 21480
rect 17224 21539 17276 21548
rect 17224 21505 17233 21539
rect 17233 21505 17267 21539
rect 17267 21505 17276 21539
rect 17224 21496 17276 21505
rect 17776 21496 17828 21548
rect 22560 21496 22612 21548
rect 24676 21496 24728 21548
rect 27712 21496 27764 21548
rect 28264 21539 28316 21548
rect 28264 21505 28273 21539
rect 28273 21505 28307 21539
rect 28307 21505 28316 21539
rect 28264 21496 28316 21505
rect 34796 21564 34848 21616
rect 20076 21428 20128 21480
rect 22652 21428 22704 21480
rect 21824 21360 21876 21412
rect 10600 21292 10652 21344
rect 16764 21335 16816 21344
rect 16764 21301 16773 21335
rect 16773 21301 16807 21335
rect 16807 21301 16816 21335
rect 16764 21292 16816 21301
rect 22100 21292 22152 21344
rect 26424 21360 26476 21412
rect 29552 21403 29604 21412
rect 29552 21369 29561 21403
rect 29561 21369 29595 21403
rect 29595 21369 29604 21403
rect 29552 21360 29604 21369
rect 33324 21496 33376 21548
rect 30104 21428 30156 21480
rect 32956 21428 33008 21480
rect 37280 21360 37332 21412
rect 23020 21292 23072 21344
rect 24676 21292 24728 21344
rect 29828 21335 29880 21344
rect 29828 21301 29837 21335
rect 29837 21301 29871 21335
rect 29871 21301 29880 21335
rect 29828 21292 29880 21301
rect 32956 21292 33008 21344
rect 38660 21496 38712 21548
rect 38936 21539 38988 21548
rect 38936 21505 38945 21539
rect 38945 21505 38979 21539
rect 38979 21505 38988 21539
rect 38936 21496 38988 21505
rect 39764 21496 39816 21548
rect 40040 21428 40092 21480
rect 40868 21428 40920 21480
rect 58164 21335 58216 21344
rect 58164 21301 58173 21335
rect 58173 21301 58207 21335
rect 58207 21301 58216 21335
rect 58164 21292 58216 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 5724 21088 5776 21140
rect 6000 21088 6052 21140
rect 8208 21088 8260 21140
rect 13084 21088 13136 21140
rect 17960 21088 18012 21140
rect 18880 21088 18932 21140
rect 20168 21088 20220 21140
rect 11152 21020 11204 21072
rect 12256 21020 12308 21072
rect 17500 21020 17552 21072
rect 21364 21088 21416 21140
rect 21824 21131 21876 21140
rect 21824 21097 21833 21131
rect 21833 21097 21867 21131
rect 21867 21097 21876 21131
rect 21824 21088 21876 21097
rect 13636 20952 13688 21004
rect 14464 20884 14516 20936
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 15568 20927 15620 20936
rect 15568 20893 15577 20927
rect 15577 20893 15611 20927
rect 15611 20893 15620 20927
rect 15568 20884 15620 20893
rect 2780 20816 2832 20868
rect 4620 20816 4672 20868
rect 6184 20816 6236 20868
rect 12716 20859 12768 20868
rect 3884 20748 3936 20800
rect 5632 20748 5684 20800
rect 6552 20748 6604 20800
rect 8484 20748 8536 20800
rect 12716 20825 12725 20859
rect 12725 20825 12759 20859
rect 12759 20825 12768 20859
rect 12716 20816 12768 20825
rect 11612 20748 11664 20800
rect 15660 20859 15712 20868
rect 15660 20825 15669 20859
rect 15669 20825 15703 20859
rect 15703 20825 15712 20859
rect 15660 20816 15712 20825
rect 12992 20748 13044 20800
rect 17408 20884 17460 20936
rect 16764 20816 16816 20868
rect 20536 21020 20588 21072
rect 17776 20791 17828 20800
rect 17776 20757 17785 20791
rect 17785 20757 17819 20791
rect 17819 20757 17828 20791
rect 17776 20748 17828 20757
rect 20168 20859 20220 20868
rect 20168 20825 20177 20859
rect 20177 20825 20211 20859
rect 20211 20825 20220 20859
rect 20168 20816 20220 20825
rect 20996 20884 21048 20936
rect 22100 20884 22152 20936
rect 22560 20927 22612 20936
rect 22560 20893 22569 20927
rect 22569 20893 22603 20927
rect 22603 20893 22612 20927
rect 22560 20884 22612 20893
rect 22836 21088 22888 21140
rect 23112 21088 23164 21140
rect 27712 21088 27764 21140
rect 32956 21088 33008 21140
rect 30196 20952 30248 21004
rect 20628 20816 20680 20868
rect 21088 20859 21140 20868
rect 21088 20825 21097 20859
rect 21097 20825 21131 20859
rect 21131 20825 21140 20859
rect 21088 20816 21140 20825
rect 23020 20884 23072 20936
rect 29276 20884 29328 20936
rect 40224 20884 40276 20936
rect 22928 20816 22980 20868
rect 20260 20748 20312 20800
rect 23940 20816 23992 20868
rect 25044 20816 25096 20868
rect 27436 20859 27488 20868
rect 24400 20748 24452 20800
rect 27436 20825 27445 20859
rect 27445 20825 27479 20859
rect 27479 20825 27488 20859
rect 27436 20816 27488 20825
rect 30840 20816 30892 20868
rect 40500 20816 40552 20868
rect 40684 20816 40736 20868
rect 27712 20748 27764 20800
rect 28172 20748 28224 20800
rect 28540 20748 28592 20800
rect 37464 20791 37516 20800
rect 37464 20757 37473 20791
rect 37473 20757 37507 20791
rect 37507 20757 37516 20791
rect 37464 20748 37516 20757
rect 41144 20748 41196 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 5816 20476 5868 20528
rect 8392 20544 8444 20596
rect 12532 20544 12584 20596
rect 13636 20587 13688 20596
rect 13636 20553 13645 20587
rect 13645 20553 13679 20587
rect 13679 20553 13688 20587
rect 13636 20544 13688 20553
rect 17224 20544 17276 20596
rect 11520 20476 11572 20528
rect 17776 20476 17828 20528
rect 6552 20408 6604 20460
rect 12532 20451 12584 20460
rect 12532 20417 12566 20451
rect 12566 20417 12584 20451
rect 6828 20340 6880 20392
rect 12532 20408 12584 20417
rect 12808 20408 12860 20460
rect 15292 20408 15344 20460
rect 15752 20408 15804 20460
rect 16580 20408 16632 20460
rect 17592 20408 17644 20460
rect 14096 20383 14148 20392
rect 14096 20349 14105 20383
rect 14105 20349 14139 20383
rect 14139 20349 14148 20383
rect 14096 20340 14148 20349
rect 15936 20340 15988 20392
rect 16948 20272 17000 20324
rect 12440 20204 12492 20256
rect 17960 20247 18012 20256
rect 17960 20213 17969 20247
rect 17969 20213 18003 20247
rect 18003 20213 18012 20247
rect 17960 20204 18012 20213
rect 18144 20247 18196 20256
rect 18144 20213 18153 20247
rect 18153 20213 18187 20247
rect 18187 20213 18196 20247
rect 18144 20204 18196 20213
rect 19616 20519 19668 20528
rect 19616 20485 19625 20519
rect 19625 20485 19659 20519
rect 19659 20485 19668 20519
rect 20168 20544 20220 20596
rect 19616 20476 19668 20485
rect 20260 20476 20312 20528
rect 19524 20451 19576 20460
rect 19524 20417 19533 20451
rect 19533 20417 19567 20451
rect 19567 20417 19576 20451
rect 19800 20451 19852 20460
rect 19524 20408 19576 20417
rect 19800 20417 19808 20451
rect 19808 20417 19842 20451
rect 19842 20417 19852 20451
rect 19800 20408 19852 20417
rect 20076 20408 20128 20460
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 20536 20476 20588 20528
rect 20720 20519 20772 20528
rect 20720 20485 20729 20519
rect 20729 20485 20763 20519
rect 20763 20485 20772 20519
rect 20720 20476 20772 20485
rect 22100 20519 22152 20528
rect 22100 20485 22109 20519
rect 22109 20485 22143 20519
rect 22143 20485 22152 20519
rect 27804 20544 27856 20596
rect 28816 20544 28868 20596
rect 29552 20544 29604 20596
rect 29828 20587 29880 20596
rect 29828 20553 29837 20587
rect 29837 20553 29871 20587
rect 29871 20553 29880 20587
rect 29828 20544 29880 20553
rect 37280 20587 37332 20596
rect 30748 20519 30800 20528
rect 22100 20476 22152 20485
rect 30748 20485 30757 20519
rect 30757 20485 30791 20519
rect 30791 20485 30800 20519
rect 30748 20476 30800 20485
rect 20628 20451 20680 20460
rect 20628 20417 20637 20451
rect 20637 20417 20671 20451
rect 20671 20417 20680 20451
rect 20628 20408 20680 20417
rect 20260 20340 20312 20392
rect 21088 20408 21140 20460
rect 23020 20451 23072 20460
rect 23020 20417 23029 20451
rect 23029 20417 23063 20451
rect 23063 20417 23072 20451
rect 23020 20408 23072 20417
rect 23296 20451 23348 20460
rect 23296 20417 23330 20451
rect 23330 20417 23348 20451
rect 23296 20408 23348 20417
rect 25780 20408 25832 20460
rect 27528 20408 27580 20460
rect 27896 20408 27948 20460
rect 28540 20408 28592 20460
rect 29000 20408 29052 20460
rect 29460 20451 29512 20460
rect 29460 20417 29469 20451
rect 29469 20417 29503 20451
rect 29503 20417 29512 20451
rect 29460 20408 29512 20417
rect 19432 20272 19484 20324
rect 19524 20272 19576 20324
rect 20168 20204 20220 20256
rect 20996 20247 21048 20256
rect 20996 20213 21005 20247
rect 21005 20213 21039 20247
rect 21039 20213 21048 20247
rect 20996 20204 21048 20213
rect 24400 20247 24452 20256
rect 24400 20213 24409 20247
rect 24409 20213 24443 20247
rect 24443 20213 24452 20247
rect 24400 20204 24452 20213
rect 27436 20272 27488 20324
rect 29644 20451 29696 20460
rect 29644 20417 29653 20451
rect 29653 20417 29687 20451
rect 29687 20417 29696 20451
rect 29644 20408 29696 20417
rect 32588 20451 32640 20460
rect 32588 20417 32597 20451
rect 32597 20417 32631 20451
rect 32631 20417 32640 20451
rect 32588 20408 32640 20417
rect 32772 20451 32824 20460
rect 32772 20417 32781 20451
rect 32781 20417 32815 20451
rect 32815 20417 32824 20451
rect 32772 20408 32824 20417
rect 33140 20476 33192 20528
rect 37280 20553 37289 20587
rect 37289 20553 37323 20587
rect 37323 20553 37332 20587
rect 37280 20544 37332 20553
rect 37372 20476 37424 20528
rect 37648 20519 37700 20528
rect 37648 20485 37657 20519
rect 37657 20485 37691 20519
rect 37691 20485 37700 20519
rect 37648 20476 37700 20485
rect 32956 20451 33008 20460
rect 32956 20417 32965 20451
rect 32965 20417 32999 20451
rect 32999 20417 33008 20451
rect 32956 20408 33008 20417
rect 37280 20408 37332 20460
rect 37556 20451 37608 20460
rect 37556 20417 37565 20451
rect 37565 20417 37599 20451
rect 37599 20417 37608 20451
rect 37832 20451 37884 20460
rect 37556 20408 37608 20417
rect 37832 20417 37841 20451
rect 37841 20417 37875 20451
rect 37875 20417 37884 20451
rect 37832 20408 37884 20417
rect 30564 20383 30616 20392
rect 30564 20349 30573 20383
rect 30573 20349 30607 20383
rect 30607 20349 30616 20383
rect 30564 20340 30616 20349
rect 32772 20272 32824 20324
rect 27068 20204 27120 20256
rect 30472 20247 30524 20256
rect 30472 20213 30481 20247
rect 30481 20213 30515 20247
rect 30515 20213 30524 20247
rect 30472 20204 30524 20213
rect 33140 20204 33192 20256
rect 34152 20204 34204 20256
rect 38752 20340 38804 20392
rect 40500 20272 40552 20324
rect 40960 20544 41012 20596
rect 40957 20408 41009 20460
rect 41236 20340 41288 20392
rect 41052 20272 41104 20324
rect 40224 20247 40276 20256
rect 40224 20213 40233 20247
rect 40233 20213 40267 20247
rect 40267 20213 40276 20247
rect 40224 20204 40276 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6276 20000 6328 20052
rect 8852 20000 8904 20052
rect 11152 20000 11204 20052
rect 12532 20000 12584 20052
rect 15200 20043 15252 20052
rect 15200 20009 15209 20043
rect 15209 20009 15243 20043
rect 15243 20009 15252 20043
rect 15200 20000 15252 20009
rect 15752 20000 15804 20052
rect 19616 20000 19668 20052
rect 20628 20000 20680 20052
rect 22100 20000 22152 20052
rect 22928 20000 22980 20052
rect 25780 20043 25832 20052
rect 25780 20009 25789 20043
rect 25789 20009 25823 20043
rect 25823 20009 25832 20043
rect 25780 20000 25832 20009
rect 27712 20043 27764 20052
rect 27712 20009 27721 20043
rect 27721 20009 27755 20043
rect 27755 20009 27764 20043
rect 27712 20000 27764 20009
rect 30472 20000 30524 20052
rect 32864 20000 32916 20052
rect 38660 20000 38712 20052
rect 12808 19932 12860 19984
rect 4620 19907 4672 19916
rect 4620 19873 4629 19907
rect 4629 19873 4663 19907
rect 4663 19873 4672 19907
rect 4620 19864 4672 19873
rect 5448 19864 5500 19916
rect 2504 19839 2556 19848
rect 2504 19805 2513 19839
rect 2513 19805 2547 19839
rect 2547 19805 2556 19839
rect 2504 19796 2556 19805
rect 6552 19796 6604 19848
rect 5080 19728 5132 19780
rect 5356 19728 5408 19780
rect 12256 19796 12308 19848
rect 9864 19771 9916 19780
rect 9864 19737 9873 19771
rect 9873 19737 9907 19771
rect 9907 19737 9916 19771
rect 9864 19728 9916 19737
rect 12992 19796 13044 19848
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 16580 19932 16632 19984
rect 15200 19907 15252 19916
rect 15200 19873 15209 19907
rect 15209 19873 15243 19907
rect 15243 19873 15252 19907
rect 15200 19864 15252 19873
rect 13084 19796 13136 19805
rect 17500 19796 17552 19848
rect 22192 19796 22244 19848
rect 26056 19839 26108 19848
rect 26056 19805 26065 19839
rect 26065 19805 26099 19839
rect 26099 19805 26108 19839
rect 26056 19796 26108 19805
rect 28264 19932 28316 19984
rect 14188 19728 14240 19780
rect 19984 19728 20036 19780
rect 24584 19728 24636 19780
rect 26516 19796 26568 19848
rect 27068 19839 27120 19848
rect 27068 19805 27077 19839
rect 27077 19805 27111 19839
rect 27111 19805 27120 19839
rect 27068 19796 27120 19805
rect 26884 19728 26936 19780
rect 28632 19864 28684 19916
rect 36268 19907 36320 19916
rect 36268 19873 36277 19907
rect 36277 19873 36311 19907
rect 36311 19873 36320 19907
rect 36268 19864 36320 19873
rect 27620 19796 27672 19848
rect 28908 19796 28960 19848
rect 29644 19796 29696 19848
rect 30012 19796 30064 19848
rect 31392 19796 31444 19848
rect 32772 19796 32824 19848
rect 33140 19839 33192 19848
rect 33140 19805 33149 19839
rect 33149 19805 33183 19839
rect 33183 19805 33192 19839
rect 33140 19796 33192 19805
rect 33324 19839 33376 19848
rect 33324 19805 33333 19839
rect 33333 19805 33367 19839
rect 33367 19805 33376 19839
rect 33324 19796 33376 19805
rect 28632 19771 28684 19780
rect 2228 19660 2280 19712
rect 5172 19703 5224 19712
rect 5172 19669 5181 19703
rect 5181 19669 5215 19703
rect 5215 19669 5224 19703
rect 5172 19660 5224 19669
rect 6828 19660 6880 19712
rect 8944 19703 8996 19712
rect 8944 19669 8953 19703
rect 8953 19669 8987 19703
rect 8987 19669 8996 19703
rect 8944 19660 8996 19669
rect 12532 19660 12584 19712
rect 12716 19660 12768 19712
rect 14924 19703 14976 19712
rect 14924 19669 14933 19703
rect 14933 19669 14967 19703
rect 14967 19669 14976 19703
rect 14924 19660 14976 19669
rect 15936 19660 15988 19712
rect 22008 19660 22060 19712
rect 25320 19660 25372 19712
rect 28632 19737 28641 19771
rect 28641 19737 28675 19771
rect 28675 19737 28684 19771
rect 28632 19728 28684 19737
rect 32680 19728 32732 19780
rect 37464 19796 37516 19848
rect 40500 19864 40552 19916
rect 40776 19839 40828 19848
rect 40776 19805 40785 19839
rect 40785 19805 40819 19839
rect 40819 19805 40828 19839
rect 40960 19839 41012 19848
rect 40776 19796 40828 19805
rect 40960 19805 40969 19839
rect 40969 19805 41003 19839
rect 41003 19805 41012 19839
rect 40960 19796 41012 19805
rect 58164 19839 58216 19848
rect 58164 19805 58173 19839
rect 58173 19805 58207 19839
rect 58207 19805 58216 19839
rect 58164 19796 58216 19805
rect 37648 19728 37700 19780
rect 32956 19660 33008 19712
rect 36084 19660 36136 19712
rect 40408 19728 40460 19780
rect 38752 19660 38804 19712
rect 40316 19703 40368 19712
rect 40316 19669 40325 19703
rect 40325 19669 40359 19703
rect 40359 19669 40368 19703
rect 40316 19660 40368 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 4620 19456 4672 19508
rect 10784 19456 10836 19508
rect 14096 19456 14148 19508
rect 15200 19456 15252 19508
rect 18972 19456 19024 19508
rect 23480 19456 23532 19508
rect 23940 19456 23992 19508
rect 26424 19499 26476 19508
rect 26424 19465 26433 19499
rect 26433 19465 26467 19499
rect 26467 19465 26476 19499
rect 26424 19456 26476 19465
rect 26976 19499 27028 19508
rect 26976 19465 26985 19499
rect 26985 19465 27019 19499
rect 27019 19465 27028 19499
rect 26976 19456 27028 19465
rect 28632 19456 28684 19508
rect 2688 19388 2740 19440
rect 5172 19388 5224 19440
rect 6552 19388 6604 19440
rect 1952 19363 2004 19372
rect 1952 19329 1961 19363
rect 1961 19329 1995 19363
rect 1995 19329 2004 19363
rect 1952 19320 2004 19329
rect 2228 19363 2280 19372
rect 2228 19329 2262 19363
rect 2262 19329 2280 19363
rect 2228 19320 2280 19329
rect 6920 19363 6972 19372
rect 6920 19329 6954 19363
rect 6954 19329 6972 19363
rect 9588 19388 9640 19440
rect 12440 19388 12492 19440
rect 13176 19388 13228 19440
rect 6368 19252 6420 19304
rect 6920 19320 6972 19329
rect 10416 19320 10468 19372
rect 10784 19320 10836 19372
rect 12716 19320 12768 19372
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14280 19320 14332 19372
rect 20996 19388 21048 19440
rect 17408 19363 17460 19372
rect 17408 19329 17417 19363
rect 17417 19329 17451 19363
rect 17451 19329 17460 19363
rect 17408 19320 17460 19329
rect 17500 19320 17552 19372
rect 20536 19320 20588 19372
rect 22100 19388 22152 19440
rect 24768 19388 24820 19440
rect 25320 19388 25372 19440
rect 25504 19431 25556 19440
rect 25504 19397 25513 19431
rect 25513 19397 25547 19431
rect 25547 19397 25556 19431
rect 25504 19388 25556 19397
rect 27252 19388 27304 19440
rect 28264 19388 28316 19440
rect 30932 19499 30984 19508
rect 29460 19388 29512 19440
rect 7748 19184 7800 19236
rect 8116 19184 8168 19236
rect 7656 19116 7708 19168
rect 8208 19116 8260 19168
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 12532 19252 12584 19304
rect 13728 19252 13780 19304
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22744 19320 22796 19372
rect 24400 19320 24452 19372
rect 25596 19363 25648 19372
rect 22008 19295 22060 19304
rect 11152 19184 11204 19236
rect 12164 19184 12216 19236
rect 10876 19116 10928 19168
rect 15476 19159 15528 19168
rect 15476 19125 15485 19159
rect 15485 19125 15519 19159
rect 15519 19125 15528 19159
rect 15476 19116 15528 19125
rect 22008 19261 22017 19295
rect 22017 19261 22051 19295
rect 22051 19261 22060 19295
rect 22008 19252 22060 19261
rect 24952 19252 25004 19304
rect 25596 19329 25605 19363
rect 25605 19329 25639 19363
rect 25639 19329 25648 19363
rect 25596 19320 25648 19329
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 27344 19320 27396 19372
rect 27252 19295 27304 19304
rect 27252 19261 27261 19295
rect 27261 19261 27295 19295
rect 27295 19261 27304 19295
rect 27252 19252 27304 19261
rect 18972 19184 19024 19236
rect 25688 19184 25740 19236
rect 22192 19116 22244 19168
rect 22468 19116 22520 19168
rect 26424 19116 26476 19168
rect 27896 19159 27948 19168
rect 27896 19125 27905 19159
rect 27905 19125 27939 19159
rect 27939 19125 27948 19159
rect 27896 19116 27948 19125
rect 29920 19295 29972 19304
rect 29920 19261 29929 19295
rect 29929 19261 29963 19295
rect 29963 19261 29972 19295
rect 29920 19252 29972 19261
rect 30012 19184 30064 19236
rect 29828 19116 29880 19168
rect 30932 19465 30941 19499
rect 30941 19465 30975 19499
rect 30975 19465 30984 19499
rect 30932 19456 30984 19465
rect 37556 19456 37608 19508
rect 31668 19388 31720 19440
rect 36084 19431 36136 19440
rect 36084 19397 36093 19431
rect 36093 19397 36127 19431
rect 36127 19397 36136 19431
rect 36084 19388 36136 19397
rect 36268 19388 36320 19440
rect 31208 19363 31260 19372
rect 31208 19329 31217 19363
rect 31217 19329 31251 19363
rect 31251 19329 31260 19363
rect 31208 19320 31260 19329
rect 33232 19320 33284 19372
rect 34152 19320 34204 19372
rect 35808 19320 35860 19372
rect 35992 19363 36044 19372
rect 35992 19329 36001 19363
rect 36001 19329 36035 19363
rect 36035 19329 36044 19363
rect 35992 19320 36044 19329
rect 38016 19388 38068 19440
rect 40316 19388 40368 19440
rect 40776 19456 40828 19508
rect 40592 19363 40644 19372
rect 40592 19329 40601 19363
rect 40601 19329 40635 19363
rect 40635 19329 40644 19363
rect 40592 19320 40644 19329
rect 37280 19295 37332 19304
rect 37280 19261 37289 19295
rect 37289 19261 37323 19295
rect 37323 19261 37332 19295
rect 37280 19252 37332 19261
rect 38752 19295 38804 19304
rect 38752 19261 38761 19295
rect 38761 19261 38795 19295
rect 38795 19261 38804 19295
rect 38752 19252 38804 19261
rect 32680 19227 32732 19236
rect 32680 19193 32689 19227
rect 32689 19193 32723 19227
rect 32723 19193 32732 19227
rect 32680 19184 32732 19193
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2504 18955 2556 18964
rect 2504 18921 2513 18955
rect 2513 18921 2547 18955
rect 2547 18921 2556 18955
rect 2504 18912 2556 18921
rect 3976 18912 4028 18964
rect 7748 18912 7800 18964
rect 8300 18955 8352 18964
rect 8300 18921 8309 18955
rect 8309 18921 8343 18955
rect 8343 18921 8352 18955
rect 8300 18912 8352 18921
rect 8392 18912 8444 18964
rect 10416 18955 10468 18964
rect 8116 18844 8168 18896
rect 10416 18921 10425 18955
rect 10425 18921 10459 18955
rect 10459 18921 10468 18955
rect 10416 18912 10468 18921
rect 13912 18912 13964 18964
rect 14188 18912 14240 18964
rect 17500 18955 17552 18964
rect 17500 18921 17509 18955
rect 17509 18921 17543 18955
rect 17543 18921 17552 18955
rect 17500 18912 17552 18921
rect 22008 18912 22060 18964
rect 27344 18912 27396 18964
rect 4804 18776 4856 18828
rect 2780 18751 2832 18760
rect 2780 18717 2789 18751
rect 2789 18717 2823 18751
rect 2823 18717 2832 18751
rect 2780 18708 2832 18717
rect 6828 18776 6880 18828
rect 8300 18819 8352 18828
rect 8300 18785 8309 18819
rect 8309 18785 8343 18819
rect 8343 18785 8352 18819
rect 8300 18776 8352 18785
rect 7012 18751 7064 18760
rect 7012 18717 7021 18751
rect 7021 18717 7055 18751
rect 7055 18717 7064 18751
rect 7012 18708 7064 18717
rect 8208 18708 8260 18760
rect 8392 18751 8444 18760
rect 8392 18717 8401 18751
rect 8401 18717 8435 18751
rect 8435 18717 8444 18751
rect 8392 18708 8444 18717
rect 13452 18844 13504 18896
rect 17960 18844 18012 18896
rect 24584 18844 24636 18896
rect 4620 18640 4672 18692
rect 5356 18683 5408 18692
rect 5356 18649 5365 18683
rect 5365 18649 5399 18683
rect 5399 18649 5408 18683
rect 5356 18640 5408 18649
rect 5908 18640 5960 18692
rect 8576 18640 8628 18692
rect 7380 18572 7432 18624
rect 8116 18572 8168 18624
rect 10876 18751 10928 18760
rect 10876 18717 10885 18751
rect 10885 18717 10919 18751
rect 10919 18717 10928 18751
rect 10876 18708 10928 18717
rect 11152 18708 11204 18760
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 15016 18776 15068 18828
rect 12164 18751 12216 18760
rect 11520 18615 11572 18624
rect 11520 18581 11529 18615
rect 11529 18581 11563 18615
rect 11563 18581 11572 18615
rect 11520 18572 11572 18581
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 12256 18708 12308 18760
rect 12900 18708 12952 18760
rect 16580 18708 16632 18760
rect 12716 18640 12768 18692
rect 18052 18708 18104 18760
rect 18328 18708 18380 18760
rect 12808 18572 12860 18624
rect 17776 18572 17828 18624
rect 20536 18640 20588 18692
rect 22376 18776 22428 18828
rect 26884 18844 26936 18896
rect 27160 18844 27212 18896
rect 30380 18844 30432 18896
rect 30656 18887 30708 18896
rect 30656 18853 30665 18887
rect 30665 18853 30699 18887
rect 30699 18853 30708 18887
rect 30656 18844 30708 18853
rect 37372 18912 37424 18964
rect 25688 18776 25740 18828
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 25504 18708 25556 18760
rect 26608 18708 26660 18760
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 29828 18708 29880 18717
rect 30012 18751 30064 18760
rect 30012 18717 30021 18751
rect 30021 18717 30055 18751
rect 30055 18717 30064 18751
rect 30012 18708 30064 18717
rect 32036 18844 32088 18896
rect 32864 18844 32916 18896
rect 34152 18819 34204 18828
rect 34152 18785 34161 18819
rect 34161 18785 34195 18819
rect 34195 18785 34204 18819
rect 34152 18776 34204 18785
rect 31116 18751 31168 18760
rect 20904 18640 20956 18692
rect 21548 18640 21600 18692
rect 26332 18640 26384 18692
rect 27068 18640 27120 18692
rect 29920 18683 29972 18692
rect 29920 18649 29929 18683
rect 29929 18649 29963 18683
rect 29963 18649 29972 18683
rect 29920 18640 29972 18649
rect 24308 18572 24360 18624
rect 25780 18615 25832 18624
rect 25780 18581 25789 18615
rect 25789 18581 25823 18615
rect 25823 18581 25832 18615
rect 25780 18572 25832 18581
rect 26056 18572 26108 18624
rect 27528 18615 27580 18624
rect 27528 18581 27537 18615
rect 27537 18581 27571 18615
rect 27571 18581 27580 18615
rect 27528 18572 27580 18581
rect 30012 18572 30064 18624
rect 31116 18717 31125 18751
rect 31125 18717 31159 18751
rect 31159 18717 31168 18751
rect 31116 18708 31168 18717
rect 32680 18708 32732 18760
rect 35992 18708 36044 18760
rect 36268 18751 36320 18760
rect 36268 18717 36277 18751
rect 36277 18717 36311 18751
rect 36311 18717 36320 18751
rect 36268 18708 36320 18717
rect 36912 18708 36964 18760
rect 37280 18708 37332 18760
rect 40224 18776 40276 18828
rect 40132 18751 40184 18760
rect 40132 18717 40141 18751
rect 40141 18717 40175 18751
rect 40175 18717 40184 18751
rect 40132 18708 40184 18717
rect 58164 18751 58216 18760
rect 58164 18717 58173 18751
rect 58173 18717 58207 18751
rect 58207 18717 58216 18751
rect 58164 18708 58216 18717
rect 33324 18640 33376 18692
rect 33508 18640 33560 18692
rect 37648 18683 37700 18692
rect 32588 18572 32640 18624
rect 37648 18649 37657 18683
rect 37657 18649 37691 18683
rect 37691 18649 37700 18683
rect 37648 18640 37700 18649
rect 38108 18640 38160 18692
rect 39396 18572 39448 18624
rect 40776 18572 40828 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 6920 18368 6972 18420
rect 8300 18368 8352 18420
rect 18052 18411 18104 18420
rect 18052 18377 18061 18411
rect 18061 18377 18095 18411
rect 18095 18377 18104 18411
rect 18052 18368 18104 18377
rect 20904 18411 20956 18420
rect 2780 18300 2832 18352
rect 4068 18232 4120 18284
rect 5080 18300 5132 18352
rect 4620 18232 4672 18284
rect 5908 18232 5960 18284
rect 7656 18300 7708 18352
rect 11520 18300 11572 18352
rect 13728 18300 13780 18352
rect 18972 18300 19024 18352
rect 20904 18377 20913 18411
rect 20913 18377 20947 18411
rect 20947 18377 20956 18411
rect 20904 18368 20956 18377
rect 7380 18275 7432 18284
rect 7380 18241 7389 18275
rect 7389 18241 7423 18275
rect 7423 18241 7432 18275
rect 7380 18232 7432 18241
rect 8116 18232 8168 18284
rect 9588 18275 9640 18284
rect 9588 18241 9597 18275
rect 9597 18241 9631 18275
rect 9631 18241 9640 18275
rect 9588 18232 9640 18241
rect 11060 18232 11112 18284
rect 14372 18232 14424 18284
rect 4804 18164 4856 18216
rect 7196 18207 7248 18216
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7196 18164 7248 18173
rect 5540 18096 5592 18148
rect 12716 18164 12768 18216
rect 18328 18164 18380 18216
rect 22008 18343 22060 18352
rect 22008 18309 22017 18343
rect 22017 18309 22051 18343
rect 22051 18309 22060 18343
rect 22008 18300 22060 18309
rect 27528 18368 27580 18420
rect 31852 18368 31904 18420
rect 32128 18368 32180 18420
rect 33232 18368 33284 18420
rect 33508 18411 33560 18420
rect 33508 18377 33517 18411
rect 33517 18377 33551 18411
rect 33551 18377 33560 18411
rect 33508 18368 33560 18377
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 2964 18071 3016 18080
rect 2964 18037 2973 18071
rect 2973 18037 3007 18071
rect 3007 18037 3016 18071
rect 2964 18028 3016 18037
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 11796 18096 11848 18148
rect 16304 18096 16356 18148
rect 18236 18096 18288 18148
rect 24216 18300 24268 18352
rect 24768 18343 24820 18352
rect 24768 18309 24777 18343
rect 24777 18309 24811 18343
rect 24811 18309 24820 18343
rect 24768 18300 24820 18309
rect 26608 18300 26660 18352
rect 29644 18300 29696 18352
rect 37924 18368 37976 18420
rect 40132 18411 40184 18420
rect 40132 18377 40141 18411
rect 40141 18377 40175 18411
rect 40175 18377 40184 18411
rect 40132 18368 40184 18377
rect 23480 18232 23532 18284
rect 24676 18232 24728 18284
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 25964 18232 26016 18284
rect 32404 18275 32456 18284
rect 25872 18207 25924 18216
rect 25872 18173 25881 18207
rect 25881 18173 25915 18207
rect 25915 18173 25924 18207
rect 25872 18164 25924 18173
rect 32404 18241 32413 18275
rect 32413 18241 32447 18275
rect 32447 18241 32456 18275
rect 32404 18232 32456 18241
rect 32588 18275 32640 18284
rect 32588 18241 32597 18275
rect 32597 18241 32631 18275
rect 32631 18241 32640 18275
rect 32588 18232 32640 18241
rect 32772 18275 32824 18284
rect 32772 18241 32781 18275
rect 32781 18241 32815 18275
rect 32815 18241 32824 18275
rect 32772 18232 32824 18241
rect 33048 18164 33100 18216
rect 34152 18275 34204 18284
rect 34152 18241 34161 18275
rect 34161 18241 34195 18275
rect 34195 18241 34204 18275
rect 34152 18232 34204 18241
rect 38108 18232 38160 18284
rect 40132 18232 40184 18284
rect 40776 18275 40828 18284
rect 40776 18241 40785 18275
rect 40785 18241 40819 18275
rect 40819 18241 40828 18275
rect 40776 18232 40828 18241
rect 41052 18300 41104 18352
rect 34336 18164 34388 18216
rect 37188 18164 37240 18216
rect 38752 18207 38804 18216
rect 38752 18173 38761 18207
rect 38761 18173 38795 18207
rect 38795 18173 38804 18207
rect 38752 18164 38804 18173
rect 40684 18164 40736 18216
rect 5632 18028 5684 18037
rect 11152 18028 11204 18080
rect 12256 18028 12308 18080
rect 13176 18071 13228 18080
rect 13176 18037 13185 18071
rect 13185 18037 13219 18071
rect 13219 18037 13228 18071
rect 13176 18028 13228 18037
rect 13820 18028 13872 18080
rect 15568 18028 15620 18080
rect 21180 18028 21232 18080
rect 22192 18028 22244 18080
rect 27068 18028 27120 18080
rect 32128 18096 32180 18148
rect 32772 18096 32824 18148
rect 38660 18096 38712 18148
rect 33600 18028 33652 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5540 17824 5592 17876
rect 6000 17824 6052 17876
rect 13268 17824 13320 17876
rect 14372 17824 14424 17876
rect 13176 17756 13228 17808
rect 4712 17688 4764 17740
rect 5540 17620 5592 17672
rect 12808 17688 12860 17740
rect 4068 17484 4120 17536
rect 5724 17484 5776 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 6276 17484 6328 17536
rect 6828 17484 6880 17536
rect 7656 17527 7708 17536
rect 7656 17493 7665 17527
rect 7665 17493 7699 17527
rect 7699 17493 7708 17527
rect 7656 17484 7708 17493
rect 11060 17484 11112 17536
rect 11796 17527 11848 17536
rect 11796 17493 11805 17527
rect 11805 17493 11839 17527
rect 11839 17493 11848 17527
rect 11796 17484 11848 17493
rect 11888 17484 11940 17536
rect 12348 17620 12400 17672
rect 12992 17620 13044 17672
rect 13820 17688 13872 17740
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 16580 17824 16632 17876
rect 25504 17824 25556 17876
rect 26608 17867 26660 17876
rect 26608 17833 26617 17867
rect 26617 17833 26651 17867
rect 26651 17833 26660 17867
rect 26608 17824 26660 17833
rect 34336 17824 34388 17876
rect 40592 17824 40644 17876
rect 13268 17620 13320 17629
rect 15016 17552 15068 17604
rect 18788 17756 18840 17808
rect 40040 17756 40092 17808
rect 41052 17756 41104 17808
rect 20812 17688 20864 17740
rect 33416 17688 33468 17740
rect 34152 17688 34204 17740
rect 38660 17688 38712 17740
rect 40684 17688 40736 17740
rect 17316 17663 17368 17672
rect 17316 17629 17325 17663
rect 17325 17629 17359 17663
rect 17359 17629 17368 17663
rect 17316 17620 17368 17629
rect 17960 17620 18012 17672
rect 19156 17620 19208 17672
rect 20352 17620 20404 17672
rect 24124 17620 24176 17672
rect 26516 17620 26568 17672
rect 27436 17620 27488 17672
rect 28816 17620 28868 17672
rect 32864 17663 32916 17672
rect 32864 17629 32873 17663
rect 32873 17629 32907 17663
rect 32907 17629 32916 17663
rect 32864 17620 32916 17629
rect 33692 17663 33744 17672
rect 33692 17629 33701 17663
rect 33701 17629 33735 17663
rect 33735 17629 33744 17663
rect 33692 17620 33744 17629
rect 38936 17663 38988 17672
rect 38936 17629 38945 17663
rect 38945 17629 38979 17663
rect 38979 17629 38988 17663
rect 38936 17620 38988 17629
rect 17776 17552 17828 17604
rect 21180 17552 21232 17604
rect 25688 17552 25740 17604
rect 26976 17552 27028 17604
rect 16948 17484 17000 17536
rect 21824 17484 21876 17536
rect 33324 17552 33376 17604
rect 36268 17595 36320 17604
rect 36268 17561 36277 17595
rect 36277 17561 36311 17595
rect 36311 17561 36320 17595
rect 36268 17552 36320 17561
rect 37188 17552 37240 17604
rect 37832 17552 37884 17604
rect 33600 17484 33652 17536
rect 36176 17484 36228 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 5448 17280 5500 17332
rect 11888 17280 11940 17332
rect 12348 17323 12400 17332
rect 12348 17289 12357 17323
rect 12357 17289 12391 17323
rect 12391 17289 12400 17323
rect 12348 17280 12400 17289
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 13912 17323 13964 17332
rect 13912 17289 13921 17323
rect 13921 17289 13955 17323
rect 13955 17289 13964 17323
rect 13912 17280 13964 17289
rect 16028 17280 16080 17332
rect 2964 17212 3016 17264
rect 7012 17144 7064 17196
rect 8944 17212 8996 17264
rect 13084 17212 13136 17264
rect 16580 17212 16632 17264
rect 8116 17187 8168 17196
rect 8116 17153 8125 17187
rect 8125 17153 8159 17187
rect 8159 17153 8168 17187
rect 8116 17144 8168 17153
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 14004 17144 14056 17196
rect 14280 17187 14332 17196
rect 14280 17153 14289 17187
rect 14289 17153 14323 17187
rect 14323 17153 14332 17187
rect 14280 17144 14332 17153
rect 14372 17187 14424 17196
rect 14372 17153 14417 17187
rect 14417 17153 14424 17187
rect 14372 17144 14424 17153
rect 14556 17187 14608 17196
rect 14556 17153 14565 17187
rect 14565 17153 14599 17187
rect 14599 17153 14608 17187
rect 14556 17144 14608 17153
rect 1952 17076 2004 17128
rect 7196 17076 7248 17128
rect 7840 17119 7892 17128
rect 7840 17085 7849 17119
rect 7849 17085 7883 17119
rect 7883 17085 7892 17119
rect 15200 17144 15252 17196
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 16764 17144 16816 17196
rect 16948 17187 17000 17196
rect 16948 17153 16982 17187
rect 16982 17153 17000 17187
rect 16948 17144 17000 17153
rect 15016 17119 15068 17128
rect 7840 17076 7892 17085
rect 3884 17008 3936 17060
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 18512 17280 18564 17332
rect 20996 17280 21048 17332
rect 25688 17323 25740 17332
rect 25688 17289 25697 17323
rect 25697 17289 25731 17323
rect 25731 17289 25740 17323
rect 25688 17280 25740 17289
rect 26976 17323 27028 17332
rect 26976 17289 26985 17323
rect 26985 17289 27019 17323
rect 27019 17289 27028 17323
rect 26976 17280 27028 17289
rect 27344 17280 27396 17332
rect 17776 17212 17828 17264
rect 18788 17187 18840 17196
rect 18788 17153 18797 17187
rect 18797 17153 18831 17187
rect 18831 17153 18840 17187
rect 18788 17144 18840 17153
rect 21824 17212 21876 17264
rect 22100 17212 22152 17264
rect 22376 17212 22428 17264
rect 25780 17212 25832 17264
rect 18972 17187 19024 17196
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 19156 17187 19208 17196
rect 18972 17144 19024 17153
rect 19156 17153 19165 17187
rect 19165 17153 19199 17187
rect 19199 17153 19208 17187
rect 19156 17144 19208 17153
rect 24216 17144 24268 17196
rect 24952 17144 25004 17196
rect 25688 17144 25740 17196
rect 20996 17076 21048 17128
rect 22928 17076 22980 17128
rect 24032 17119 24084 17128
rect 24032 17085 24041 17119
rect 24041 17085 24075 17119
rect 24075 17085 24084 17119
rect 24032 17076 24084 17085
rect 26700 17144 26752 17196
rect 27160 17144 27212 17196
rect 27436 17187 27488 17196
rect 27436 17153 27445 17187
rect 27445 17153 27479 17187
rect 27479 17153 27488 17187
rect 32404 17280 32456 17332
rect 36268 17280 36320 17332
rect 37372 17280 37424 17332
rect 40500 17280 40552 17332
rect 29920 17212 29972 17264
rect 27436 17144 27488 17153
rect 26240 17076 26292 17128
rect 10876 17008 10928 17060
rect 4620 16940 4672 16992
rect 4712 16940 4764 16992
rect 5356 16940 5408 16992
rect 5908 16940 5960 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 9680 16940 9732 16992
rect 16028 16940 16080 16992
rect 19340 17008 19392 17060
rect 29000 17144 29052 17196
rect 33048 17144 33100 17196
rect 33416 17187 33468 17196
rect 33416 17153 33425 17187
rect 33425 17153 33459 17187
rect 33459 17153 33468 17187
rect 33416 17144 33468 17153
rect 33600 17187 33652 17196
rect 33600 17153 33609 17187
rect 33609 17153 33643 17187
rect 33643 17153 33652 17187
rect 33600 17144 33652 17153
rect 35624 17187 35676 17196
rect 35624 17153 35658 17187
rect 35658 17153 35676 17187
rect 32128 17119 32180 17128
rect 32128 17085 32137 17119
rect 32137 17085 32171 17119
rect 32171 17085 32180 17119
rect 32128 17076 32180 17085
rect 28080 17008 28132 17060
rect 18144 16940 18196 16992
rect 18328 16940 18380 16992
rect 21732 16940 21784 16992
rect 25044 16940 25096 16992
rect 29184 16940 29236 16992
rect 30472 16940 30524 16992
rect 31300 17008 31352 17060
rect 33324 17008 33376 17060
rect 35624 17144 35676 17153
rect 39948 17144 40000 17196
rect 34520 17076 34572 17128
rect 58164 17051 58216 17060
rect 34060 16983 34112 16992
rect 34060 16949 34069 16983
rect 34069 16949 34103 16983
rect 34103 16949 34112 16983
rect 34060 16940 34112 16949
rect 58164 17017 58173 17051
rect 58173 17017 58207 17051
rect 58207 17017 58216 17051
rect 58164 17008 58216 17017
rect 36360 16940 36412 16992
rect 38200 16940 38252 16992
rect 40132 16940 40184 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 9956 16736 10008 16788
rect 16304 16779 16356 16788
rect 16304 16745 16313 16779
rect 16313 16745 16347 16779
rect 16347 16745 16356 16779
rect 16304 16736 16356 16745
rect 17316 16736 17368 16788
rect 18972 16736 19024 16788
rect 21180 16779 21232 16788
rect 21180 16745 21189 16779
rect 21189 16745 21223 16779
rect 21223 16745 21232 16779
rect 21180 16736 21232 16745
rect 9496 16668 9548 16720
rect 10324 16668 10376 16720
rect 20904 16668 20956 16720
rect 24584 16736 24636 16788
rect 4620 16600 4672 16652
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 9588 16600 9640 16652
rect 2504 16532 2556 16584
rect 5540 16532 5592 16584
rect 7380 16532 7432 16584
rect 11244 16600 11296 16652
rect 16304 16532 16356 16584
rect 17776 16600 17828 16652
rect 17408 16532 17460 16584
rect 17960 16600 18012 16652
rect 18052 16532 18104 16584
rect 18236 16532 18288 16584
rect 21548 16668 21600 16720
rect 24492 16668 24544 16720
rect 25412 16668 25464 16720
rect 27436 16736 27488 16788
rect 28908 16736 28960 16788
rect 30564 16736 30616 16788
rect 33324 16779 33376 16788
rect 33324 16745 33333 16779
rect 33333 16745 33367 16779
rect 33367 16745 33376 16779
rect 33324 16736 33376 16745
rect 35624 16736 35676 16788
rect 25688 16668 25740 16720
rect 21732 16600 21784 16652
rect 26056 16600 26108 16652
rect 27252 16600 27304 16652
rect 27344 16600 27396 16652
rect 32128 16600 32180 16652
rect 14556 16464 14608 16516
rect 18144 16507 18196 16516
rect 18144 16473 18153 16507
rect 18153 16473 18187 16507
rect 18187 16473 18196 16507
rect 18144 16464 18196 16473
rect 19432 16507 19484 16516
rect 19432 16473 19441 16507
rect 19441 16473 19475 16507
rect 19475 16473 19484 16507
rect 19432 16464 19484 16473
rect 26608 16532 26660 16584
rect 29828 16532 29880 16584
rect 35624 16532 35676 16584
rect 26332 16507 26384 16516
rect 2228 16439 2280 16448
rect 2228 16405 2237 16439
rect 2237 16405 2271 16439
rect 2271 16405 2280 16439
rect 2228 16396 2280 16405
rect 5724 16396 5776 16448
rect 7012 16439 7064 16448
rect 7012 16405 7021 16439
rect 7021 16405 7055 16439
rect 7055 16405 7064 16439
rect 7012 16396 7064 16405
rect 8852 16396 8904 16448
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 11244 16396 11296 16448
rect 12164 16396 12216 16448
rect 16856 16439 16908 16448
rect 16856 16405 16865 16439
rect 16865 16405 16899 16439
rect 16899 16405 16908 16439
rect 16856 16396 16908 16405
rect 19340 16396 19392 16448
rect 26332 16473 26341 16507
rect 26341 16473 26375 16507
rect 26375 16473 26384 16507
rect 26332 16464 26384 16473
rect 26700 16464 26752 16516
rect 27160 16464 27212 16516
rect 30564 16464 30616 16516
rect 36176 16575 36228 16584
rect 36176 16541 36185 16575
rect 36185 16541 36219 16575
rect 36219 16541 36228 16575
rect 36176 16532 36228 16541
rect 36360 16575 36412 16584
rect 36360 16541 36369 16575
rect 36369 16541 36403 16575
rect 36403 16541 36412 16575
rect 36360 16532 36412 16541
rect 37832 16600 37884 16652
rect 37004 16575 37056 16584
rect 37004 16541 37013 16575
rect 37013 16541 37047 16575
rect 37047 16541 37056 16575
rect 37004 16532 37056 16541
rect 37372 16575 37424 16584
rect 37372 16541 37381 16575
rect 37381 16541 37415 16575
rect 37415 16541 37424 16575
rect 37372 16532 37424 16541
rect 38936 16532 38988 16584
rect 22468 16396 22520 16448
rect 22652 16396 22704 16448
rect 29184 16396 29236 16448
rect 30380 16396 30432 16448
rect 37648 16464 37700 16516
rect 40040 16507 40092 16516
rect 40040 16473 40049 16507
rect 40049 16473 40083 16507
rect 40083 16473 40092 16507
rect 40040 16464 40092 16473
rect 37372 16396 37424 16448
rect 40224 16439 40276 16448
rect 40224 16405 40233 16439
rect 40233 16405 40267 16439
rect 40267 16405 40276 16439
rect 40224 16396 40276 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 2228 16167 2280 16176
rect 2228 16133 2262 16167
rect 2262 16133 2280 16167
rect 2228 16124 2280 16133
rect 7840 16192 7892 16244
rect 10692 16192 10744 16244
rect 11980 16192 12032 16244
rect 17408 16235 17460 16244
rect 17408 16201 17417 16235
rect 17417 16201 17451 16235
rect 17451 16201 17460 16235
rect 17408 16192 17460 16201
rect 5724 16124 5776 16176
rect 9496 16124 9548 16176
rect 1952 16031 2004 16040
rect 1952 15997 1961 16031
rect 1961 15997 1995 16031
rect 1995 15997 2004 16031
rect 1952 15988 2004 15997
rect 3792 15895 3844 15904
rect 3792 15861 3801 15895
rect 3801 15861 3835 15895
rect 3835 15861 3844 15895
rect 3792 15852 3844 15861
rect 5540 15988 5592 16040
rect 6828 15988 6880 16040
rect 4804 15920 4856 15972
rect 5356 15920 5408 15972
rect 8116 16056 8168 16108
rect 9680 16099 9732 16108
rect 9680 16065 9689 16099
rect 9689 16065 9723 16099
rect 9723 16065 9732 16099
rect 9680 16056 9732 16065
rect 12348 16124 12400 16176
rect 12532 16167 12584 16176
rect 12532 16133 12541 16167
rect 12541 16133 12575 16167
rect 12575 16133 12584 16167
rect 12532 16124 12584 16133
rect 10508 16099 10560 16108
rect 10508 16065 10512 16099
rect 10512 16065 10546 16099
rect 10546 16065 10560 16099
rect 10508 16056 10560 16065
rect 10692 16099 10744 16108
rect 10692 16065 10701 16099
rect 10701 16065 10735 16099
rect 10735 16065 10744 16099
rect 10692 16056 10744 16065
rect 10784 16099 10836 16108
rect 10784 16065 10829 16099
rect 10829 16065 10836 16099
rect 10784 16056 10836 16065
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 12164 16056 12216 16108
rect 14188 16056 14240 16108
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 15016 16056 15068 16108
rect 4620 15852 4672 15904
rect 6920 15852 6972 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 7472 15895 7524 15904
rect 7472 15861 7481 15895
rect 7481 15861 7515 15895
rect 7515 15861 7524 15895
rect 7472 15852 7524 15861
rect 8116 15852 8168 15904
rect 8852 15852 8904 15904
rect 9220 15852 9272 15904
rect 12532 15988 12584 16040
rect 14280 15920 14332 15972
rect 18052 16056 18104 16108
rect 19248 16124 19300 16176
rect 20812 16192 20864 16244
rect 26884 16124 26936 16176
rect 28264 16167 28316 16176
rect 28264 16133 28273 16167
rect 28273 16133 28307 16167
rect 28307 16133 28316 16167
rect 28264 16124 28316 16133
rect 17960 15920 18012 15972
rect 17040 15852 17092 15904
rect 19340 16056 19392 16108
rect 20536 16056 20588 16108
rect 20996 16056 21048 16108
rect 21272 16056 21324 16108
rect 21640 16056 21692 16108
rect 22744 16099 22796 16108
rect 22744 16065 22753 16099
rect 22753 16065 22787 16099
rect 22787 16065 22796 16099
rect 22744 16056 22796 16065
rect 22928 16056 22980 16108
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 24032 16056 24084 16108
rect 26424 16056 26476 16108
rect 28172 16056 28224 16108
rect 29000 16192 29052 16244
rect 29920 16192 29972 16244
rect 33692 16192 33744 16244
rect 30564 16124 30616 16176
rect 38568 16192 38620 16244
rect 34060 16167 34112 16176
rect 34060 16133 34078 16167
rect 34078 16133 34112 16167
rect 34060 16124 34112 16133
rect 40040 16124 40092 16176
rect 23296 15988 23348 16040
rect 19892 15852 19944 15904
rect 22652 15852 22704 15904
rect 26332 15895 26384 15904
rect 26332 15861 26341 15895
rect 26341 15861 26375 15895
rect 26375 15861 26384 15895
rect 27436 15988 27488 16040
rect 29276 16099 29328 16108
rect 29276 16065 29285 16099
rect 29285 16065 29319 16099
rect 29319 16065 29328 16099
rect 29276 16056 29328 16065
rect 29920 16056 29972 16108
rect 30380 16056 30432 16108
rect 37004 16056 37056 16108
rect 37280 16056 37332 16108
rect 37648 16099 37700 16108
rect 37648 16065 37657 16099
rect 37657 16065 37691 16099
rect 37691 16065 37700 16099
rect 37648 16056 37700 16065
rect 38660 16056 38712 16108
rect 38752 16056 38804 16108
rect 39856 16056 39908 16108
rect 29460 15988 29512 16040
rect 31760 15988 31812 16040
rect 34520 15988 34572 16040
rect 35532 16031 35584 16040
rect 35532 15997 35541 16031
rect 35541 15997 35575 16031
rect 35575 15997 35584 16031
rect 35532 15988 35584 15997
rect 40684 16031 40736 16040
rect 40684 15997 40693 16031
rect 40693 15997 40727 16031
rect 40727 15997 40736 16031
rect 40684 15988 40736 15997
rect 40960 16031 41012 16040
rect 40960 15997 40969 16031
rect 40969 15997 41003 16031
rect 41003 15997 41012 16031
rect 40960 15988 41012 15997
rect 26700 15920 26752 15972
rect 28816 15920 28868 15972
rect 37280 15963 37332 15972
rect 37280 15929 37289 15963
rect 37289 15929 37323 15963
rect 37323 15929 37332 15963
rect 37280 15920 37332 15929
rect 29552 15895 29604 15904
rect 26332 15852 26384 15861
rect 29552 15861 29561 15895
rect 29561 15861 29595 15895
rect 29595 15861 29604 15895
rect 29552 15852 29604 15861
rect 58164 15895 58216 15904
rect 58164 15861 58173 15895
rect 58173 15861 58207 15895
rect 58207 15861 58216 15895
rect 58164 15852 58216 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 9772 15648 9824 15700
rect 10600 15580 10652 15632
rect 2780 15512 2832 15564
rect 10048 15555 10100 15564
rect 10048 15521 10057 15555
rect 10057 15521 10091 15555
rect 10091 15521 10100 15555
rect 10048 15512 10100 15521
rect 10692 15512 10744 15564
rect 13176 15648 13228 15700
rect 14464 15691 14516 15700
rect 14464 15657 14473 15691
rect 14473 15657 14507 15691
rect 14507 15657 14516 15691
rect 14464 15648 14516 15657
rect 14556 15648 14608 15700
rect 13084 15623 13136 15632
rect 13084 15589 13093 15623
rect 13093 15589 13127 15623
rect 13127 15589 13136 15623
rect 13084 15580 13136 15589
rect 14188 15580 14240 15632
rect 18420 15648 18472 15700
rect 19340 15691 19392 15700
rect 19340 15657 19349 15691
rect 19349 15657 19383 15691
rect 19383 15657 19392 15691
rect 19340 15648 19392 15657
rect 19892 15691 19944 15700
rect 19892 15657 19901 15691
rect 19901 15657 19935 15691
rect 19935 15657 19944 15691
rect 19892 15648 19944 15657
rect 20352 15691 20404 15700
rect 20352 15657 20361 15691
rect 20361 15657 20395 15691
rect 20395 15657 20404 15691
rect 20352 15648 20404 15657
rect 22928 15648 22980 15700
rect 23480 15648 23532 15700
rect 26240 15648 26292 15700
rect 28264 15648 28316 15700
rect 36176 15648 36228 15700
rect 37464 15648 37516 15700
rect 39856 15691 39908 15700
rect 39856 15657 39865 15691
rect 39865 15657 39899 15691
rect 39899 15657 39908 15691
rect 39856 15648 39908 15657
rect 3792 15444 3844 15496
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 10784 15487 10836 15496
rect 7288 15376 7340 15428
rect 4620 15308 4672 15360
rect 4804 15308 4856 15360
rect 6920 15351 6972 15360
rect 6920 15317 6929 15351
rect 6929 15317 6963 15351
rect 6963 15317 6972 15351
rect 6920 15308 6972 15317
rect 8484 15308 8536 15360
rect 10784 15453 10788 15487
rect 10788 15453 10822 15487
rect 10822 15453 10836 15487
rect 10784 15444 10836 15453
rect 11152 15487 11204 15496
rect 11152 15453 11160 15487
rect 11160 15453 11194 15487
rect 11194 15453 11204 15487
rect 11152 15444 11204 15453
rect 11796 15444 11848 15496
rect 13176 15444 13228 15496
rect 12624 15376 12676 15428
rect 14188 15376 14240 15428
rect 14556 15444 14608 15496
rect 22008 15580 22060 15632
rect 29000 15623 29052 15632
rect 18420 15444 18472 15496
rect 16028 15376 16080 15428
rect 19892 15376 19944 15428
rect 20352 15487 20404 15496
rect 20352 15453 20361 15487
rect 20361 15453 20395 15487
rect 20395 15453 20404 15487
rect 20536 15487 20588 15496
rect 20352 15444 20404 15453
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 22652 15512 22704 15564
rect 21456 15376 21508 15428
rect 22192 15444 22244 15496
rect 22008 15376 22060 15428
rect 22376 15376 22428 15428
rect 24308 15444 24360 15496
rect 26240 15487 26292 15496
rect 26240 15453 26249 15487
rect 26249 15453 26283 15487
rect 26283 15453 26292 15487
rect 26240 15444 26292 15453
rect 26424 15487 26476 15496
rect 26424 15453 26433 15487
rect 26433 15453 26467 15487
rect 26467 15453 26476 15487
rect 26424 15444 26476 15453
rect 14096 15308 14148 15360
rect 16304 15351 16356 15360
rect 16304 15317 16313 15351
rect 16313 15317 16347 15351
rect 16347 15317 16356 15351
rect 16304 15308 16356 15317
rect 16672 15308 16724 15360
rect 17776 15351 17828 15360
rect 17776 15317 17785 15351
rect 17785 15317 17819 15351
rect 17819 15317 17828 15351
rect 17776 15308 17828 15317
rect 19340 15308 19392 15360
rect 20352 15308 20404 15360
rect 21364 15351 21416 15360
rect 21364 15317 21373 15351
rect 21373 15317 21407 15351
rect 21407 15317 21416 15351
rect 21364 15308 21416 15317
rect 21640 15308 21692 15360
rect 26608 15376 26660 15428
rect 27252 15419 27304 15428
rect 27252 15385 27261 15419
rect 27261 15385 27295 15419
rect 27295 15385 27304 15419
rect 27252 15376 27304 15385
rect 29000 15589 29009 15623
rect 29009 15589 29043 15623
rect 29043 15589 29052 15623
rect 29000 15580 29052 15589
rect 37832 15580 37884 15632
rect 37648 15512 37700 15564
rect 28816 15487 28868 15496
rect 28816 15453 28825 15487
rect 28825 15453 28859 15487
rect 28859 15453 28868 15487
rect 28816 15444 28868 15453
rect 29552 15444 29604 15496
rect 31760 15444 31812 15496
rect 33324 15487 33376 15496
rect 33324 15453 33333 15487
rect 33333 15453 33367 15487
rect 33367 15453 33376 15487
rect 33324 15444 33376 15453
rect 33692 15444 33744 15496
rect 38200 15487 38252 15496
rect 38200 15453 38209 15487
rect 38209 15453 38243 15487
rect 38243 15453 38252 15487
rect 38200 15444 38252 15453
rect 38568 15487 38620 15496
rect 38568 15453 38577 15487
rect 38577 15453 38611 15487
rect 38611 15453 38620 15487
rect 38568 15444 38620 15453
rect 35440 15376 35492 15428
rect 37188 15376 37240 15428
rect 38660 15376 38712 15428
rect 39948 15376 40000 15428
rect 40960 15444 41012 15496
rect 27528 15308 27580 15360
rect 33324 15308 33376 15360
rect 33600 15308 33652 15360
rect 38844 15351 38896 15360
rect 38844 15317 38853 15351
rect 38853 15317 38887 15351
rect 38887 15317 38896 15351
rect 38844 15308 38896 15317
rect 40224 15308 40276 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 4988 15104 5040 15156
rect 6920 15104 6972 15156
rect 7288 15147 7340 15156
rect 5448 15036 5500 15088
rect 1952 14968 2004 15020
rect 3700 15011 3752 15020
rect 3700 14977 3734 15011
rect 3734 14977 3752 15011
rect 7288 15113 7297 15147
rect 7297 15113 7331 15147
rect 7331 15113 7340 15147
rect 7288 15104 7340 15113
rect 12716 15104 12768 15156
rect 14556 15104 14608 15156
rect 3700 14968 3752 14977
rect 5632 14764 5684 14816
rect 7196 14900 7248 14952
rect 10232 15011 10284 15020
rect 10232 14977 10241 15011
rect 10241 14977 10275 15011
rect 10275 14977 10284 15011
rect 10232 14968 10284 14977
rect 10324 14943 10376 14952
rect 10324 14909 10333 14943
rect 10333 14909 10367 14943
rect 10367 14909 10376 14943
rect 10324 14900 10376 14909
rect 6920 14764 6972 14816
rect 7932 14807 7984 14816
rect 7932 14773 7941 14807
rect 7941 14773 7975 14807
rect 7975 14773 7984 14807
rect 7932 14764 7984 14773
rect 8760 14764 8812 14816
rect 10416 14832 10468 14884
rect 12072 14968 12124 15020
rect 13084 15036 13136 15088
rect 12808 15011 12860 15020
rect 12808 14977 12817 15011
rect 12817 14977 12851 15011
rect 12851 14977 12860 15011
rect 12808 14968 12860 14977
rect 12992 14968 13044 15020
rect 12532 14832 12584 14884
rect 14004 14900 14056 14952
rect 16028 15079 16080 15088
rect 16028 15045 16037 15079
rect 16037 15045 16071 15079
rect 16071 15045 16080 15079
rect 16028 15036 16080 15045
rect 16764 15036 16816 15088
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 19248 15036 19300 15088
rect 18328 15011 18380 15020
rect 18328 14977 18362 15011
rect 18362 14977 18380 15011
rect 16304 14900 16356 14952
rect 18328 14968 18380 14977
rect 20168 14968 20220 15020
rect 20996 15104 21048 15156
rect 21548 15104 21600 15156
rect 21180 14968 21232 15020
rect 26240 15104 26292 15156
rect 12716 14832 12768 14884
rect 17132 14832 17184 14884
rect 19432 14875 19484 14884
rect 19432 14841 19441 14875
rect 19441 14841 19475 14875
rect 19475 14841 19484 14875
rect 22192 14968 22244 15020
rect 22652 14968 22704 15020
rect 22836 15036 22888 15088
rect 23112 15079 23164 15088
rect 23112 15045 23121 15079
rect 23121 15045 23155 15079
rect 23155 15045 23164 15079
rect 23112 15036 23164 15045
rect 26608 15036 26660 15088
rect 27252 15036 27304 15088
rect 28172 15036 28224 15088
rect 28632 15036 28684 15088
rect 30380 15104 30432 15156
rect 38660 15104 38712 15156
rect 37832 15079 37884 15088
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 24400 14968 24452 15020
rect 23204 14900 23256 14952
rect 25044 14943 25096 14952
rect 25044 14909 25053 14943
rect 25053 14909 25087 14943
rect 25087 14909 25096 14943
rect 25044 14900 25096 14909
rect 25504 14900 25556 14952
rect 29552 14968 29604 15020
rect 28356 14900 28408 14952
rect 29920 14900 29972 14952
rect 30472 15011 30524 15020
rect 30472 14977 30481 15011
rect 30481 14977 30515 15011
rect 30515 14977 30524 15011
rect 30472 14968 30524 14977
rect 19432 14832 19484 14841
rect 27988 14832 28040 14884
rect 29460 14832 29512 14884
rect 10232 14764 10284 14816
rect 12624 14764 12676 14816
rect 14372 14764 14424 14816
rect 18420 14764 18472 14816
rect 21364 14764 21416 14816
rect 22192 14764 22244 14816
rect 22560 14764 22612 14816
rect 23296 14764 23348 14816
rect 23480 14807 23532 14816
rect 23480 14773 23489 14807
rect 23489 14773 23523 14807
rect 23523 14773 23532 14807
rect 23480 14764 23532 14773
rect 24032 14807 24084 14816
rect 24032 14773 24041 14807
rect 24041 14773 24075 14807
rect 24075 14773 24084 14807
rect 24032 14764 24084 14773
rect 24216 14807 24268 14816
rect 24216 14773 24225 14807
rect 24225 14773 24259 14807
rect 24259 14773 24268 14807
rect 24216 14764 24268 14773
rect 24308 14764 24360 14816
rect 27804 14764 27856 14816
rect 29552 14807 29604 14816
rect 29552 14773 29561 14807
rect 29561 14773 29595 14807
rect 29595 14773 29604 14807
rect 29552 14764 29604 14773
rect 33416 14968 33468 15020
rect 35440 15011 35492 15020
rect 35440 14977 35449 15011
rect 35449 14977 35483 15011
rect 35483 14977 35492 15011
rect 35440 14968 35492 14977
rect 37832 15045 37841 15079
rect 37841 15045 37875 15079
rect 37875 15045 37884 15079
rect 37832 15036 37884 15045
rect 38844 15036 38896 15088
rect 33692 14900 33744 14952
rect 36728 14968 36780 15020
rect 38660 14900 38712 14952
rect 35440 14832 35492 14884
rect 37648 14875 37700 14884
rect 37648 14841 37657 14875
rect 37657 14841 37691 14875
rect 37691 14841 37700 14875
rect 37648 14832 37700 14841
rect 35992 14764 36044 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2780 14560 2832 14612
rect 3700 14560 3752 14612
rect 12808 14560 12860 14612
rect 14464 14560 14516 14612
rect 17960 14603 18012 14612
rect 17960 14569 17969 14603
rect 17969 14569 18003 14603
rect 18003 14569 18012 14603
rect 17960 14560 18012 14569
rect 1584 14492 1636 14544
rect 7656 14492 7708 14544
rect 10416 14492 10468 14544
rect 14372 14492 14424 14544
rect 18144 14492 18196 14544
rect 18420 14424 18472 14476
rect 20168 14467 20220 14476
rect 3976 14399 4028 14408
rect 3976 14365 3985 14399
rect 3985 14365 4019 14399
rect 4019 14365 4028 14399
rect 3976 14356 4028 14365
rect 4804 14288 4856 14340
rect 8944 14288 8996 14340
rect 11796 14356 11848 14408
rect 16672 14356 16724 14408
rect 16856 14399 16908 14408
rect 16856 14365 16890 14399
rect 16890 14365 16908 14399
rect 16856 14356 16908 14365
rect 19340 14356 19392 14408
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 21456 14467 21508 14476
rect 21456 14433 21465 14467
rect 21465 14433 21499 14467
rect 21499 14433 21508 14467
rect 21456 14424 21508 14433
rect 19984 14356 20036 14408
rect 20076 14356 20128 14408
rect 20260 14356 20312 14408
rect 22744 14424 22796 14476
rect 22560 14356 22612 14408
rect 24216 14560 24268 14612
rect 24492 14603 24544 14612
rect 24492 14569 24501 14603
rect 24501 14569 24535 14603
rect 24535 14569 24544 14603
rect 24492 14560 24544 14569
rect 26608 14560 26660 14612
rect 27712 14560 27764 14612
rect 30380 14560 30432 14612
rect 23664 14492 23716 14544
rect 28356 14535 28408 14544
rect 28356 14501 28365 14535
rect 28365 14501 28399 14535
rect 28399 14501 28408 14535
rect 28356 14492 28408 14501
rect 29184 14492 29236 14544
rect 23112 14356 23164 14408
rect 25504 14424 25556 14476
rect 26516 14467 26568 14476
rect 26516 14433 26525 14467
rect 26525 14433 26559 14467
rect 26559 14433 26568 14467
rect 26516 14424 26568 14433
rect 27988 14424 28040 14476
rect 35532 14424 35584 14476
rect 37740 14560 37792 14612
rect 38936 14560 38988 14612
rect 40132 14560 40184 14612
rect 38936 14424 38988 14476
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 24860 14356 24912 14408
rect 29828 14356 29880 14408
rect 15200 14331 15252 14340
rect 6920 14220 6972 14272
rect 7288 14220 7340 14272
rect 10232 14220 10284 14272
rect 12900 14220 12952 14272
rect 15200 14297 15218 14331
rect 15218 14297 15252 14331
rect 15200 14288 15252 14297
rect 21364 14288 21416 14340
rect 20168 14220 20220 14272
rect 23112 14220 23164 14272
rect 27068 14288 27120 14340
rect 27252 14331 27304 14340
rect 27252 14297 27286 14331
rect 27286 14297 27304 14331
rect 27252 14288 27304 14297
rect 27436 14288 27488 14340
rect 35164 14356 35216 14408
rect 35348 14399 35400 14408
rect 35348 14365 35357 14399
rect 35357 14365 35391 14399
rect 35391 14365 35400 14399
rect 35348 14356 35400 14365
rect 36176 14399 36228 14408
rect 36176 14365 36185 14399
rect 36185 14365 36219 14399
rect 36219 14365 36228 14399
rect 36176 14356 36228 14365
rect 40684 14356 40736 14408
rect 58164 14399 58216 14408
rect 58164 14365 58173 14399
rect 58173 14365 58207 14399
rect 58207 14365 58216 14399
rect 58164 14356 58216 14365
rect 30380 14288 30432 14340
rect 28816 14220 28868 14272
rect 31760 14220 31812 14272
rect 34520 14220 34572 14272
rect 38660 14220 38712 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 3976 14016 4028 14068
rect 6552 14016 6604 14068
rect 11060 14016 11112 14068
rect 12532 14016 12584 14068
rect 4804 13948 4856 14000
rect 8944 13948 8996 14000
rect 14464 13991 14516 14000
rect 14464 13957 14473 13991
rect 14473 13957 14507 13991
rect 14507 13957 14516 13991
rect 14464 13948 14516 13957
rect 15844 13948 15896 14000
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 5172 13880 5224 13932
rect 5632 13880 5684 13932
rect 13912 13880 13964 13932
rect 17776 13948 17828 14000
rect 19340 13991 19392 14000
rect 19340 13957 19349 13991
rect 19349 13957 19383 13991
rect 19383 13957 19392 13991
rect 19340 13948 19392 13957
rect 20076 13923 20128 13932
rect 20076 13889 20085 13923
rect 20085 13889 20119 13923
rect 20119 13889 20128 13923
rect 20076 13880 20128 13889
rect 5724 13812 5776 13864
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 8024 13812 8076 13864
rect 8576 13812 8628 13864
rect 16304 13812 16356 13864
rect 17500 13812 17552 13864
rect 12072 13744 12124 13796
rect 15568 13744 15620 13796
rect 20168 13812 20220 13864
rect 22100 13880 22152 13932
rect 22376 13948 22428 14000
rect 23664 14016 23716 14068
rect 23940 14059 23992 14068
rect 23940 14025 23949 14059
rect 23949 14025 23983 14059
rect 23983 14025 23992 14059
rect 23940 14016 23992 14025
rect 25136 14016 25188 14068
rect 27252 14059 27304 14068
rect 27252 14025 27261 14059
rect 27261 14025 27295 14059
rect 27295 14025 27304 14059
rect 27252 14016 27304 14025
rect 29828 14016 29880 14068
rect 23296 13855 23348 13864
rect 23296 13821 23305 13855
rect 23305 13821 23339 13855
rect 23339 13821 23348 13855
rect 23296 13812 23348 13821
rect 24032 13880 24084 13932
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 23664 13812 23716 13864
rect 26332 13948 26384 14000
rect 28632 13991 28684 14000
rect 28632 13957 28641 13991
rect 28641 13957 28675 13991
rect 28675 13957 28684 13991
rect 28632 13948 28684 13957
rect 28816 13991 28868 14000
rect 28816 13957 28825 13991
rect 28825 13957 28859 13991
rect 28859 13957 28868 13991
rect 28816 13948 28868 13957
rect 26424 13923 26476 13932
rect 26424 13889 26433 13923
rect 26433 13889 26467 13923
rect 26467 13889 26476 13923
rect 26424 13880 26476 13889
rect 27804 13880 27856 13932
rect 28080 13880 28132 13932
rect 29460 13923 29512 13932
rect 29460 13889 29469 13923
rect 29469 13889 29503 13923
rect 29503 13889 29512 13923
rect 29460 13880 29512 13889
rect 30656 13991 30708 14000
rect 30656 13957 30665 13991
rect 30665 13957 30699 13991
rect 30699 13957 30708 13991
rect 31484 14016 31536 14068
rect 35992 14016 36044 14068
rect 39764 14059 39816 14068
rect 30656 13948 30708 13957
rect 37188 13948 37240 14000
rect 37648 13948 37700 14000
rect 39764 14025 39773 14059
rect 39773 14025 39807 14059
rect 39807 14025 39816 14059
rect 39764 14016 39816 14025
rect 31300 13880 31352 13932
rect 33140 13880 33192 13932
rect 34612 13880 34664 13932
rect 35164 13923 35216 13932
rect 35164 13889 35173 13923
rect 35173 13889 35207 13923
rect 35207 13889 35216 13923
rect 35164 13880 35216 13889
rect 35440 13880 35492 13932
rect 38752 13923 38804 13932
rect 29920 13812 29972 13864
rect 30564 13812 30616 13864
rect 35900 13812 35952 13864
rect 27436 13744 27488 13796
rect 35348 13744 35400 13796
rect 37280 13855 37332 13864
rect 37280 13821 37289 13855
rect 37289 13821 37323 13855
rect 37323 13821 37332 13855
rect 37280 13812 37332 13821
rect 37556 13855 37608 13864
rect 37556 13821 37565 13855
rect 37565 13821 37599 13855
rect 37599 13821 37608 13855
rect 37556 13812 37608 13821
rect 38752 13889 38761 13923
rect 38761 13889 38795 13923
rect 38795 13889 38804 13923
rect 38752 13880 38804 13889
rect 40684 13948 40736 14000
rect 38936 13923 38988 13932
rect 38936 13889 38945 13923
rect 38945 13889 38979 13923
rect 38979 13889 38988 13923
rect 38936 13880 38988 13889
rect 39764 13812 39816 13864
rect 4896 13676 4948 13728
rect 7012 13676 7064 13728
rect 15016 13676 15068 13728
rect 19156 13676 19208 13728
rect 21824 13676 21876 13728
rect 23112 13676 23164 13728
rect 23480 13676 23532 13728
rect 33324 13719 33376 13728
rect 33324 13685 33333 13719
rect 33333 13685 33367 13719
rect 33367 13685 33376 13719
rect 33324 13676 33376 13685
rect 37740 13676 37792 13728
rect 39212 13719 39264 13728
rect 39212 13685 39221 13719
rect 39221 13685 39255 13719
rect 39255 13685 39264 13719
rect 39212 13676 39264 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 12256 13472 12308 13524
rect 15200 13472 15252 13524
rect 21180 13472 21232 13524
rect 22192 13515 22244 13524
rect 22192 13481 22201 13515
rect 22201 13481 22235 13515
rect 22235 13481 22244 13515
rect 22192 13472 22244 13481
rect 27068 13515 27120 13524
rect 27068 13481 27077 13515
rect 27077 13481 27111 13515
rect 27111 13481 27120 13515
rect 27068 13472 27120 13481
rect 27712 13472 27764 13524
rect 28816 13472 28868 13524
rect 31300 13472 31352 13524
rect 33140 13515 33192 13524
rect 14832 13404 14884 13456
rect 17960 13404 18012 13456
rect 2780 13336 2832 13388
rect 5632 13379 5684 13388
rect 5632 13345 5641 13379
rect 5641 13345 5675 13379
rect 5675 13345 5684 13379
rect 5632 13336 5684 13345
rect 6184 13336 6236 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 8944 13379 8996 13388
rect 8944 13345 8953 13379
rect 8953 13345 8987 13379
rect 8987 13345 8996 13379
rect 8944 13336 8996 13345
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 6552 13268 6604 13320
rect 8208 13268 8260 13320
rect 8392 13268 8444 13320
rect 10048 13268 10100 13320
rect 11428 13268 11480 13320
rect 2044 13132 2096 13184
rect 4620 13175 4672 13184
rect 4620 13141 4629 13175
rect 4629 13141 4663 13175
rect 4663 13141 4672 13175
rect 4620 13132 4672 13141
rect 5540 13175 5592 13184
rect 5540 13141 5549 13175
rect 5549 13141 5583 13175
rect 5583 13141 5592 13175
rect 5540 13132 5592 13141
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 15016 13336 15068 13388
rect 15384 13268 15436 13320
rect 15660 13268 15712 13320
rect 15568 13243 15620 13252
rect 15568 13209 15577 13243
rect 15577 13209 15611 13243
rect 15611 13209 15620 13243
rect 15568 13200 15620 13209
rect 17500 13243 17552 13252
rect 17500 13209 17509 13243
rect 17509 13209 17543 13243
rect 17543 13209 17552 13243
rect 17500 13200 17552 13209
rect 20904 13404 20956 13456
rect 23848 13379 23900 13388
rect 23848 13345 23857 13379
rect 23857 13345 23891 13379
rect 23891 13345 23900 13379
rect 23848 13336 23900 13345
rect 19432 13268 19484 13320
rect 26240 13336 26292 13388
rect 26516 13379 26568 13388
rect 26516 13345 26525 13379
rect 26525 13345 26559 13379
rect 26559 13345 26568 13379
rect 26516 13336 26568 13345
rect 31760 13336 31812 13388
rect 33140 13481 33149 13515
rect 33149 13481 33183 13515
rect 33183 13481 33192 13515
rect 33140 13472 33192 13481
rect 35900 13472 35952 13524
rect 38752 13472 38804 13524
rect 20720 13200 20772 13252
rect 27252 13268 27304 13320
rect 27436 13311 27488 13320
rect 27436 13277 27445 13311
rect 27445 13277 27479 13311
rect 27479 13277 27488 13311
rect 27436 13268 27488 13277
rect 27528 13311 27580 13320
rect 27528 13277 27537 13311
rect 27537 13277 27571 13311
rect 27571 13277 27580 13311
rect 27528 13268 27580 13277
rect 28080 13268 28132 13320
rect 32496 13311 32548 13320
rect 32496 13277 32505 13311
rect 32505 13277 32539 13311
rect 32539 13277 32548 13311
rect 32496 13268 32548 13277
rect 32680 13311 32732 13320
rect 32680 13277 32689 13311
rect 32689 13277 32723 13311
rect 32723 13277 32732 13311
rect 32680 13268 32732 13277
rect 35348 13336 35400 13388
rect 35716 13311 35768 13320
rect 25228 13200 25280 13252
rect 30564 13200 30616 13252
rect 31024 13200 31076 13252
rect 35716 13277 35725 13311
rect 35725 13277 35759 13311
rect 35759 13277 35768 13311
rect 35716 13268 35768 13277
rect 35992 13311 36044 13320
rect 35992 13277 36001 13311
rect 36001 13277 36035 13311
rect 36035 13277 36044 13311
rect 35992 13268 36044 13277
rect 36728 13311 36780 13320
rect 36728 13277 36737 13311
rect 36737 13277 36771 13311
rect 36771 13277 36780 13311
rect 36728 13268 36780 13277
rect 38016 13311 38068 13320
rect 38016 13277 38025 13311
rect 38025 13277 38059 13311
rect 38059 13277 38068 13311
rect 38016 13268 38068 13277
rect 58164 13311 58216 13320
rect 58164 13277 58173 13311
rect 58173 13277 58207 13311
rect 58207 13277 58216 13311
rect 58164 13268 58216 13277
rect 15292 13132 15344 13184
rect 19156 13132 19208 13184
rect 24400 13132 24452 13184
rect 34704 13200 34756 13252
rect 37280 13200 37332 13252
rect 37556 13200 37608 13252
rect 33600 13175 33652 13184
rect 33600 13141 33609 13175
rect 33609 13141 33643 13175
rect 33643 13141 33652 13175
rect 33600 13132 33652 13141
rect 36360 13132 36412 13184
rect 39488 13132 39540 13184
rect 39948 13132 40000 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 2320 12928 2372 12980
rect 5540 12928 5592 12980
rect 9404 12928 9456 12980
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 3792 12860 3844 12912
rect 4620 12792 4672 12844
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 6736 12792 6788 12844
rect 7564 12792 7616 12844
rect 8300 12792 8352 12844
rect 9680 12860 9732 12912
rect 9772 12860 9824 12912
rect 10876 12928 10928 12980
rect 21824 12971 21876 12980
rect 13912 12903 13964 12912
rect 13912 12869 13921 12903
rect 13921 12869 13955 12903
rect 13955 12869 13964 12903
rect 13912 12860 13964 12869
rect 14096 12903 14148 12912
rect 14096 12869 14105 12903
rect 14105 12869 14139 12903
rect 14139 12869 14148 12903
rect 14096 12860 14148 12869
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 11704 12835 11756 12844
rect 10048 12792 10100 12801
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 21824 12937 21833 12971
rect 21833 12937 21867 12971
rect 21867 12937 21876 12971
rect 21824 12928 21876 12937
rect 23848 12928 23900 12980
rect 24032 12928 24084 12980
rect 24216 12928 24268 12980
rect 32680 12971 32732 12980
rect 32680 12937 32689 12971
rect 32689 12937 32723 12971
rect 32723 12937 32732 12971
rect 32680 12928 32732 12937
rect 35900 12928 35952 12980
rect 16764 12860 16816 12912
rect 11888 12767 11940 12776
rect 9588 12656 9640 12708
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 9864 12656 9916 12708
rect 11888 12733 11897 12767
rect 11897 12733 11931 12767
rect 11931 12733 11940 12767
rect 11888 12724 11940 12733
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 10048 12656 10100 12708
rect 15384 12835 15436 12844
rect 15384 12801 15393 12835
rect 15393 12801 15427 12835
rect 15427 12801 15436 12835
rect 23112 12860 23164 12912
rect 23756 12860 23808 12912
rect 33140 12860 33192 12912
rect 33324 12860 33376 12912
rect 36728 12928 36780 12980
rect 38016 12928 38068 12980
rect 37372 12860 37424 12912
rect 37740 12860 37792 12912
rect 39212 12860 39264 12912
rect 15384 12792 15436 12801
rect 15292 12724 15344 12776
rect 16120 12724 16172 12776
rect 16764 12724 16816 12776
rect 15752 12656 15804 12708
rect 11612 12588 11664 12640
rect 15200 12588 15252 12640
rect 15660 12588 15712 12640
rect 19156 12792 19208 12844
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 20996 12835 21048 12844
rect 19248 12792 19300 12801
rect 20996 12801 21005 12835
rect 21005 12801 21039 12835
rect 21039 12801 21048 12835
rect 20996 12792 21048 12801
rect 22928 12835 22980 12844
rect 22928 12801 22937 12835
rect 22937 12801 22971 12835
rect 22971 12801 22980 12835
rect 22928 12792 22980 12801
rect 31668 12792 31720 12844
rect 33600 12792 33652 12844
rect 35716 12792 35768 12844
rect 33416 12767 33468 12776
rect 18972 12656 19024 12708
rect 33416 12733 33425 12767
rect 33425 12733 33459 12767
rect 33459 12733 33468 12767
rect 33416 12724 33468 12733
rect 25596 12656 25648 12708
rect 29184 12656 29236 12708
rect 36360 12835 36412 12844
rect 36360 12801 36369 12835
rect 36369 12801 36403 12835
rect 36403 12801 36412 12835
rect 36360 12792 36412 12801
rect 36544 12792 36596 12844
rect 38660 12835 38712 12844
rect 38660 12801 38669 12835
rect 38669 12801 38703 12835
rect 38703 12801 38712 12835
rect 38660 12792 38712 12801
rect 19156 12588 19208 12640
rect 27252 12588 27304 12640
rect 36728 12631 36780 12640
rect 36728 12597 36737 12631
rect 36737 12597 36771 12631
rect 36771 12597 36780 12631
rect 36728 12588 36780 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 7564 12427 7616 12436
rect 7564 12393 7573 12427
rect 7573 12393 7607 12427
rect 7607 12393 7616 12427
rect 7564 12384 7616 12393
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 5540 12248 5592 12300
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 8024 12291 8076 12300
rect 6184 12248 6236 12257
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 2596 12223 2648 12232
rect 2596 12189 2605 12223
rect 2605 12189 2639 12223
rect 2639 12189 2648 12223
rect 2596 12180 2648 12189
rect 3056 12112 3108 12164
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 5540 12044 5592 12096
rect 7012 12180 7064 12232
rect 14096 12427 14148 12436
rect 8300 12316 8352 12368
rect 9128 12316 9180 12368
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 18236 12384 18288 12436
rect 21180 12384 21232 12436
rect 22192 12384 22244 12436
rect 22376 12384 22428 12436
rect 27160 12384 27212 12436
rect 35624 12384 35676 12436
rect 36544 12384 36596 12436
rect 37464 12384 37516 12436
rect 16120 12248 16172 12300
rect 18144 12316 18196 12368
rect 19248 12316 19300 12368
rect 29368 12316 29420 12368
rect 30840 12316 30892 12368
rect 31484 12316 31536 12368
rect 8392 12180 8444 12232
rect 9772 12223 9824 12232
rect 9772 12189 9806 12223
rect 9806 12189 9824 12223
rect 9772 12180 9824 12189
rect 11428 12180 11480 12232
rect 11612 12223 11664 12232
rect 11612 12189 11646 12223
rect 11646 12189 11664 12223
rect 11612 12180 11664 12189
rect 13912 12180 13964 12232
rect 15200 12223 15252 12232
rect 15200 12189 15218 12223
rect 15218 12189 15252 12223
rect 15200 12180 15252 12189
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 16028 12180 16080 12232
rect 9588 12112 9640 12164
rect 12348 12112 12400 12164
rect 13728 12112 13780 12164
rect 16764 12180 16816 12232
rect 17500 12180 17552 12232
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 18972 12248 19024 12300
rect 7104 12044 7156 12096
rect 9680 12044 9732 12096
rect 11704 12044 11756 12096
rect 12716 12087 12768 12096
rect 12716 12053 12725 12087
rect 12725 12053 12759 12087
rect 12759 12053 12768 12087
rect 12716 12044 12768 12053
rect 16672 12112 16724 12164
rect 14832 12044 14884 12096
rect 18144 12044 18196 12096
rect 18328 12044 18380 12096
rect 18696 12180 18748 12232
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 20628 12180 20680 12232
rect 20720 12180 20772 12232
rect 20996 12223 21048 12232
rect 20996 12189 21005 12223
rect 21005 12189 21039 12223
rect 21039 12189 21048 12223
rect 20996 12180 21048 12189
rect 24584 12248 24636 12300
rect 25320 12223 25372 12232
rect 19984 12155 20036 12164
rect 19984 12121 19993 12155
rect 19993 12121 20027 12155
rect 20027 12121 20036 12155
rect 19984 12112 20036 12121
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 25320 12189 25329 12223
rect 25329 12189 25363 12223
rect 25363 12189 25372 12223
rect 25320 12180 25372 12189
rect 25780 12248 25832 12300
rect 25504 12180 25556 12232
rect 31760 12248 31812 12300
rect 32496 12248 32548 12300
rect 31300 12223 31352 12232
rect 31300 12189 31309 12223
rect 31309 12189 31343 12223
rect 31343 12189 31352 12223
rect 31300 12180 31352 12189
rect 21732 12112 21784 12164
rect 28264 12155 28316 12164
rect 28264 12121 28273 12155
rect 28273 12121 28307 12155
rect 28307 12121 28316 12155
rect 28264 12112 28316 12121
rect 31024 12112 31076 12164
rect 31484 12223 31536 12232
rect 31484 12189 31493 12223
rect 31493 12189 31527 12223
rect 31527 12189 31536 12223
rect 31484 12180 31536 12189
rect 34520 12180 34572 12232
rect 38384 12180 38436 12232
rect 36728 12112 36780 12164
rect 22468 12044 22520 12096
rect 23480 12044 23532 12096
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 32404 12044 32456 12096
rect 34612 12044 34664 12096
rect 35808 12044 35860 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 3056 11883 3108 11892
rect 3056 11849 3065 11883
rect 3065 11849 3099 11883
rect 3099 11849 3108 11883
rect 3056 11840 3108 11849
rect 9864 11840 9916 11892
rect 13728 11883 13780 11892
rect 13728 11849 13737 11883
rect 13737 11849 13771 11883
rect 13771 11849 13780 11883
rect 13728 11840 13780 11849
rect 14740 11840 14792 11892
rect 15016 11840 15068 11892
rect 15568 11840 15620 11892
rect 16672 11840 16724 11892
rect 6828 11772 6880 11824
rect 14832 11815 14884 11824
rect 14832 11781 14850 11815
rect 14850 11781 14884 11815
rect 19984 11840 20036 11892
rect 14832 11772 14884 11781
rect 2872 11747 2924 11756
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 2872 11704 2924 11713
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 6644 11704 6696 11756
rect 8024 11704 8076 11756
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 2596 11636 2648 11688
rect 5540 11568 5592 11620
rect 5724 11568 5776 11620
rect 6736 11636 6788 11688
rect 11336 11636 11388 11688
rect 6920 11500 6972 11552
rect 7564 11500 7616 11552
rect 7840 11500 7892 11552
rect 8208 11500 8260 11552
rect 12256 11500 12308 11552
rect 15476 11704 15528 11756
rect 20444 11772 20496 11824
rect 20628 11772 20680 11824
rect 25320 11840 25372 11892
rect 29644 11883 29696 11892
rect 29644 11849 29653 11883
rect 29653 11849 29687 11883
rect 29687 11849 29696 11883
rect 29644 11840 29696 11849
rect 31300 11840 31352 11892
rect 34704 11840 34756 11892
rect 18144 11747 18196 11756
rect 18144 11713 18162 11747
rect 18162 11713 18196 11747
rect 18144 11704 18196 11713
rect 18328 11704 18380 11756
rect 19340 11704 19392 11756
rect 20536 11704 20588 11756
rect 20720 11704 20772 11756
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 24952 11772 25004 11824
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 22744 11747 22796 11756
rect 22744 11713 22753 11747
rect 22753 11713 22787 11747
rect 22787 11713 22796 11747
rect 22744 11704 22796 11713
rect 23112 11704 23164 11756
rect 23388 11747 23440 11756
rect 23388 11713 23397 11747
rect 23397 11713 23431 11747
rect 23431 11713 23440 11747
rect 23388 11704 23440 11713
rect 23480 11704 23532 11756
rect 21548 11636 21600 11688
rect 24860 11679 24912 11688
rect 24860 11645 24869 11679
rect 24869 11645 24903 11679
rect 24903 11645 24912 11679
rect 24860 11636 24912 11645
rect 19156 11611 19208 11620
rect 19156 11577 19165 11611
rect 19165 11577 19199 11611
rect 19199 11577 19208 11611
rect 19156 11568 19208 11577
rect 16028 11500 16080 11552
rect 16764 11500 16816 11552
rect 22744 11568 22796 11620
rect 28264 11704 28316 11756
rect 30840 11772 30892 11824
rect 31668 11772 31720 11824
rect 36268 11772 36320 11824
rect 39488 11815 39540 11824
rect 39488 11781 39497 11815
rect 39497 11781 39531 11815
rect 39531 11781 39540 11815
rect 39488 11772 39540 11781
rect 30564 11747 30616 11756
rect 30564 11713 30573 11747
rect 30573 11713 30607 11747
rect 30607 11713 30616 11747
rect 30564 11704 30616 11713
rect 31760 11704 31812 11756
rect 32404 11704 32456 11756
rect 33232 11704 33284 11756
rect 33416 11704 33468 11756
rect 35348 11747 35400 11756
rect 35348 11713 35357 11747
rect 35357 11713 35391 11747
rect 35391 11713 35400 11747
rect 35348 11704 35400 11713
rect 35532 11747 35584 11756
rect 35532 11713 35541 11747
rect 35541 11713 35575 11747
rect 35575 11713 35584 11747
rect 35532 11704 35584 11713
rect 35624 11704 35676 11756
rect 37740 11704 37792 11756
rect 38292 11679 38344 11688
rect 38292 11645 38301 11679
rect 38301 11645 38335 11679
rect 38335 11645 38344 11679
rect 38292 11636 38344 11645
rect 33968 11568 34020 11620
rect 35716 11568 35768 11620
rect 39120 11568 39172 11620
rect 58164 11611 58216 11620
rect 58164 11577 58173 11611
rect 58173 11577 58207 11611
rect 58207 11577 58216 11611
rect 58164 11568 58216 11577
rect 21824 11500 21876 11552
rect 22192 11500 22244 11552
rect 23112 11500 23164 11552
rect 25044 11500 25096 11552
rect 30288 11500 30340 11552
rect 38108 11500 38160 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 8024 11339 8076 11348
rect 8024 11305 8033 11339
rect 8033 11305 8067 11339
rect 8067 11305 8076 11339
rect 8024 11296 8076 11305
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 20536 11339 20588 11348
rect 20536 11305 20545 11339
rect 20545 11305 20579 11339
rect 20579 11305 20588 11339
rect 20536 11296 20588 11305
rect 7196 11228 7248 11280
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 11612 11228 11664 11280
rect 21548 11203 21600 11212
rect 21548 11169 21557 11203
rect 21557 11169 21591 11203
rect 21591 11169 21600 11203
rect 21548 11160 21600 11169
rect 24860 11160 24912 11212
rect 26240 11296 26292 11348
rect 36268 11339 36320 11348
rect 36268 11305 36277 11339
rect 36277 11305 36311 11339
rect 36311 11305 36320 11339
rect 36268 11296 36320 11305
rect 38108 11339 38160 11348
rect 38108 11305 38117 11339
rect 38117 11305 38151 11339
rect 38151 11305 38160 11339
rect 38108 11296 38160 11305
rect 39304 11296 39356 11348
rect 29920 11228 29972 11280
rect 30196 11228 30248 11280
rect 32496 11160 32548 11212
rect 33232 11160 33284 11212
rect 34520 11160 34572 11212
rect 39120 11228 39172 11280
rect 7288 11135 7340 11144
rect 7288 11101 7297 11135
rect 7297 11101 7331 11135
rect 7331 11101 7340 11135
rect 7288 11092 7340 11101
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 21824 11135 21876 11144
rect 21824 11101 21858 11135
rect 21858 11101 21876 11135
rect 21824 11092 21876 11101
rect 23112 11092 23164 11144
rect 23388 11092 23440 11144
rect 23756 11135 23808 11144
rect 23756 11101 23765 11135
rect 23765 11101 23799 11135
rect 23799 11101 23808 11135
rect 23756 11092 23808 11101
rect 24952 11092 25004 11144
rect 25320 11135 25372 11144
rect 25320 11101 25329 11135
rect 25329 11101 25363 11135
rect 25363 11101 25372 11135
rect 25320 11092 25372 11101
rect 30196 11135 30248 11144
rect 30196 11101 30205 11135
rect 30205 11101 30239 11135
rect 30239 11101 30248 11135
rect 30196 11092 30248 11101
rect 30288 11092 30340 11144
rect 38936 11135 38988 11144
rect 38936 11101 38945 11135
rect 38945 11101 38979 11135
rect 38979 11101 38988 11135
rect 38936 11092 38988 11101
rect 39304 11135 39356 11144
rect 39304 11101 39313 11135
rect 39313 11101 39347 11135
rect 39347 11101 39356 11135
rect 39304 11092 39356 11101
rect 40408 11092 40460 11144
rect 4804 11024 4856 11076
rect 7012 11024 7064 11076
rect 8116 11024 8168 11076
rect 9864 11024 9916 11076
rect 14924 11024 14976 11076
rect 18236 11024 18288 11076
rect 18788 11024 18840 11076
rect 19156 11024 19208 11076
rect 25596 11024 25648 11076
rect 26240 11067 26292 11076
rect 26240 11033 26274 11067
rect 26274 11033 26292 11067
rect 26240 11024 26292 11033
rect 27712 11024 27764 11076
rect 30012 11024 30064 11076
rect 35164 11067 35216 11076
rect 35164 11033 35198 11067
rect 35198 11033 35216 11067
rect 35164 11024 35216 11033
rect 38292 11024 38344 11076
rect 5448 10956 5500 11008
rect 7840 10956 7892 11008
rect 22468 10956 22520 11008
rect 22928 10999 22980 11008
rect 22928 10965 22937 10999
rect 22937 10965 22971 10999
rect 22971 10965 22980 10999
rect 22928 10956 22980 10965
rect 23388 10999 23440 11008
rect 23388 10965 23397 10999
rect 23397 10965 23431 10999
rect 23431 10965 23440 10999
rect 23388 10956 23440 10965
rect 27344 10999 27396 11008
rect 27344 10965 27353 10999
rect 27353 10965 27387 10999
rect 27387 10965 27396 10999
rect 27344 10956 27396 10965
rect 28448 10999 28500 11008
rect 28448 10965 28457 10999
rect 28457 10965 28491 10999
rect 28491 10965 28500 10999
rect 28448 10956 28500 10965
rect 31024 10956 31076 11008
rect 38660 10999 38712 11008
rect 38660 10965 38669 10999
rect 38669 10965 38703 10999
rect 38703 10965 38712 10999
rect 38660 10956 38712 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 15660 10752 15712 10804
rect 15936 10752 15988 10804
rect 17040 10727 17092 10736
rect 17040 10693 17049 10727
rect 17049 10693 17083 10727
rect 17083 10693 17092 10727
rect 17040 10684 17092 10693
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 6736 10548 6788 10600
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 6184 10480 6236 10532
rect 13268 10548 13320 10600
rect 16212 10548 16264 10600
rect 23756 10752 23808 10804
rect 25780 10752 25832 10804
rect 26240 10752 26292 10804
rect 26424 10752 26476 10804
rect 22284 10684 22336 10736
rect 28448 10684 28500 10736
rect 22468 10659 22520 10668
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 22468 10616 22520 10625
rect 23388 10616 23440 10668
rect 22560 10548 22612 10600
rect 17132 10480 17184 10532
rect 23572 10480 23624 10532
rect 9772 10412 9824 10464
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 19340 10455 19392 10464
rect 19340 10421 19349 10455
rect 19349 10421 19383 10455
rect 19383 10421 19392 10455
rect 19340 10412 19392 10421
rect 25044 10616 25096 10668
rect 25228 10659 25280 10668
rect 25228 10625 25237 10659
rect 25237 10625 25271 10659
rect 25271 10625 25280 10659
rect 25228 10616 25280 10625
rect 25412 10659 25464 10668
rect 25412 10625 25421 10659
rect 25421 10625 25455 10659
rect 25455 10625 25464 10659
rect 25412 10616 25464 10625
rect 24952 10480 25004 10532
rect 25596 10659 25648 10668
rect 25596 10625 25605 10659
rect 25605 10625 25639 10659
rect 25639 10625 25648 10659
rect 25596 10616 25648 10625
rect 27436 10616 27488 10668
rect 27620 10659 27672 10668
rect 27620 10625 27629 10659
rect 27629 10625 27663 10659
rect 27663 10625 27672 10659
rect 27620 10616 27672 10625
rect 27804 10659 27856 10668
rect 27804 10625 27813 10659
rect 27813 10625 27847 10659
rect 27847 10625 27856 10659
rect 27804 10616 27856 10625
rect 27344 10548 27396 10600
rect 28080 10616 28132 10668
rect 30564 10752 30616 10804
rect 33968 10752 34020 10804
rect 31024 10727 31076 10736
rect 31024 10693 31033 10727
rect 31033 10693 31067 10727
rect 31067 10693 31076 10727
rect 31024 10684 31076 10693
rect 31300 10684 31352 10736
rect 31668 10684 31720 10736
rect 35164 10752 35216 10804
rect 34796 10616 34848 10668
rect 40408 10752 40460 10804
rect 36268 10684 36320 10736
rect 38660 10684 38712 10736
rect 30472 10548 30524 10600
rect 31208 10480 31260 10532
rect 26976 10455 27028 10464
rect 26976 10421 26985 10455
rect 26985 10421 27019 10455
rect 27019 10421 27028 10455
rect 26976 10412 27028 10421
rect 38292 10616 38344 10668
rect 38384 10548 38436 10600
rect 39120 10412 39172 10464
rect 58164 10455 58216 10464
rect 58164 10421 58173 10455
rect 58173 10421 58207 10455
rect 58207 10421 58216 10455
rect 58164 10412 58216 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5356 10208 5408 10260
rect 11060 10208 11112 10260
rect 13544 10208 13596 10260
rect 15844 10208 15896 10260
rect 17040 10208 17092 10260
rect 25412 10208 25464 10260
rect 33784 10208 33836 10260
rect 11980 10140 12032 10192
rect 12808 10140 12860 10192
rect 14740 10140 14792 10192
rect 25596 10140 25648 10192
rect 4068 10072 4120 10124
rect 4528 10072 4580 10124
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 2596 10004 2648 10056
rect 9772 10047 9824 10056
rect 4344 9936 4396 9988
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 10692 10072 10744 10124
rect 25320 10072 25372 10124
rect 11796 9936 11848 9988
rect 1400 9868 1452 9920
rect 6828 9911 6880 9920
rect 6828 9877 6837 9911
rect 6837 9877 6871 9911
rect 6871 9877 6880 9911
rect 6828 9868 6880 9877
rect 9220 9868 9272 9920
rect 9404 9868 9456 9920
rect 11704 9868 11756 9920
rect 12532 10004 12584 10056
rect 15844 10004 15896 10056
rect 12164 9979 12216 9988
rect 12164 9945 12173 9979
rect 12173 9945 12207 9979
rect 12207 9945 12216 9979
rect 22284 10004 22336 10056
rect 27344 10004 27396 10056
rect 27436 10004 27488 10056
rect 31760 10072 31812 10124
rect 12164 9936 12216 9945
rect 12808 9868 12860 9920
rect 12992 9868 13044 9920
rect 15384 9911 15436 9920
rect 15384 9877 15393 9911
rect 15393 9877 15427 9911
rect 15427 9877 15436 9911
rect 15384 9868 15436 9877
rect 15476 9868 15528 9920
rect 15936 9868 15988 9920
rect 26240 9936 26292 9988
rect 26976 9936 27028 9988
rect 30932 10004 30984 10056
rect 31208 10047 31260 10056
rect 31208 10013 31217 10047
rect 31217 10013 31251 10047
rect 31251 10013 31260 10047
rect 31208 10004 31260 10013
rect 31852 10004 31904 10056
rect 32036 10004 32088 10056
rect 32588 10047 32640 10056
rect 32588 10013 32597 10047
rect 32597 10013 32631 10047
rect 32631 10013 32640 10047
rect 32588 10004 32640 10013
rect 35624 10004 35676 10056
rect 37280 10004 37332 10056
rect 39396 10004 39448 10056
rect 31668 9936 31720 9988
rect 30380 9868 30432 9920
rect 30840 9868 30892 9920
rect 31484 9911 31536 9920
rect 31484 9877 31493 9911
rect 31493 9877 31527 9911
rect 31527 9877 31536 9911
rect 31484 9868 31536 9877
rect 32220 9868 32272 9920
rect 33140 9936 33192 9988
rect 38292 9936 38344 9988
rect 35440 9868 35492 9920
rect 38752 9911 38804 9920
rect 38752 9877 38761 9911
rect 38761 9877 38795 9911
rect 38795 9877 38804 9911
rect 38752 9868 38804 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 8208 9596 8260 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 3516 9528 3568 9580
rect 4344 9571 4396 9580
rect 4344 9537 4353 9571
rect 4353 9537 4387 9571
rect 4387 9537 4396 9571
rect 4344 9528 4396 9537
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 6736 9528 6788 9580
rect 9772 9664 9824 9716
rect 10232 9664 10284 9716
rect 10692 9664 10744 9716
rect 12164 9664 12216 9716
rect 13544 9664 13596 9716
rect 17040 9664 17092 9716
rect 19432 9664 19484 9716
rect 11428 9596 11480 9648
rect 15752 9596 15804 9648
rect 11704 9571 11756 9580
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 5724 9460 5776 9512
rect 7012 9460 7064 9512
rect 7288 9392 7340 9444
rect 8116 9392 8168 9444
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 11796 9528 11848 9580
rect 13360 9571 13412 9580
rect 13360 9537 13369 9571
rect 13369 9537 13403 9571
rect 13403 9537 13412 9571
rect 13360 9528 13412 9537
rect 14740 9528 14792 9580
rect 11980 9460 12032 9512
rect 15200 9460 15252 9512
rect 15384 9460 15436 9512
rect 18420 9528 18472 9580
rect 18972 9596 19024 9648
rect 20076 9596 20128 9648
rect 20536 9596 20588 9648
rect 20260 9528 20312 9580
rect 22928 9596 22980 9648
rect 28540 9664 28592 9716
rect 29184 9664 29236 9716
rect 31024 9664 31076 9716
rect 23572 9596 23624 9648
rect 24768 9596 24820 9648
rect 25044 9596 25096 9648
rect 29000 9596 29052 9648
rect 30932 9596 30984 9648
rect 39396 9664 39448 9716
rect 31668 9596 31720 9648
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 3976 9324 4028 9376
rect 6184 9324 6236 9376
rect 6920 9367 6972 9376
rect 6920 9333 6929 9367
rect 6929 9333 6963 9367
rect 6963 9333 6972 9367
rect 6920 9324 6972 9333
rect 7656 9324 7708 9376
rect 9404 9324 9456 9376
rect 13084 9324 13136 9376
rect 14464 9324 14516 9376
rect 15016 9324 15068 9376
rect 20352 9392 20404 9444
rect 23480 9571 23532 9580
rect 21824 9503 21876 9512
rect 21824 9469 21833 9503
rect 21833 9469 21867 9503
rect 21867 9469 21876 9503
rect 21824 9460 21876 9469
rect 22192 9460 22244 9512
rect 23480 9537 23489 9571
rect 23489 9537 23523 9571
rect 23523 9537 23532 9571
rect 23480 9528 23532 9537
rect 25228 9571 25280 9580
rect 25228 9537 25237 9571
rect 25237 9537 25271 9571
rect 25271 9537 25280 9571
rect 25228 9528 25280 9537
rect 25412 9571 25464 9580
rect 25412 9537 25421 9571
rect 25421 9537 25455 9571
rect 25455 9537 25464 9571
rect 25412 9528 25464 9537
rect 28080 9528 28132 9580
rect 23112 9392 23164 9444
rect 18420 9324 18472 9376
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 30380 9528 30432 9580
rect 31024 9571 31076 9580
rect 31024 9537 31033 9571
rect 31033 9537 31067 9571
rect 31067 9537 31076 9571
rect 31024 9528 31076 9537
rect 31208 9571 31260 9580
rect 31208 9537 31217 9571
rect 31217 9537 31251 9571
rect 31251 9537 31260 9571
rect 31208 9528 31260 9537
rect 25688 9392 25740 9444
rect 26056 9392 26108 9444
rect 28724 9392 28776 9444
rect 31116 9460 31168 9512
rect 31760 9528 31812 9580
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 32956 9596 33008 9648
rect 35348 9596 35400 9648
rect 38660 9571 38712 9580
rect 38660 9537 38694 9571
rect 38694 9537 38712 9571
rect 38660 9528 38712 9537
rect 32588 9460 32640 9512
rect 34704 9460 34756 9512
rect 37924 9460 37976 9512
rect 38384 9503 38436 9512
rect 38384 9469 38393 9503
rect 38393 9469 38427 9503
rect 38427 9469 38436 9503
rect 38384 9460 38436 9469
rect 31576 9435 31628 9444
rect 31576 9401 31585 9435
rect 31585 9401 31619 9435
rect 31619 9401 31628 9435
rect 31576 9392 31628 9401
rect 25412 9324 25464 9376
rect 30380 9324 30432 9376
rect 31300 9324 31352 9376
rect 33140 9324 33192 9376
rect 35624 9324 35676 9376
rect 37556 9324 37608 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2320 9120 2372 9172
rect 2964 9120 3016 9172
rect 13544 9163 13596 9172
rect 5172 9052 5224 9104
rect 3976 8984 4028 9036
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 3424 8848 3476 8900
rect 5540 8916 5592 8968
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 2780 8780 2832 8789
rect 3976 8780 4028 8832
rect 5632 8848 5684 8900
rect 6000 8984 6052 9036
rect 6184 8984 6236 9036
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 8484 9052 8536 9104
rect 7196 8984 7248 9036
rect 7288 8959 7340 8968
rect 5816 8848 5868 8900
rect 7288 8925 7297 8959
rect 7297 8925 7331 8959
rect 7331 8925 7340 8959
rect 7288 8916 7340 8925
rect 13544 9129 13553 9163
rect 13553 9129 13587 9163
rect 13587 9129 13596 9163
rect 13544 9120 13596 9129
rect 15476 9120 15528 9172
rect 16028 9120 16080 9172
rect 11428 9095 11480 9104
rect 11428 9061 11437 9095
rect 11437 9061 11471 9095
rect 11471 9061 11480 9095
rect 11428 9052 11480 9061
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 14004 8984 14056 9036
rect 19432 9120 19484 9172
rect 20352 9120 20404 9172
rect 20628 9163 20680 9172
rect 20628 9129 20637 9163
rect 20637 9129 20671 9163
rect 20671 9129 20680 9163
rect 20628 9120 20680 9129
rect 25228 9120 25280 9172
rect 27712 9163 27764 9172
rect 27712 9129 27721 9163
rect 27721 9129 27755 9163
rect 27755 9129 27764 9163
rect 27712 9120 27764 9129
rect 30104 9163 30156 9172
rect 30104 9129 30113 9163
rect 30113 9129 30147 9163
rect 30147 9129 30156 9163
rect 30104 9120 30156 9129
rect 32312 9120 32364 9172
rect 34244 9120 34296 9172
rect 35348 9120 35400 9172
rect 20260 9052 20312 9104
rect 24492 9052 24544 9104
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 14464 8916 14516 8968
rect 18328 8916 18380 8968
rect 21824 8984 21876 9036
rect 8300 8848 8352 8900
rect 11888 8848 11940 8900
rect 5264 8780 5316 8832
rect 6092 8823 6144 8832
rect 6092 8789 6101 8823
rect 6101 8789 6135 8823
rect 6135 8789 6144 8823
rect 6092 8780 6144 8789
rect 6184 8780 6236 8832
rect 11980 8780 12032 8832
rect 12164 8780 12216 8832
rect 17408 8848 17460 8900
rect 19064 8848 19116 8900
rect 20536 8916 20588 8968
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 21364 8916 21416 8968
rect 23480 8916 23532 8968
rect 27804 9052 27856 9104
rect 35440 9052 35492 9104
rect 28724 8984 28776 9036
rect 28080 8916 28132 8968
rect 24032 8848 24084 8900
rect 16580 8823 16632 8832
rect 16580 8789 16589 8823
rect 16589 8789 16623 8823
rect 16623 8789 16632 8823
rect 16580 8780 16632 8789
rect 18788 8780 18840 8832
rect 25964 8848 26016 8900
rect 27436 8891 27488 8900
rect 27436 8857 27445 8891
rect 27445 8857 27479 8891
rect 27479 8857 27488 8891
rect 28540 8916 28592 8968
rect 31208 8984 31260 9036
rect 32220 8984 32272 9036
rect 31300 8959 31352 8968
rect 31300 8925 31309 8959
rect 31309 8925 31343 8959
rect 31343 8925 31352 8959
rect 31300 8916 31352 8925
rect 32128 8959 32180 8968
rect 32128 8925 32137 8959
rect 32137 8925 32171 8959
rect 32171 8925 32180 8959
rect 32128 8916 32180 8925
rect 32404 8959 32456 8968
rect 32404 8925 32413 8959
rect 32413 8925 32447 8959
rect 32447 8925 32456 8959
rect 32404 8916 32456 8925
rect 32588 8916 32640 8968
rect 34796 8916 34848 8968
rect 35624 8959 35676 8968
rect 35624 8925 35633 8959
rect 35633 8925 35667 8959
rect 35667 8925 35676 8959
rect 35624 8916 35676 8925
rect 35808 8916 35860 8968
rect 27436 8848 27488 8857
rect 24492 8823 24544 8832
rect 24492 8789 24501 8823
rect 24501 8789 24535 8823
rect 24535 8789 24544 8823
rect 24492 8780 24544 8789
rect 25412 8780 25464 8832
rect 28080 8780 28132 8832
rect 31576 8848 31628 8900
rect 32220 8848 32272 8900
rect 37648 8984 37700 9036
rect 36912 8959 36964 8968
rect 36912 8925 36921 8959
rect 36921 8925 36955 8959
rect 36955 8925 36964 8959
rect 36912 8916 36964 8925
rect 37556 8959 37608 8968
rect 37556 8925 37565 8959
rect 37565 8925 37599 8959
rect 37599 8925 37608 8959
rect 37556 8916 37608 8925
rect 58164 8959 58216 8968
rect 58164 8925 58173 8959
rect 58173 8925 58207 8959
rect 58207 8925 58216 8959
rect 58164 8916 58216 8925
rect 37280 8848 37332 8900
rect 35348 8780 35400 8832
rect 37096 8823 37148 8832
rect 37096 8789 37105 8823
rect 37105 8789 37139 8823
rect 37139 8789 37148 8823
rect 37096 8780 37148 8789
rect 37924 8780 37976 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 1952 8576 2004 8628
rect 5632 8576 5684 8628
rect 5816 8619 5868 8628
rect 5816 8585 5825 8619
rect 5825 8585 5859 8619
rect 5859 8585 5868 8619
rect 5816 8576 5868 8585
rect 5908 8576 5960 8628
rect 8668 8576 8720 8628
rect 9588 8576 9640 8628
rect 9680 8576 9732 8628
rect 12992 8576 13044 8628
rect 13360 8576 13412 8628
rect 14004 8619 14056 8628
rect 14004 8585 14013 8619
rect 14013 8585 14047 8619
rect 14047 8585 14056 8619
rect 14004 8576 14056 8585
rect 15476 8576 15528 8628
rect 17408 8576 17460 8628
rect 3424 8508 3476 8560
rect 2044 8440 2096 8492
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3792 8440 3844 8492
rect 5816 8440 5868 8492
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 2044 8347 2096 8356
rect 2044 8313 2053 8347
rect 2053 8313 2087 8347
rect 2087 8313 2096 8347
rect 2044 8304 2096 8313
rect 5264 8304 5316 8356
rect 8392 8440 8444 8492
rect 9772 8440 9824 8492
rect 8024 8415 8076 8424
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 8208 8415 8260 8424
rect 8208 8381 8217 8415
rect 8217 8381 8251 8415
rect 8251 8381 8260 8415
rect 8208 8372 8260 8381
rect 12348 8508 12400 8560
rect 13084 8508 13136 8560
rect 16764 8551 16816 8560
rect 16764 8517 16773 8551
rect 16773 8517 16807 8551
rect 16807 8517 16816 8551
rect 16764 8508 16816 8517
rect 11796 8440 11848 8492
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 12624 8440 12676 8492
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 7656 8304 7708 8356
rect 13268 8372 13320 8424
rect 12256 8304 12308 8356
rect 12440 8304 12492 8356
rect 12992 8347 13044 8356
rect 12992 8313 13001 8347
rect 13001 8313 13035 8347
rect 13035 8313 13044 8347
rect 16028 8440 16080 8492
rect 17960 8576 18012 8628
rect 19064 8619 19116 8628
rect 19064 8585 19073 8619
rect 19073 8585 19107 8619
rect 19107 8585 19116 8619
rect 19064 8576 19116 8585
rect 21272 8576 21324 8628
rect 24492 8576 24544 8628
rect 28908 8619 28960 8628
rect 17960 8483 18012 8492
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 20628 8508 20680 8560
rect 17960 8440 18012 8449
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 18972 8440 19024 8492
rect 19984 8440 20036 8492
rect 24952 8508 25004 8560
rect 25504 8508 25556 8560
rect 24860 8483 24912 8492
rect 24860 8449 24869 8483
rect 24869 8449 24903 8483
rect 24903 8449 24912 8483
rect 24860 8440 24912 8449
rect 25136 8440 25188 8492
rect 19248 8372 19300 8424
rect 25688 8372 25740 8424
rect 28908 8585 28917 8619
rect 28917 8585 28951 8619
rect 28951 8585 28960 8619
rect 28908 8576 28960 8585
rect 30012 8576 30064 8628
rect 30196 8576 30248 8628
rect 30472 8576 30524 8628
rect 27436 8508 27488 8560
rect 28080 8508 28132 8560
rect 29000 8508 29052 8560
rect 37556 8576 37608 8628
rect 38660 8576 38712 8628
rect 34796 8551 34848 8560
rect 34796 8517 34805 8551
rect 34805 8517 34839 8551
rect 34839 8517 34848 8551
rect 34796 8508 34848 8517
rect 37096 8508 37148 8560
rect 38752 8508 38804 8560
rect 26240 8483 26292 8492
rect 26240 8449 26249 8483
rect 26249 8449 26283 8483
rect 26283 8449 26292 8483
rect 26240 8440 26292 8449
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 28724 8483 28776 8492
rect 28724 8449 28733 8483
rect 28733 8449 28767 8483
rect 28767 8449 28776 8483
rect 28724 8440 28776 8449
rect 31116 8483 31168 8492
rect 31116 8449 31125 8483
rect 31125 8449 31159 8483
rect 31159 8449 31168 8483
rect 31116 8440 31168 8449
rect 26424 8372 26476 8424
rect 12992 8304 13044 8313
rect 18696 8304 18748 8356
rect 25964 8304 26016 8356
rect 29552 8304 29604 8356
rect 37280 8440 37332 8492
rect 35532 8372 35584 8424
rect 37740 8483 37792 8492
rect 37740 8449 37749 8483
rect 37749 8449 37783 8483
rect 37783 8449 37792 8483
rect 37740 8440 37792 8449
rect 38844 8483 38896 8492
rect 38844 8449 38853 8483
rect 38853 8449 38887 8483
rect 38887 8449 38896 8483
rect 38844 8440 38896 8449
rect 38660 8372 38712 8424
rect 39120 8372 39172 8424
rect 34704 8304 34756 8356
rect 37924 8304 37976 8356
rect 39304 8440 39356 8492
rect 6736 8236 6788 8288
rect 6920 8236 6972 8288
rect 11520 8279 11572 8288
rect 11520 8245 11529 8279
rect 11529 8245 11563 8279
rect 11563 8245 11572 8279
rect 11520 8236 11572 8245
rect 16028 8279 16080 8288
rect 16028 8245 16037 8279
rect 16037 8245 16071 8279
rect 16071 8245 16080 8279
rect 16028 8236 16080 8245
rect 17684 8236 17736 8288
rect 18972 8236 19024 8288
rect 22928 8236 22980 8288
rect 25596 8236 25648 8288
rect 36084 8236 36136 8288
rect 38200 8236 38252 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 7472 8032 7524 8084
rect 8024 8032 8076 8084
rect 17684 8075 17736 8084
rect 2504 7896 2556 7948
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 6092 7828 6144 7880
rect 7012 7828 7064 7880
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 17960 8032 18012 8084
rect 19248 8075 19300 8084
rect 19248 8041 19257 8075
rect 19257 8041 19291 8075
rect 19291 8041 19300 8075
rect 19248 8032 19300 8041
rect 23204 8075 23256 8084
rect 23204 8041 23213 8075
rect 23213 8041 23247 8075
rect 23247 8041 23256 8075
rect 23204 8032 23256 8041
rect 24860 8032 24912 8084
rect 11888 7896 11940 7948
rect 11428 7828 11480 7880
rect 11704 7828 11756 7880
rect 13452 7896 13504 7948
rect 16856 7964 16908 8016
rect 18696 7896 18748 7948
rect 3056 7760 3108 7812
rect 6368 7760 6420 7812
rect 7288 7760 7340 7812
rect 11520 7760 11572 7812
rect 12164 7760 12216 7812
rect 15292 7828 15344 7880
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 19432 7871 19484 7880
rect 19432 7837 19441 7871
rect 19441 7837 19475 7871
rect 19475 7837 19484 7871
rect 19432 7828 19484 7837
rect 15384 7760 15436 7812
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 3700 7692 3752 7744
rect 7196 7692 7248 7744
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 8668 7692 8720 7744
rect 11796 7692 11848 7744
rect 12532 7692 12584 7744
rect 12624 7692 12676 7744
rect 13544 7692 13596 7744
rect 13912 7692 13964 7744
rect 19984 7760 20036 7812
rect 24124 7964 24176 8016
rect 27436 8032 27488 8084
rect 29000 8032 29052 8084
rect 36084 8075 36136 8084
rect 36084 8041 36093 8075
rect 36093 8041 36127 8075
rect 36127 8041 36136 8075
rect 36084 8032 36136 8041
rect 37280 8075 37332 8084
rect 37280 8041 37289 8075
rect 37289 8041 37323 8075
rect 37323 8041 37332 8075
rect 37280 8032 37332 8041
rect 36912 7964 36964 8016
rect 25688 7939 25740 7948
rect 22928 7871 22980 7880
rect 22928 7837 22937 7871
rect 22937 7837 22971 7871
rect 22971 7837 22980 7871
rect 22928 7828 22980 7837
rect 23204 7828 23256 7880
rect 25688 7905 25697 7939
rect 25697 7905 25731 7939
rect 25731 7905 25740 7939
rect 25688 7896 25740 7905
rect 37924 7939 37976 7948
rect 21732 7692 21784 7744
rect 22560 7760 22612 7812
rect 24308 7760 24360 7812
rect 26240 7828 26292 7880
rect 31484 7828 31536 7880
rect 33876 7828 33928 7880
rect 26056 7760 26108 7812
rect 25780 7692 25832 7744
rect 35624 7828 35676 7880
rect 35440 7760 35492 7812
rect 37924 7905 37933 7939
rect 37933 7905 37967 7939
rect 37967 7905 37976 7939
rect 37924 7896 37976 7905
rect 38200 7871 38252 7880
rect 38200 7837 38234 7871
rect 38234 7837 38252 7871
rect 38200 7828 38252 7837
rect 58164 7871 58216 7880
rect 58164 7837 58173 7871
rect 58173 7837 58207 7871
rect 58207 7837 58216 7871
rect 58164 7828 58216 7837
rect 38844 7760 38896 7812
rect 35716 7692 35768 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 5724 7352 5776 7404
rect 9680 7488 9732 7540
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 6920 7420 6972 7472
rect 8024 7352 8076 7404
rect 9772 7420 9824 7472
rect 8392 7352 8444 7404
rect 11888 7488 11940 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 15660 7488 15712 7540
rect 15292 7420 15344 7472
rect 16856 7463 16908 7472
rect 16856 7429 16865 7463
rect 16865 7429 16899 7463
rect 16899 7429 16908 7463
rect 16856 7420 16908 7429
rect 17316 7420 17368 7472
rect 5632 7284 5684 7336
rect 5816 7327 5868 7336
rect 5816 7293 5825 7327
rect 5825 7293 5859 7327
rect 5859 7293 5868 7327
rect 5816 7284 5868 7293
rect 6460 7327 6512 7336
rect 6460 7293 6469 7327
rect 6469 7293 6503 7327
rect 6503 7293 6512 7327
rect 6460 7284 6512 7293
rect 6736 7327 6788 7336
rect 6736 7293 6745 7327
rect 6745 7293 6779 7327
rect 6779 7293 6788 7327
rect 6736 7284 6788 7293
rect 11336 7284 11388 7336
rect 11612 7352 11664 7404
rect 7840 7216 7892 7268
rect 15016 7216 15068 7268
rect 16764 7216 16816 7268
rect 18696 7352 18748 7404
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 23296 7488 23348 7540
rect 24216 7488 24268 7540
rect 26056 7531 26108 7540
rect 23848 7420 23900 7472
rect 24400 7420 24452 7472
rect 26056 7497 26065 7531
rect 26065 7497 26099 7531
rect 26099 7497 26108 7531
rect 26056 7488 26108 7497
rect 27712 7488 27764 7540
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 23204 7352 23256 7404
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 25136 7352 25188 7404
rect 25596 7395 25648 7404
rect 25596 7361 25605 7395
rect 25605 7361 25639 7395
rect 25639 7361 25648 7395
rect 25596 7352 25648 7361
rect 25504 7284 25556 7336
rect 25964 7352 26016 7404
rect 19984 7216 20036 7268
rect 27620 7352 27672 7404
rect 28356 7352 28408 7404
rect 31024 7420 31076 7472
rect 31208 7352 31260 7404
rect 33140 7420 33192 7472
rect 35440 7420 35492 7472
rect 38844 7463 38896 7472
rect 38844 7429 38853 7463
rect 38853 7429 38887 7463
rect 38887 7429 38896 7463
rect 38844 7420 38896 7429
rect 33876 7395 33928 7404
rect 33876 7361 33885 7395
rect 33885 7361 33919 7395
rect 33919 7361 33928 7395
rect 33876 7352 33928 7361
rect 31576 7216 31628 7268
rect 1768 7191 1820 7200
rect 1768 7157 1777 7191
rect 1777 7157 1811 7191
rect 1811 7157 1820 7191
rect 1768 7148 1820 7157
rect 3148 7148 3200 7200
rect 3976 7148 4028 7200
rect 7748 7148 7800 7200
rect 9220 7148 9272 7200
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 14280 7148 14332 7200
rect 14740 7148 14792 7200
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 17960 7148 18012 7200
rect 19340 7191 19392 7200
rect 19340 7157 19349 7191
rect 19349 7157 19383 7191
rect 19383 7157 19392 7191
rect 19340 7148 19392 7157
rect 23480 7191 23532 7200
rect 23480 7157 23489 7191
rect 23489 7157 23523 7191
rect 23523 7157 23532 7191
rect 23480 7148 23532 7157
rect 24584 7148 24636 7200
rect 25964 7148 26016 7200
rect 27988 7148 28040 7200
rect 29828 7148 29880 7200
rect 30932 7148 30984 7200
rect 35256 7395 35308 7404
rect 35256 7361 35265 7395
rect 35265 7361 35299 7395
rect 35299 7361 35308 7395
rect 35256 7352 35308 7361
rect 35532 7395 35584 7404
rect 35532 7361 35541 7395
rect 35541 7361 35575 7395
rect 35575 7361 35584 7395
rect 35532 7352 35584 7361
rect 35716 7352 35768 7404
rect 36268 7395 36320 7404
rect 36268 7361 36277 7395
rect 36277 7361 36311 7395
rect 36311 7361 36320 7395
rect 36268 7352 36320 7361
rect 37096 7352 37148 7404
rect 38292 7352 38344 7404
rect 36912 7284 36964 7336
rect 36176 7216 36228 7268
rect 34796 7148 34848 7200
rect 38936 7148 38988 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2504 6944 2556 6996
rect 3240 6944 3292 6996
rect 15384 6987 15436 6996
rect 15384 6953 15393 6987
rect 15393 6953 15427 6987
rect 15427 6953 15436 6987
rect 15384 6944 15436 6953
rect 27620 6987 27672 6996
rect 27620 6953 27629 6987
rect 27629 6953 27663 6987
rect 27663 6953 27672 6987
rect 27620 6944 27672 6953
rect 3884 6876 3936 6928
rect 2596 6808 2648 6860
rect 4068 6808 4120 6860
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 3884 6740 3936 6792
rect 5540 6808 5592 6860
rect 6736 6808 6788 6860
rect 3608 6672 3660 6724
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 3332 6604 3384 6656
rect 3424 6604 3476 6656
rect 6368 6740 6420 6792
rect 7196 6740 7248 6792
rect 7840 6740 7892 6792
rect 9864 6876 9916 6928
rect 9220 6851 9272 6860
rect 9220 6817 9229 6851
rect 9229 6817 9263 6851
rect 9263 6817 9272 6851
rect 9220 6808 9272 6817
rect 5080 6672 5132 6724
rect 5816 6672 5868 6724
rect 8300 6672 8352 6724
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 11060 6740 11112 6792
rect 15200 6808 15252 6860
rect 12256 6672 12308 6724
rect 12532 6740 12584 6792
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 16672 6808 16724 6860
rect 17040 6808 17092 6860
rect 19432 6808 19484 6860
rect 22192 6851 22244 6860
rect 22192 6817 22201 6851
rect 22201 6817 22235 6851
rect 22235 6817 22244 6851
rect 22192 6808 22244 6817
rect 16028 6783 16080 6792
rect 12624 6672 12676 6724
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 18788 6740 18840 6792
rect 21824 6740 21876 6792
rect 23480 6876 23532 6928
rect 30932 6944 30984 6996
rect 31024 6944 31076 6996
rect 36912 6987 36964 6996
rect 36912 6953 36921 6987
rect 36921 6953 36955 6987
rect 36955 6953 36964 6987
rect 36912 6944 36964 6953
rect 15936 6672 15988 6724
rect 18328 6672 18380 6724
rect 20168 6672 20220 6724
rect 23756 6740 23808 6792
rect 25136 6808 25188 6860
rect 25780 6851 25832 6860
rect 25780 6817 25789 6851
rect 25789 6817 25823 6851
rect 25823 6817 25832 6851
rect 25780 6808 25832 6817
rect 24584 6783 24636 6792
rect 24584 6749 24593 6783
rect 24593 6749 24627 6783
rect 24627 6749 24636 6783
rect 24584 6740 24636 6749
rect 24768 6783 24820 6792
rect 24768 6749 24777 6783
rect 24777 6749 24811 6783
rect 24811 6749 24820 6783
rect 27252 6808 27304 6860
rect 24768 6740 24820 6749
rect 27436 6740 27488 6792
rect 30012 6851 30064 6860
rect 30012 6817 30021 6851
rect 30021 6817 30055 6851
rect 30055 6817 30064 6851
rect 30012 6808 30064 6817
rect 37004 6876 37056 6928
rect 35440 6808 35492 6860
rect 38384 6808 38436 6860
rect 38660 6808 38712 6860
rect 25504 6672 25556 6724
rect 27528 6672 27580 6724
rect 30380 6672 30432 6724
rect 6644 6647 6696 6656
rect 6644 6613 6653 6647
rect 6653 6613 6687 6647
rect 6687 6613 6696 6647
rect 6644 6604 6696 6613
rect 6828 6604 6880 6656
rect 8024 6604 8076 6656
rect 8944 6604 8996 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 11520 6604 11572 6656
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 16856 6604 16908 6656
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 20720 6647 20772 6656
rect 20720 6613 20729 6647
rect 20729 6613 20763 6647
rect 20763 6613 20772 6647
rect 20720 6604 20772 6613
rect 20996 6604 21048 6656
rect 23572 6604 23624 6656
rect 25044 6647 25096 6656
rect 25044 6613 25053 6647
rect 25053 6613 25087 6647
rect 25087 6613 25096 6647
rect 25044 6604 25096 6613
rect 27068 6647 27120 6656
rect 27068 6613 27077 6647
rect 27077 6613 27111 6647
rect 27111 6613 27120 6647
rect 27068 6604 27120 6613
rect 30656 6604 30708 6656
rect 31116 6604 31168 6656
rect 34612 6604 34664 6656
rect 35532 6740 35584 6792
rect 35992 6783 36044 6792
rect 35992 6749 36001 6783
rect 36001 6749 36035 6783
rect 36035 6749 36044 6783
rect 35992 6740 36044 6749
rect 35900 6672 35952 6724
rect 36176 6783 36228 6792
rect 36176 6749 36185 6783
rect 36185 6749 36219 6783
rect 36219 6749 36228 6783
rect 36176 6740 36228 6749
rect 37004 6740 37056 6792
rect 37096 6715 37148 6724
rect 37096 6681 37105 6715
rect 37105 6681 37139 6715
rect 37139 6681 37148 6715
rect 37096 6672 37148 6681
rect 37372 6672 37424 6724
rect 38936 6783 38988 6792
rect 38936 6749 38945 6783
rect 38945 6749 38979 6783
rect 38979 6749 38988 6783
rect 38936 6740 38988 6749
rect 39304 6740 39356 6792
rect 35348 6604 35400 6656
rect 36084 6604 36136 6656
rect 38568 6604 38620 6656
rect 39304 6604 39356 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 11244 6400 11296 6452
rect 14832 6400 14884 6452
rect 3240 6375 3292 6384
rect 3240 6341 3249 6375
rect 3249 6341 3283 6375
rect 3283 6341 3292 6375
rect 3240 6332 3292 6341
rect 3332 6332 3384 6384
rect 6552 6332 6604 6384
rect 2136 6264 2188 6316
rect 6276 6264 6328 6316
rect 5356 6196 5408 6248
rect 7288 6264 7340 6316
rect 8024 6264 8076 6316
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 11428 6332 11480 6384
rect 9680 6264 9732 6316
rect 4712 6128 4764 6180
rect 8392 6128 8444 6180
rect 1676 6103 1728 6112
rect 1676 6069 1685 6103
rect 1685 6069 1719 6103
rect 1719 6069 1728 6103
rect 1676 6060 1728 6069
rect 2228 6103 2280 6112
rect 2228 6069 2237 6103
rect 2237 6069 2271 6103
rect 2271 6069 2280 6103
rect 2228 6060 2280 6069
rect 2688 6060 2740 6112
rect 4620 6060 4672 6112
rect 5632 6103 5684 6112
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 7564 6060 7616 6112
rect 9036 6060 9088 6112
rect 12900 6196 12952 6248
rect 13084 6332 13136 6384
rect 15568 6332 15620 6384
rect 17316 6400 17368 6452
rect 20536 6400 20588 6452
rect 21916 6400 21968 6452
rect 23664 6443 23716 6452
rect 23664 6409 23673 6443
rect 23673 6409 23707 6443
rect 23707 6409 23716 6443
rect 23664 6400 23716 6409
rect 24032 6400 24084 6452
rect 24768 6400 24820 6452
rect 25136 6443 25188 6452
rect 25136 6409 25145 6443
rect 25145 6409 25179 6443
rect 25179 6409 25188 6443
rect 25136 6400 25188 6409
rect 25688 6400 25740 6452
rect 27528 6443 27580 6452
rect 27528 6409 27537 6443
rect 27537 6409 27571 6443
rect 27571 6409 27580 6443
rect 27528 6400 27580 6409
rect 29184 6443 29236 6452
rect 29184 6409 29193 6443
rect 29193 6409 29227 6443
rect 29227 6409 29236 6443
rect 29184 6400 29236 6409
rect 30104 6400 30156 6452
rect 30380 6443 30432 6452
rect 30380 6409 30389 6443
rect 30389 6409 30423 6443
rect 30423 6409 30432 6443
rect 30380 6400 30432 6409
rect 37096 6400 37148 6452
rect 38844 6400 38896 6452
rect 17040 6375 17092 6384
rect 17040 6341 17049 6375
rect 17049 6341 17083 6375
rect 17083 6341 17092 6375
rect 17040 6332 17092 6341
rect 19340 6332 19392 6384
rect 14464 6264 14516 6316
rect 14648 6264 14700 6316
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 19432 6307 19484 6316
rect 19432 6273 19441 6307
rect 19441 6273 19475 6307
rect 19475 6273 19484 6307
rect 19432 6264 19484 6273
rect 19524 6264 19576 6316
rect 22560 6332 22612 6384
rect 24400 6332 24452 6384
rect 27068 6332 27120 6384
rect 27436 6332 27488 6384
rect 13728 6128 13780 6180
rect 11060 6060 11112 6112
rect 11428 6060 11480 6112
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 12992 6060 13044 6112
rect 13452 6103 13504 6112
rect 13452 6069 13461 6103
rect 13461 6069 13495 6103
rect 13495 6069 13504 6103
rect 13452 6060 13504 6069
rect 18420 6196 18472 6248
rect 18604 6196 18656 6248
rect 19248 6196 19300 6248
rect 21824 6239 21876 6248
rect 21824 6205 21833 6239
rect 21833 6205 21867 6239
rect 21867 6205 21876 6239
rect 21824 6196 21876 6205
rect 18512 6128 18564 6180
rect 23204 6264 23256 6316
rect 26976 6307 27028 6316
rect 26976 6273 26985 6307
rect 26985 6273 27019 6307
rect 27019 6273 27028 6307
rect 26976 6264 27028 6273
rect 27988 6307 28040 6316
rect 27988 6273 27997 6307
rect 27997 6273 28031 6307
rect 28031 6273 28040 6307
rect 27988 6264 28040 6273
rect 28172 6307 28224 6316
rect 28172 6273 28181 6307
rect 28181 6273 28215 6307
rect 28215 6273 28224 6307
rect 28172 6264 28224 6273
rect 29828 6264 29880 6316
rect 30104 6307 30156 6316
rect 30104 6273 30133 6307
rect 30133 6273 30156 6307
rect 31208 6307 31260 6316
rect 30104 6264 30156 6273
rect 31208 6273 31217 6307
rect 31217 6273 31251 6307
rect 31251 6273 31260 6307
rect 31208 6264 31260 6273
rect 34796 6332 34848 6384
rect 36176 6332 36228 6384
rect 32036 6264 32088 6316
rect 34704 6307 34756 6316
rect 34704 6273 34713 6307
rect 34713 6273 34747 6307
rect 34747 6273 34756 6307
rect 34704 6264 34756 6273
rect 36084 6264 36136 6316
rect 38660 6332 38712 6384
rect 37924 6264 37976 6316
rect 38568 6307 38620 6316
rect 38568 6273 38602 6307
rect 38602 6273 38620 6307
rect 38568 6264 38620 6273
rect 30104 6128 30156 6180
rect 14924 6060 14976 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 18236 6060 18288 6112
rect 20260 6103 20312 6112
rect 20260 6069 20269 6103
rect 20269 6069 20303 6103
rect 20303 6069 20312 6103
rect 20260 6060 20312 6069
rect 20812 6103 20864 6112
rect 20812 6069 20821 6103
rect 20821 6069 20855 6103
rect 20855 6069 20864 6103
rect 20812 6060 20864 6069
rect 30012 6060 30064 6112
rect 58164 6171 58216 6180
rect 58164 6137 58173 6171
rect 58173 6137 58207 6171
rect 58207 6137 58216 6171
rect 58164 6128 58216 6137
rect 30380 6060 30432 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 4068 5856 4120 5908
rect 2872 5720 2924 5772
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 2504 5652 2556 5704
rect 3332 5652 3384 5704
rect 3884 5652 3936 5704
rect 7656 5856 7708 5908
rect 8116 5856 8168 5908
rect 14464 5899 14516 5908
rect 6184 5788 6236 5840
rect 6552 5788 6604 5840
rect 8208 5788 8260 5840
rect 5724 5720 5776 5772
rect 8668 5720 8720 5772
rect 4712 5652 4764 5704
rect 5816 5652 5868 5704
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6736 5652 6788 5704
rect 7748 5652 7800 5704
rect 8300 5652 8352 5704
rect 8944 5652 8996 5704
rect 14464 5865 14473 5899
rect 14473 5865 14507 5899
rect 14507 5865 14516 5899
rect 14464 5856 14516 5865
rect 12900 5788 12952 5840
rect 18144 5856 18196 5908
rect 16672 5788 16724 5840
rect 18328 5788 18380 5840
rect 14648 5720 14700 5772
rect 10508 5652 10560 5704
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11612 5652 11664 5704
rect 12440 5652 12492 5704
rect 13268 5652 13320 5704
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 15752 5720 15804 5772
rect 1676 5584 1728 5636
rect 7932 5584 7984 5636
rect 10876 5584 10928 5636
rect 15292 5652 15344 5704
rect 16028 5720 16080 5772
rect 15936 5584 15988 5636
rect 16120 5584 16172 5636
rect 16672 5695 16724 5704
rect 16672 5661 16681 5695
rect 16681 5661 16715 5695
rect 16715 5661 16724 5695
rect 16672 5652 16724 5661
rect 18052 5695 18104 5704
rect 18052 5661 18061 5695
rect 18061 5661 18095 5695
rect 18095 5661 18104 5695
rect 18052 5652 18104 5661
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 19432 5856 19484 5908
rect 23756 5856 23808 5908
rect 29920 5856 29972 5908
rect 30564 5856 30616 5908
rect 33876 5899 33928 5908
rect 33876 5865 33885 5899
rect 33885 5865 33919 5899
rect 33919 5865 33928 5899
rect 33876 5856 33928 5865
rect 35348 5856 35400 5908
rect 35992 5899 36044 5908
rect 35992 5865 36001 5899
rect 36001 5865 36035 5899
rect 36035 5865 36044 5899
rect 35992 5856 36044 5865
rect 27804 5788 27856 5840
rect 30196 5788 30248 5840
rect 18788 5652 18840 5704
rect 19248 5695 19300 5704
rect 19248 5661 19257 5695
rect 19257 5661 19291 5695
rect 19291 5661 19300 5695
rect 19248 5652 19300 5661
rect 27344 5720 27396 5772
rect 30012 5720 30064 5772
rect 25412 5652 25464 5704
rect 4620 5516 4672 5568
rect 5356 5516 5408 5568
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 6184 5516 6236 5568
rect 6552 5516 6604 5568
rect 8116 5516 8168 5568
rect 8484 5516 8536 5568
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 9036 5516 9088 5568
rect 15476 5516 15528 5568
rect 18512 5584 18564 5636
rect 23848 5584 23900 5636
rect 27712 5695 27764 5704
rect 27712 5661 27721 5695
rect 27721 5661 27755 5695
rect 27755 5661 27764 5695
rect 30104 5695 30156 5704
rect 27712 5652 27764 5661
rect 30104 5661 30113 5695
rect 30113 5661 30147 5695
rect 30147 5661 30156 5695
rect 30104 5652 30156 5661
rect 30196 5652 30248 5704
rect 19340 5516 19392 5568
rect 21640 5559 21692 5568
rect 21640 5525 21649 5559
rect 21649 5525 21683 5559
rect 21683 5525 21692 5559
rect 21640 5516 21692 5525
rect 22192 5559 22244 5568
rect 22192 5525 22201 5559
rect 22201 5525 22235 5559
rect 22235 5525 22244 5559
rect 22192 5516 22244 5525
rect 22652 5559 22704 5568
rect 22652 5525 22661 5559
rect 22661 5525 22695 5559
rect 22695 5525 22704 5559
rect 22652 5516 22704 5525
rect 23204 5559 23256 5568
rect 23204 5525 23213 5559
rect 23213 5525 23247 5559
rect 23247 5525 23256 5559
rect 23204 5516 23256 5525
rect 24308 5516 24360 5568
rect 27436 5516 27488 5568
rect 28172 5584 28224 5636
rect 30656 5652 30708 5704
rect 31668 5652 31720 5704
rect 35624 5652 35676 5704
rect 36268 5652 36320 5704
rect 38292 5652 38344 5704
rect 30564 5584 30616 5636
rect 31208 5627 31260 5636
rect 31208 5593 31217 5627
rect 31217 5593 31251 5627
rect 31251 5593 31260 5627
rect 31208 5584 31260 5593
rect 32128 5584 32180 5636
rect 28540 5516 28592 5568
rect 29552 5559 29604 5568
rect 29552 5525 29561 5559
rect 29561 5525 29595 5559
rect 29595 5525 29604 5559
rect 29552 5516 29604 5525
rect 29920 5516 29972 5568
rect 31116 5516 31168 5568
rect 37372 5516 37424 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 2320 5312 2372 5364
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 4620 5312 4672 5364
rect 5080 5312 5132 5364
rect 5540 5312 5592 5364
rect 21824 5312 21876 5364
rect 25412 5355 25464 5364
rect 25412 5321 25421 5355
rect 25421 5321 25455 5355
rect 25455 5321 25464 5355
rect 25412 5312 25464 5321
rect 2228 5244 2280 5296
rect 2780 5219 2832 5228
rect 2780 5185 2789 5219
rect 2789 5185 2823 5219
rect 2823 5185 2832 5219
rect 3700 5219 3752 5228
rect 2780 5176 2832 5185
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 6000 5244 6052 5296
rect 8852 5244 8904 5296
rect 9772 5244 9824 5296
rect 5356 5176 5408 5228
rect 5448 5176 5500 5228
rect 6092 5176 6144 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 3516 5108 3568 5160
rect 7656 5108 7708 5160
rect 8484 5176 8536 5228
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 8116 5108 8168 5160
rect 14280 5176 14332 5228
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 15292 5219 15344 5228
rect 15292 5185 15301 5219
rect 15301 5185 15335 5219
rect 15335 5185 15344 5219
rect 15292 5176 15344 5185
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 15936 5244 15988 5296
rect 13452 5108 13504 5160
rect 18052 5176 18104 5228
rect 19432 5244 19484 5296
rect 18328 5108 18380 5160
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 21364 5176 21416 5228
rect 21088 5108 21140 5160
rect 29092 5312 29144 5364
rect 29736 5355 29788 5364
rect 29736 5321 29745 5355
rect 29745 5321 29779 5355
rect 29779 5321 29788 5355
rect 29736 5312 29788 5321
rect 26424 5287 26476 5296
rect 26424 5253 26433 5287
rect 26433 5253 26467 5287
rect 26467 5253 26476 5287
rect 26424 5244 26476 5253
rect 27896 5244 27948 5296
rect 27436 5219 27488 5228
rect 27436 5185 27445 5219
rect 27445 5185 27479 5219
rect 27479 5185 27488 5219
rect 27436 5176 27488 5185
rect 28172 5176 28224 5228
rect 30104 5176 30156 5228
rect 30380 5219 30432 5228
rect 30380 5185 30389 5219
rect 30389 5185 30423 5219
rect 30423 5185 30432 5219
rect 30380 5176 30432 5185
rect 30748 5312 30800 5364
rect 31668 5312 31720 5364
rect 36268 5312 36320 5364
rect 37924 5244 37976 5296
rect 30012 5108 30064 5160
rect 38384 5219 38436 5228
rect 38384 5185 38402 5219
rect 38402 5185 38436 5219
rect 38384 5176 38436 5185
rect 53748 5108 53800 5160
rect 5724 5083 5776 5092
rect 5724 5049 5733 5083
rect 5733 5049 5767 5083
rect 5767 5049 5776 5083
rect 5724 5040 5776 5049
rect 6552 5040 6604 5092
rect 3516 4972 3568 5024
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 6736 4972 6788 5024
rect 16948 5040 17000 5092
rect 19432 5040 19484 5092
rect 22100 5040 22152 5092
rect 27344 5040 27396 5092
rect 54116 5040 54168 5092
rect 10232 4972 10284 5024
rect 10784 4972 10836 5024
rect 11336 4972 11388 5024
rect 11888 4972 11940 5024
rect 13820 4972 13872 5024
rect 14096 5015 14148 5024
rect 14096 4981 14105 5015
rect 14105 4981 14139 5015
rect 14139 4981 14148 5015
rect 14096 4972 14148 4981
rect 14740 5015 14792 5024
rect 14740 4981 14749 5015
rect 14749 4981 14783 5015
rect 14783 4981 14792 5015
rect 14740 4972 14792 4981
rect 16764 4972 16816 5024
rect 18420 4972 18472 5024
rect 20076 4972 20128 5024
rect 20904 4972 20956 5024
rect 21732 4972 21784 5024
rect 22560 4972 22612 5024
rect 23480 4972 23532 5024
rect 27252 4972 27304 5024
rect 30840 5015 30892 5024
rect 30840 4981 30849 5015
rect 30849 4981 30883 5015
rect 30883 4981 30892 5015
rect 30840 4972 30892 4981
rect 53656 4972 53708 5024
rect 58164 5015 58216 5024
rect 58164 4981 58173 5015
rect 58173 4981 58207 5015
rect 58207 4981 58216 5015
rect 58164 4972 58216 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 5908 4700 5960 4752
rect 6092 4811 6144 4820
rect 6092 4777 6101 4811
rect 6101 4777 6135 4811
rect 6135 4777 6144 4811
rect 7472 4811 7524 4820
rect 6092 4768 6144 4777
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 8116 4768 8168 4820
rect 7012 4700 7064 4752
rect 9404 4811 9456 4820
rect 9404 4777 9413 4811
rect 9413 4777 9447 4811
rect 9447 4777 9456 4811
rect 9404 4768 9456 4777
rect 9772 4768 9824 4820
rect 23848 4768 23900 4820
rect 24400 4811 24452 4820
rect 24400 4777 24409 4811
rect 24409 4777 24443 4811
rect 24443 4777 24452 4811
rect 24400 4768 24452 4777
rect 9864 4700 9916 4752
rect 10140 4700 10192 4752
rect 18144 4700 18196 4752
rect 22008 4700 22060 4752
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 5724 4632 5776 4684
rect 5264 4564 5316 4616
rect 5540 4564 5592 4616
rect 8484 4632 8536 4684
rect 10416 4632 10468 4684
rect 13452 4632 13504 4684
rect 18972 4632 19024 4684
rect 46756 4768 46808 4820
rect 32128 4700 32180 4752
rect 52184 4700 52236 4752
rect 53932 4700 53984 4752
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 6736 4564 6788 4616
rect 7564 4607 7616 4616
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 6552 4496 6604 4548
rect 6828 4496 6880 4548
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 9128 4564 9180 4616
rect 2780 4428 2832 4437
rect 5264 4428 5316 4480
rect 6920 4428 6972 4480
rect 10968 4564 11020 4616
rect 12164 4564 12216 4616
rect 12992 4564 13044 4616
rect 13912 4564 13964 4616
rect 14188 4564 14240 4616
rect 15384 4564 15436 4616
rect 16028 4564 16080 4616
rect 16488 4564 16540 4616
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 19156 4564 19208 4616
rect 19340 4564 19392 4616
rect 20628 4564 20680 4616
rect 21180 4564 21232 4616
rect 22284 4564 22336 4616
rect 23572 4607 23624 4616
rect 23572 4573 23590 4607
rect 23590 4573 23624 4607
rect 23572 4564 23624 4573
rect 10600 4496 10652 4548
rect 10876 4539 10928 4548
rect 10876 4505 10885 4539
rect 10885 4505 10919 4539
rect 10919 4505 10928 4539
rect 10876 4496 10928 4505
rect 22376 4496 22428 4548
rect 53196 4632 53248 4684
rect 54300 4632 54352 4684
rect 25136 4564 25188 4616
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 30932 4564 30984 4616
rect 31116 4564 31168 4616
rect 52092 4564 52144 4616
rect 52644 4564 52696 4616
rect 25044 4496 25096 4548
rect 14004 4428 14056 4480
rect 18328 4428 18380 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 3608 4224 3660 4276
rect 4068 4224 4120 4276
rect 6276 4224 6328 4276
rect 7104 4224 7156 4276
rect 9404 4224 9456 4276
rect 29736 4224 29788 4276
rect 3884 4156 3936 4208
rect 6552 4199 6604 4208
rect 6552 4165 6561 4199
rect 6561 4165 6595 4199
rect 6595 4165 6604 4199
rect 6552 4156 6604 4165
rect 1768 4088 1820 4140
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 3792 4088 3844 4140
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 4620 4088 4672 4140
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 3240 3884 3292 3936
rect 4620 3884 4672 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 7472 4088 7524 4140
rect 6828 4020 6880 4072
rect 7380 4020 7432 4072
rect 8392 4063 8444 4072
rect 5080 3884 5132 3936
rect 5540 3884 5592 3936
rect 7472 3952 7524 4004
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8576 4063 8628 4072
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 9956 4088 10008 4140
rect 11520 4088 11572 4140
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 10416 4063 10468 4072
rect 10416 4029 10425 4063
rect 10425 4029 10459 4063
rect 10459 4029 10468 4063
rect 10968 4063 11020 4072
rect 10416 4020 10468 4029
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 8300 3995 8352 4004
rect 8300 3961 8309 3995
rect 8309 3961 8343 3995
rect 8343 3961 8352 3995
rect 8300 3952 8352 3961
rect 10600 3995 10652 4004
rect 10600 3961 10609 3995
rect 10609 3961 10643 3995
rect 10643 3961 10652 3995
rect 10600 3952 10652 3961
rect 10692 3952 10744 4004
rect 12256 4088 12308 4140
rect 14280 4088 14332 4140
rect 15568 4088 15620 4140
rect 16948 4131 17000 4140
rect 16948 4097 16982 4131
rect 16982 4097 17000 4131
rect 16948 4088 17000 4097
rect 19432 4156 19484 4208
rect 27252 4199 27304 4208
rect 19248 4088 19300 4140
rect 27252 4165 27286 4199
rect 27286 4165 27304 4199
rect 27252 4156 27304 4165
rect 25780 4088 25832 4140
rect 30932 4088 30984 4140
rect 33876 4088 33928 4140
rect 34704 4088 34756 4140
rect 53012 4088 53064 4140
rect 16212 4020 16264 4072
rect 51816 4020 51868 4072
rect 54024 4020 54076 4072
rect 6644 3884 6696 3936
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 7564 3884 7616 3936
rect 8484 3884 8536 3936
rect 9036 3884 9088 3936
rect 9128 3884 9180 3936
rect 10140 3884 10192 3936
rect 11980 3884 12032 3936
rect 13176 3884 13228 3936
rect 13544 3927 13596 3936
rect 13544 3893 13553 3927
rect 13553 3893 13587 3927
rect 13587 3893 13596 3927
rect 13544 3884 13596 3893
rect 15200 3952 15252 4004
rect 16672 3952 16724 4004
rect 18512 3952 18564 4004
rect 21364 3952 21416 4004
rect 22468 3952 22520 4004
rect 28540 3952 28592 4004
rect 35624 3952 35676 4004
rect 52828 3952 52880 4004
rect 15936 3884 15988 3936
rect 17684 3884 17736 3936
rect 19432 3884 19484 3936
rect 22928 3884 22980 3936
rect 23112 3884 23164 3936
rect 23388 3884 23440 3936
rect 24216 3884 24268 3936
rect 25504 3927 25556 3936
rect 25504 3893 25513 3927
rect 25513 3893 25547 3927
rect 25547 3893 25556 3927
rect 25504 3884 25556 3893
rect 51080 3884 51132 3936
rect 51356 3884 51408 3936
rect 52460 3884 52512 3936
rect 55312 3927 55364 3936
rect 55312 3893 55321 3927
rect 55321 3893 55355 3927
rect 55355 3893 55364 3927
rect 55312 3884 55364 3893
rect 58440 3884 58492 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4804 3680 4856 3732
rect 7012 3680 7064 3732
rect 8300 3680 8352 3732
rect 9312 3680 9364 3732
rect 9772 3723 9824 3732
rect 9772 3689 9781 3723
rect 9781 3689 9815 3723
rect 9815 3689 9824 3723
rect 9772 3680 9824 3689
rect 12072 3680 12124 3732
rect 14648 3680 14700 3732
rect 17040 3723 17092 3732
rect 17040 3689 17049 3723
rect 17049 3689 17083 3723
rect 17083 3689 17092 3723
rect 17040 3680 17092 3689
rect 18880 3680 18932 3732
rect 20444 3680 20496 3732
rect 21088 3723 21140 3732
rect 21088 3689 21097 3723
rect 21097 3689 21131 3723
rect 21131 3689 21140 3723
rect 21088 3680 21140 3689
rect 21916 3723 21968 3732
rect 21916 3689 21925 3723
rect 21925 3689 21959 3723
rect 21959 3689 21968 3723
rect 21916 3680 21968 3689
rect 32036 3680 32088 3732
rect 52736 3680 52788 3732
rect 2964 3612 3016 3664
rect 3608 3612 3660 3664
rect 6276 3612 6328 3664
rect 6736 3612 6788 3664
rect 7472 3655 7524 3664
rect 7472 3621 7481 3655
rect 7481 3621 7515 3655
rect 7515 3621 7524 3655
rect 7472 3612 7524 3621
rect 8484 3612 8536 3664
rect 6184 3587 6236 3596
rect 6184 3553 6193 3587
rect 6193 3553 6227 3587
rect 6227 3553 6236 3587
rect 6184 3544 6236 3553
rect 8024 3587 8076 3596
rect 8024 3553 8033 3587
rect 8033 3553 8067 3587
rect 8067 3553 8076 3587
rect 8024 3544 8076 3553
rect 8760 3544 8812 3596
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 2412 3476 2464 3528
rect 3424 3408 3476 3460
rect 5816 3476 5868 3528
rect 10140 3544 10192 3596
rect 10416 3544 10468 3596
rect 10692 3544 10744 3596
rect 10968 3655 11020 3664
rect 10968 3621 10977 3655
rect 10977 3621 11011 3655
rect 11011 3621 11020 3655
rect 10968 3612 11020 3621
rect 16396 3612 16448 3664
rect 17868 3655 17920 3664
rect 17868 3621 17877 3655
rect 17877 3621 17911 3655
rect 17911 3621 17920 3655
rect 17868 3612 17920 3621
rect 19064 3612 19116 3664
rect 25504 3612 25556 3664
rect 46296 3612 46348 3664
rect 51448 3612 51500 3664
rect 11980 3544 12032 3596
rect 14372 3544 14424 3596
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 15936 3544 15988 3596
rect 9220 3519 9272 3528
rect 9220 3485 9229 3519
rect 9229 3485 9263 3519
rect 9263 3485 9272 3519
rect 9220 3476 9272 3485
rect 9588 3476 9640 3528
rect 10324 3476 10376 3528
rect 10600 3476 10652 3528
rect 11704 3476 11756 3528
rect 5080 3408 5132 3460
rect 3332 3340 3384 3392
rect 3516 3340 3568 3392
rect 8484 3340 8536 3392
rect 8576 3340 8628 3392
rect 9404 3340 9456 3392
rect 13912 3476 13964 3528
rect 14004 3476 14056 3528
rect 14924 3476 14976 3528
rect 15752 3476 15804 3528
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 17408 3544 17460 3596
rect 18696 3544 18748 3596
rect 21456 3544 21508 3596
rect 30932 3587 30984 3596
rect 30932 3553 30941 3587
rect 30941 3553 30975 3587
rect 30975 3553 30984 3587
rect 30932 3544 30984 3553
rect 50804 3544 50856 3596
rect 51632 3544 51684 3596
rect 53840 3544 53892 3596
rect 17500 3476 17552 3528
rect 18328 3476 18380 3528
rect 19524 3476 19576 3528
rect 20812 3476 20864 3528
rect 21640 3476 21692 3528
rect 23664 3476 23716 3528
rect 23940 3476 23992 3528
rect 24768 3476 24820 3528
rect 25596 3476 25648 3528
rect 26700 3476 26752 3528
rect 27528 3476 27580 3528
rect 28632 3476 28684 3528
rect 30840 3476 30892 3528
rect 34704 3476 34756 3528
rect 35348 3476 35400 3528
rect 35808 3476 35860 3528
rect 36636 3476 36688 3528
rect 37464 3476 37516 3528
rect 38568 3476 38620 3528
rect 39948 3476 40000 3528
rect 40500 3476 40552 3528
rect 41052 3476 41104 3528
rect 42432 3476 42484 3528
rect 42708 3476 42760 3528
rect 44364 3476 44416 3528
rect 45192 3476 45244 3528
rect 46020 3476 46072 3528
rect 47676 3476 47728 3528
rect 48228 3476 48280 3528
rect 50160 3476 50212 3528
rect 50620 3476 50672 3528
rect 51172 3476 51224 3528
rect 52276 3476 52328 3528
rect 13544 3408 13596 3460
rect 14832 3408 14884 3460
rect 15292 3408 15344 3460
rect 17776 3408 17828 3460
rect 23480 3408 23532 3460
rect 53288 3408 53340 3460
rect 57520 3519 57572 3528
rect 57520 3485 57529 3519
rect 57529 3485 57563 3519
rect 57563 3485 57572 3519
rect 57520 3476 57572 3485
rect 58164 3519 58216 3528
rect 58164 3485 58173 3519
rect 58173 3485 58207 3519
rect 58207 3485 58216 3519
rect 58164 3476 58216 3485
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 19524 3340 19576 3392
rect 22836 3340 22888 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 3792 3179 3844 3188
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 4712 3136 4764 3188
rect 1952 3111 2004 3120
rect 1952 3077 1961 3111
rect 1961 3077 1995 3111
rect 1995 3077 2004 3111
rect 1952 3068 2004 3077
rect 2780 3068 2832 3120
rect 3240 3068 3292 3120
rect 6828 3136 6880 3188
rect 6920 3136 6972 3188
rect 8024 3136 8076 3188
rect 8576 3136 8628 3188
rect 8852 3136 8904 3188
rect 14464 3179 14516 3188
rect 14464 3145 14473 3179
rect 14473 3145 14507 3179
rect 14507 3145 14516 3179
rect 14464 3136 14516 3145
rect 1492 3000 1544 3052
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 4804 3000 4856 3052
rect 5264 3000 5316 3052
rect 6460 3000 6512 3052
rect 7380 3068 7432 3120
rect 13728 3068 13780 3120
rect 15108 3111 15160 3120
rect 3700 2932 3752 2984
rect 6092 2932 6144 2984
rect 7564 3000 7616 3052
rect 8208 3000 8260 3052
rect 8484 3000 8536 3052
rect 8760 3000 8812 3052
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 15108 3077 15117 3111
rect 15117 3077 15151 3111
rect 15151 3077 15160 3111
rect 15108 3068 15160 3077
rect 16304 3068 16356 3120
rect 16672 3136 16724 3188
rect 17040 3136 17092 3188
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 18880 3179 18932 3188
rect 18880 3145 18889 3179
rect 18889 3145 18923 3179
rect 18923 3145 18932 3179
rect 18880 3136 18932 3145
rect 20352 3179 20404 3188
rect 20352 3145 20361 3179
rect 20361 3145 20395 3179
rect 20395 3145 20404 3179
rect 20352 3136 20404 3145
rect 21088 3179 21140 3188
rect 21088 3145 21097 3179
rect 21097 3145 21131 3179
rect 21131 3145 21140 3179
rect 21088 3136 21140 3145
rect 21272 3136 21324 3188
rect 22652 3136 22704 3188
rect 23020 3179 23072 3188
rect 23020 3145 23029 3179
rect 23029 3145 23063 3179
rect 23063 3145 23072 3179
rect 23020 3136 23072 3145
rect 17316 3068 17368 3120
rect 17592 3111 17644 3120
rect 17592 3077 17601 3111
rect 17601 3077 17635 3111
rect 17635 3077 17644 3111
rect 17592 3068 17644 3077
rect 14832 3000 14884 3052
rect 15016 3000 15068 3052
rect 15568 3000 15620 3052
rect 16580 3000 16632 3052
rect 17776 3000 17828 3052
rect 17960 3000 18012 3052
rect 18604 3000 18656 3052
rect 18880 3000 18932 3052
rect 19064 3043 19116 3052
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 19984 3000 20036 3052
rect 20260 3068 20312 3120
rect 20536 3068 20588 3120
rect 22192 3068 22244 3120
rect 51908 3068 51960 3120
rect 2596 2796 2648 2848
rect 5356 2864 5408 2916
rect 7748 2864 7800 2916
rect 5632 2839 5684 2848
rect 5632 2805 5641 2839
rect 5641 2805 5675 2839
rect 5675 2805 5684 2839
rect 5632 2796 5684 2805
rect 6552 2796 6604 2848
rect 8024 2864 8076 2916
rect 10416 2932 10468 2984
rect 15660 2932 15712 2984
rect 21364 3000 21416 3052
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22836 3043 22888 3052
rect 22100 3000 22152 3009
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 23204 2932 23256 2984
rect 24492 2932 24544 2984
rect 9404 2864 9456 2916
rect 14924 2864 14976 2916
rect 9496 2796 9548 2848
rect 9680 2796 9732 2848
rect 14740 2796 14792 2848
rect 17868 2864 17920 2916
rect 17960 2864 18012 2916
rect 18880 2864 18932 2916
rect 34520 3000 34572 3052
rect 51724 3000 51776 3052
rect 54760 3000 54812 3052
rect 32772 2932 32824 2984
rect 38292 2932 38344 2984
rect 42156 2932 42208 2984
rect 53104 2932 53156 2984
rect 56600 2975 56652 2984
rect 56600 2941 56609 2975
rect 56609 2941 56643 2975
rect 56643 2941 56652 2975
rect 56600 2932 56652 2941
rect 33876 2864 33928 2916
rect 37188 2864 37240 2916
rect 39120 2864 39172 2916
rect 40224 2864 40276 2916
rect 42984 2864 43036 2916
rect 44088 2864 44140 2916
rect 19432 2796 19484 2848
rect 22376 2796 22428 2848
rect 25044 2796 25096 2848
rect 25320 2796 25372 2848
rect 26148 2796 26200 2848
rect 26884 2796 26936 2848
rect 27804 2796 27856 2848
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 29184 2796 29236 2848
rect 29736 2796 29788 2848
rect 30012 2839 30064 2848
rect 30012 2805 30021 2839
rect 30021 2805 30055 2839
rect 30055 2805 30064 2839
rect 30012 2796 30064 2805
rect 30564 2796 30616 2848
rect 31668 2796 31720 2848
rect 32220 2796 32272 2848
rect 33324 2796 33376 2848
rect 34428 2796 34480 2848
rect 35440 2796 35492 2848
rect 36360 2796 36412 2848
rect 37740 2796 37792 2848
rect 39672 2796 39724 2848
rect 41604 2796 41656 2848
rect 43536 2796 43588 2848
rect 44916 2796 44968 2848
rect 47400 2864 47452 2916
rect 48780 2864 48832 2916
rect 49884 2864 49936 2916
rect 50988 2864 51040 2916
rect 54208 2864 54260 2916
rect 45468 2796 45520 2848
rect 46848 2796 46900 2848
rect 47952 2796 48004 2848
rect 49332 2796 49384 2848
rect 50712 2796 50764 2848
rect 51540 2796 51592 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 6276 2592 6328 2644
rect 8576 2592 8628 2644
rect 14740 2592 14792 2644
rect 2688 2524 2740 2576
rect 7380 2524 7432 2576
rect 9680 2524 9732 2576
rect 14556 2524 14608 2576
rect 7656 2456 7708 2508
rect 12624 2456 12676 2508
rect 15844 2592 15896 2644
rect 16120 2592 16172 2644
rect 17132 2635 17184 2644
rect 17132 2601 17141 2635
rect 17141 2601 17175 2635
rect 17175 2601 17184 2635
rect 17132 2592 17184 2601
rect 17684 2592 17736 2644
rect 19616 2592 19668 2644
rect 20444 2592 20496 2644
rect 27344 2592 27396 2644
rect 16304 2524 16356 2576
rect 18512 2567 18564 2576
rect 18512 2533 18521 2567
rect 18521 2533 18555 2567
rect 18555 2533 18564 2567
rect 18512 2524 18564 2533
rect 20352 2524 20404 2576
rect 22652 2524 22704 2576
rect 23572 2567 23624 2576
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 3056 2388 3108 2440
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 4988 2388 5040 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 7104 2388 7156 2440
rect 11520 2431 11572 2440
rect 3700 2320 3752 2372
rect 4252 2295 4304 2304
rect 4252 2261 4261 2295
rect 4261 2261 4295 2295
rect 4295 2261 4304 2295
rect 4252 2252 4304 2261
rect 5816 2252 5868 2304
rect 8668 2320 8720 2372
rect 9036 2363 9088 2372
rect 9036 2329 9045 2363
rect 9045 2329 9079 2363
rect 9079 2329 9088 2363
rect 9036 2320 9088 2329
rect 9220 2320 9272 2372
rect 11520 2397 11529 2431
rect 11529 2397 11563 2431
rect 11563 2397 11572 2431
rect 11520 2388 11572 2397
rect 12716 2388 12768 2440
rect 17224 2456 17276 2508
rect 19984 2456 20036 2508
rect 20168 2456 20220 2508
rect 17960 2431 18012 2440
rect 15476 2320 15528 2372
rect 17960 2397 17969 2431
rect 17969 2397 18003 2431
rect 18003 2397 18012 2431
rect 17960 2388 18012 2397
rect 19524 2388 19576 2440
rect 20996 2456 21048 2508
rect 23572 2533 23581 2567
rect 23581 2533 23615 2567
rect 23615 2533 23624 2567
rect 23572 2524 23624 2533
rect 26424 2524 26476 2576
rect 28356 2524 28408 2576
rect 35624 2592 35676 2644
rect 36728 2524 36780 2576
rect 42892 2592 42944 2644
rect 52000 2592 52052 2644
rect 31944 2456 31996 2508
rect 33048 2456 33100 2508
rect 35624 2456 35676 2508
rect 38016 2524 38068 2576
rect 41880 2524 41932 2576
rect 45744 2524 45796 2576
rect 49608 2524 49660 2576
rect 36912 2456 36964 2508
rect 38844 2456 38896 2508
rect 40776 2456 40828 2508
rect 43260 2456 43312 2508
rect 46572 2456 46624 2508
rect 48504 2456 48556 2508
rect 51264 2456 51316 2508
rect 54392 2524 54444 2576
rect 52552 2456 52604 2508
rect 53564 2456 53616 2508
rect 20720 2388 20772 2440
rect 21272 2431 21324 2440
rect 21272 2397 21281 2431
rect 21281 2397 21315 2431
rect 21315 2397 21324 2431
rect 21272 2388 21324 2397
rect 22468 2388 22520 2440
rect 18052 2320 18104 2372
rect 20260 2320 20312 2372
rect 8024 2252 8076 2304
rect 10048 2252 10100 2304
rect 10416 2295 10468 2304
rect 10416 2261 10425 2295
rect 10425 2261 10459 2295
rect 10459 2261 10468 2295
rect 10416 2252 10468 2261
rect 16028 2295 16080 2304
rect 16028 2261 16037 2295
rect 16037 2261 16071 2295
rect 16071 2261 16080 2295
rect 16028 2252 16080 2261
rect 20352 2295 20404 2304
rect 20352 2261 20361 2295
rect 20361 2261 20395 2295
rect 20395 2261 20404 2295
rect 20352 2252 20404 2261
rect 23296 2388 23348 2440
rect 25872 2388 25924 2440
rect 27252 2388 27304 2440
rect 27344 2388 27396 2440
rect 23572 2320 23624 2372
rect 28908 2388 28960 2440
rect 29460 2388 29512 2440
rect 30288 2388 30340 2440
rect 30840 2388 30892 2440
rect 31116 2388 31168 2440
rect 31392 2388 31444 2440
rect 32496 2388 32548 2440
rect 33600 2388 33652 2440
rect 35716 2388 35768 2440
rect 36084 2388 36136 2440
rect 39396 2388 39448 2440
rect 41328 2388 41380 2440
rect 43812 2388 43864 2440
rect 23020 2252 23072 2304
rect 36544 2320 36596 2372
rect 36728 2320 36780 2372
rect 43168 2320 43220 2372
rect 44640 2320 44692 2372
rect 47124 2388 47176 2440
rect 49056 2388 49108 2440
rect 50896 2388 50948 2440
rect 52368 2320 52420 2372
rect 56324 2252 56376 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 5816 2048 5868 2100
rect 8300 2048 8352 2100
rect 4068 1980 4120 2032
rect 7656 1980 7708 2032
rect 6828 1912 6880 1964
rect 7104 1912 7156 1964
rect 4252 1844 4304 1896
rect 18788 2048 18840 2100
rect 22652 2048 22704 2100
rect 35624 2048 35676 2100
rect 36544 2048 36596 2100
rect 44732 2048 44784 2100
rect 52736 2048 52788 2100
rect 52920 2048 52972 2100
rect 54392 2048 54444 2100
rect 10048 1980 10100 2032
rect 12900 1980 12952 2032
rect 20352 1980 20404 2032
rect 43444 1980 43496 2032
rect 10416 1844 10468 1896
rect 29552 1844 29604 1896
rect 5908 1776 5960 1828
rect 6644 1776 6696 1828
rect 15476 1708 15528 1760
rect 16396 1708 16448 1760
rect 20720 1708 20772 1760
rect 21088 1708 21140 1760
rect 21272 1708 21324 1760
rect 21916 1708 21968 1760
rect 5356 1572 5408 1624
rect 5908 1572 5960 1624
rect 14004 1436 14056 1488
rect 15016 1436 15068 1488
rect 19340 1436 19392 1488
rect 19800 1436 19852 1488
rect 4620 1368 4672 1420
rect 5724 1368 5776 1420
rect 14280 1368 14332 1420
rect 14740 1368 14792 1420
rect 19708 1368 19760 1420
rect 20168 1368 20220 1420
rect 34152 1368 34204 1420
rect 35716 1368 35768 1420
rect 4804 1300 4856 1352
rect 6184 1300 6236 1352
rect 19432 1300 19484 1352
rect 19616 1300 19668 1352
rect 52828 1436 52880 1488
rect 53012 1436 53064 1488
rect 53012 1300 53064 1352
rect 52552 1096 52604 1148
rect 52552 960 52604 1012
rect 54760 960 54812 1012
rect 50988 892 51040 944
<< metal2 >>
rect 1766 59200 1822 60000
rect 3330 59200 3386 60000
rect 4894 59200 4950 60000
rect 6458 59200 6514 60000
rect 8022 59200 8078 60000
rect 9586 59200 9642 60000
rect 11150 59200 11206 60000
rect 12714 59200 12770 60000
rect 14278 59200 14334 60000
rect 15842 59200 15898 60000
rect 17406 59200 17462 60000
rect 18970 59200 19026 60000
rect 19076 59214 19288 59242
rect 1780 57458 1808 59200
rect 3344 57458 3372 59200
rect 4908 57458 4936 59200
rect 6472 57458 6500 59200
rect 8036 57458 8064 59200
rect 1768 57452 1820 57458
rect 1768 57394 1820 57400
rect 3332 57452 3384 57458
rect 3332 57394 3384 57400
rect 4896 57452 4948 57458
rect 4896 57394 4948 57400
rect 6460 57452 6512 57458
rect 6460 57394 6512 57400
rect 8024 57452 8076 57458
rect 9600 57440 9628 59200
rect 11164 57458 11192 59200
rect 12728 57594 12756 59200
rect 14292 57594 14320 59200
rect 15856 57594 15884 59200
rect 17420 57594 17448 59200
rect 18984 59106 19012 59200
rect 19076 59106 19104 59214
rect 18984 59078 19104 59106
rect 19260 57610 19288 59214
rect 20534 59200 20590 60000
rect 22098 59200 22154 60000
rect 23662 59200 23718 60000
rect 25226 59200 25282 60000
rect 26790 59200 26846 60000
rect 28354 59200 28410 60000
rect 29918 59200 29974 60000
rect 31482 59200 31538 60000
rect 33046 59200 33102 60000
rect 34610 59200 34666 60000
rect 36174 59200 36230 60000
rect 37738 59200 37794 60000
rect 39302 59200 39358 60000
rect 40866 59200 40922 60000
rect 42430 59200 42486 60000
rect 43994 59200 44050 60000
rect 45558 59200 45614 60000
rect 47122 59200 47178 60000
rect 48686 59200 48742 60000
rect 50250 59200 50306 60000
rect 51814 59200 51870 60000
rect 53378 59200 53434 60000
rect 54942 59200 54998 60000
rect 56506 59200 56562 60000
rect 58070 59200 58126 60000
rect 58438 59256 58494 59265
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 20548 57610 20576 59200
rect 19260 57594 19380 57610
rect 20548 57594 20760 57610
rect 22112 57594 22140 59200
rect 23676 57594 23704 59200
rect 25240 57594 25268 59200
rect 26804 57594 26832 59200
rect 28368 57594 28396 59200
rect 29932 57594 29960 59200
rect 31496 57594 31524 59200
rect 12716 57588 12768 57594
rect 12716 57530 12768 57536
rect 14280 57588 14332 57594
rect 14280 57530 14332 57536
rect 15844 57588 15896 57594
rect 15844 57530 15896 57536
rect 17408 57588 17460 57594
rect 19260 57588 19392 57594
rect 19260 57582 19340 57588
rect 17408 57530 17460 57536
rect 20548 57588 20772 57594
rect 20548 57582 20720 57588
rect 19340 57530 19392 57536
rect 20720 57530 20772 57536
rect 22100 57588 22152 57594
rect 22100 57530 22152 57536
rect 23664 57588 23716 57594
rect 23664 57530 23716 57536
rect 25228 57588 25280 57594
rect 25228 57530 25280 57536
rect 26792 57588 26844 57594
rect 26792 57530 26844 57536
rect 28356 57588 28408 57594
rect 28356 57530 28408 57536
rect 29920 57588 29972 57594
rect 29920 57530 29972 57536
rect 31484 57588 31536 57594
rect 33060 57576 33088 59200
rect 34624 57594 34652 59200
rect 36188 57594 36216 59200
rect 37752 57594 37780 59200
rect 39316 57594 39344 59200
rect 40880 57594 40908 59200
rect 42444 57594 42472 59200
rect 33140 57588 33192 57594
rect 33060 57548 33140 57576
rect 31484 57530 31536 57536
rect 33140 57530 33192 57536
rect 34612 57588 34664 57594
rect 34612 57530 34664 57536
rect 36176 57588 36228 57594
rect 36176 57530 36228 57536
rect 37740 57588 37792 57594
rect 37740 57530 37792 57536
rect 39304 57588 39356 57594
rect 39304 57530 39356 57536
rect 40868 57588 40920 57594
rect 40868 57530 40920 57536
rect 42432 57588 42484 57594
rect 44008 57576 44036 59200
rect 45572 57594 45600 59200
rect 47136 57594 47164 59200
rect 48700 57594 48728 59200
rect 50264 57882 50292 59200
rect 50172 57854 50292 57882
rect 50172 57594 50200 57854
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 51828 57594 51856 59200
rect 53392 57594 53420 59200
rect 54956 57594 54984 59200
rect 56520 57610 56548 59200
rect 57518 57896 57574 57905
rect 57518 57831 57574 57840
rect 56520 57594 56640 57610
rect 44180 57588 44232 57594
rect 44008 57548 44180 57576
rect 42432 57530 42484 57536
rect 44180 57530 44232 57536
rect 45560 57588 45612 57594
rect 45560 57530 45612 57536
rect 47124 57588 47176 57594
rect 47124 57530 47176 57536
rect 48688 57588 48740 57594
rect 48688 57530 48740 57536
rect 50160 57588 50212 57594
rect 50160 57530 50212 57536
rect 51816 57588 51868 57594
rect 51816 57530 51868 57536
rect 53380 57588 53432 57594
rect 53380 57530 53432 57536
rect 54944 57588 54996 57594
rect 56520 57588 56652 57594
rect 56520 57582 56600 57588
rect 54944 57530 54996 57536
rect 56600 57530 56652 57536
rect 20904 57520 20956 57526
rect 20904 57462 20956 57468
rect 31760 57520 31812 57526
rect 31760 57462 31812 57468
rect 46204 57520 46256 57526
rect 46204 57462 46256 57468
rect 9680 57452 9732 57458
rect 9600 57412 9680 57440
rect 8024 57394 8076 57400
rect 9680 57394 9732 57400
rect 11152 57452 11204 57458
rect 11152 57394 11204 57400
rect 13084 57452 13136 57458
rect 13084 57394 13136 57400
rect 14648 57452 14700 57458
rect 14648 57394 14700 57400
rect 16672 57452 16724 57458
rect 16672 57394 16724 57400
rect 17500 57452 17552 57458
rect 17500 57394 17552 57400
rect 19248 57452 19300 57458
rect 19248 57394 19300 57400
rect 20628 57452 20680 57458
rect 20628 57394 20680 57400
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 13096 56506 13124 57394
rect 14660 56506 14688 57394
rect 16488 56704 16540 56710
rect 16488 56646 16540 56652
rect 13084 56500 13136 56506
rect 13084 56442 13136 56448
rect 14648 56500 14700 56506
rect 14648 56442 14700 56448
rect 16500 56370 16528 56646
rect 16684 56506 16712 57394
rect 17512 56506 17540 57394
rect 16672 56500 16724 56506
rect 16672 56442 16724 56448
rect 17500 56500 17552 56506
rect 17500 56442 17552 56448
rect 14188 56364 14240 56370
rect 14188 56306 14240 56312
rect 15108 56364 15160 56370
rect 15108 56306 15160 56312
rect 16488 56364 16540 56370
rect 16488 56306 16540 56312
rect 16580 56364 16632 56370
rect 16580 56306 16632 56312
rect 17224 56364 17276 56370
rect 17224 56306 17276 56312
rect 17868 56364 17920 56370
rect 17868 56306 17920 56312
rect 18604 56364 18656 56370
rect 18604 56306 18656 56312
rect 19064 56364 19116 56370
rect 19064 56306 19116 56312
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 14200 55622 14228 56306
rect 15120 55622 15148 56306
rect 16396 55684 16448 55690
rect 16396 55626 16448 55632
rect 14188 55616 14240 55622
rect 14186 55584 14188 55593
rect 15108 55616 15160 55622
rect 14240 55584 14242 55593
rect 15108 55558 15160 55564
rect 14186 55519 14242 55528
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 12532 42220 12584 42226
rect 12532 42162 12584 42168
rect 15016 42220 15068 42226
rect 15016 42162 15068 42168
rect 12440 42084 12492 42090
rect 12440 42026 12492 42032
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 11520 41744 11572 41750
rect 11518 41712 11520 41721
rect 11572 41712 11574 41721
rect 11518 41647 11574 41656
rect 11704 41540 11756 41546
rect 11704 41482 11756 41488
rect 9680 41472 9732 41478
rect 9680 41414 9732 41420
rect 9404 41132 9456 41138
rect 9404 41074 9456 41080
rect 8944 40928 8996 40934
rect 8944 40870 8996 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4896 40656 4948 40662
rect 4896 40598 4948 40604
rect 4252 40520 4304 40526
rect 4252 40462 4304 40468
rect 4804 40520 4856 40526
rect 4804 40462 4856 40468
rect 3792 40384 3844 40390
rect 3792 40326 3844 40332
rect 3804 40118 3832 40326
rect 4264 40186 4292 40462
rect 4252 40180 4304 40186
rect 4252 40122 4304 40128
rect 3792 40112 3844 40118
rect 3792 40054 3844 40060
rect 4816 40050 4844 40462
rect 4908 40458 4936 40598
rect 6092 40520 6144 40526
rect 6092 40462 6144 40468
rect 4896 40452 4948 40458
rect 4896 40394 4948 40400
rect 5816 40452 5868 40458
rect 5816 40394 5868 40400
rect 4712 40044 4764 40050
rect 4712 39986 4764 39992
rect 4804 40044 4856 40050
rect 4804 39986 4856 39992
rect 1860 39976 1912 39982
rect 1860 39918 1912 39924
rect 1872 39438 1900 39918
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 1860 39432 1912 39438
rect 1860 39374 1912 39380
rect 1872 38350 1900 39374
rect 4724 39001 4752 39986
rect 4710 38992 4766 39001
rect 3053 38956 3105 38962
rect 3053 38898 3105 38904
rect 3148 38956 3200 38962
rect 3148 38898 3200 38904
rect 3332 38956 3384 38962
rect 4710 38927 4766 38936
rect 3332 38898 3384 38904
rect 2872 38820 2924 38826
rect 2872 38762 2924 38768
rect 2688 38752 2740 38758
rect 2688 38694 2740 38700
rect 2700 38350 2728 38694
rect 1860 38344 1912 38350
rect 1860 38286 1912 38292
rect 2688 38344 2740 38350
rect 2688 38286 2740 38292
rect 1872 37330 1900 38286
rect 2780 37868 2832 37874
rect 2780 37810 2832 37816
rect 2688 37664 2740 37670
rect 2688 37606 2740 37612
rect 1860 37324 1912 37330
rect 1860 37266 1912 37272
rect 1872 36242 1900 37266
rect 2700 37262 2728 37606
rect 2792 37466 2820 37810
rect 2780 37460 2832 37466
rect 2780 37402 2832 37408
rect 2688 37256 2740 37262
rect 2688 37198 2740 37204
rect 1860 36236 1912 36242
rect 1860 36178 1912 36184
rect 2688 35148 2740 35154
rect 2688 35090 2740 35096
rect 2412 34536 2464 34542
rect 2412 34478 2464 34484
rect 2424 33454 2452 34478
rect 2412 33448 2464 33454
rect 2412 33390 2464 33396
rect 2424 31822 2452 33390
rect 2412 31816 2464 31822
rect 2412 31758 2464 31764
rect 2136 31748 2188 31754
rect 2136 31690 2188 31696
rect 2148 31482 2176 31690
rect 2136 31476 2188 31482
rect 2136 31418 2188 31424
rect 2424 30802 2452 31758
rect 2700 31414 2728 35090
rect 2780 34604 2832 34610
rect 2780 34546 2832 34552
rect 2792 34202 2820 34546
rect 2780 34196 2832 34202
rect 2780 34138 2832 34144
rect 2884 33998 2912 38762
rect 3068 38010 3096 38898
rect 3160 38010 3188 38898
rect 3344 38758 3372 38898
rect 3332 38752 3384 38758
rect 3332 38694 3384 38700
rect 3056 38004 3108 38010
rect 3056 37946 3108 37952
rect 3148 38004 3200 38010
rect 3148 37946 3200 37952
rect 3344 37874 3372 38694
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4724 37942 4752 38927
rect 4816 38758 4844 39986
rect 4804 38752 4856 38758
rect 4804 38694 4856 38700
rect 4712 37936 4764 37942
rect 4712 37878 4764 37884
rect 3332 37868 3384 37874
rect 3332 37810 3384 37816
rect 3424 37868 3476 37874
rect 3424 37810 3476 37816
rect 3436 37754 3464 37810
rect 3344 37726 3464 37754
rect 3344 37126 3372 37726
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4068 37460 4120 37466
rect 4068 37402 4120 37408
rect 3332 37120 3384 37126
rect 3332 37062 3384 37068
rect 2964 34944 3016 34950
rect 2964 34886 3016 34892
rect 2872 33992 2924 33998
rect 2872 33934 2924 33940
rect 2688 31408 2740 31414
rect 2688 31350 2740 31356
rect 2412 30796 2464 30802
rect 2412 30738 2464 30744
rect 2424 30258 2452 30738
rect 2412 30252 2464 30258
rect 2412 30194 2464 30200
rect 2504 30252 2556 30258
rect 2504 30194 2556 30200
rect 2516 29850 2544 30194
rect 2504 29844 2556 29850
rect 2504 29786 2556 29792
rect 2596 29640 2648 29646
rect 2700 29628 2728 31350
rect 2872 31340 2924 31346
rect 2976 31328 3004 34886
rect 3148 34400 3200 34406
rect 3148 34342 3200 34348
rect 3160 33998 3188 34342
rect 3148 33992 3200 33998
rect 3148 33934 3200 33940
rect 3240 33856 3292 33862
rect 3240 33798 3292 33804
rect 2924 31300 3004 31328
rect 2872 31282 2924 31288
rect 2780 31204 2832 31210
rect 2780 31146 2832 31152
rect 2792 30598 2820 31146
rect 2780 30592 2832 30598
rect 2780 30534 2832 30540
rect 2648 29600 2728 29628
rect 2596 29582 2648 29588
rect 2608 29238 2636 29582
rect 2688 29504 2740 29510
rect 2688 29446 2740 29452
rect 2596 29232 2648 29238
rect 2596 29174 2648 29180
rect 2700 28762 2728 29446
rect 2688 28756 2740 28762
rect 2688 28698 2740 28704
rect 2596 28008 2648 28014
rect 2596 27950 2648 27956
rect 2608 25906 2636 27950
rect 2792 27130 2820 30534
rect 2884 29646 2912 31282
rect 2964 29776 3016 29782
rect 2964 29718 3016 29724
rect 2872 29640 2924 29646
rect 2872 29582 2924 29588
rect 2884 29306 2912 29582
rect 2872 29300 2924 29306
rect 2872 29242 2924 29248
rect 2872 28960 2924 28966
rect 2872 28902 2924 28908
rect 2884 28082 2912 28902
rect 2872 28076 2924 28082
rect 2872 28018 2924 28024
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 2792 26382 2820 27066
rect 2780 26376 2832 26382
rect 2780 26318 2832 26324
rect 2596 25900 2648 25906
rect 2596 25842 2648 25848
rect 2608 25294 2636 25842
rect 2596 25288 2648 25294
rect 2596 25230 2648 25236
rect 2608 24818 2636 25230
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 2240 23050 2268 23666
rect 2504 23520 2556 23526
rect 2504 23462 2556 23468
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2240 22710 2268 22986
rect 2228 22704 2280 22710
rect 2228 22646 2280 22652
rect 2516 22094 2544 23462
rect 2608 22710 2636 24754
rect 2792 24698 2820 26318
rect 2872 26240 2924 26246
rect 2872 26182 2924 26188
rect 2884 25974 2912 26182
rect 2872 25968 2924 25974
rect 2872 25910 2924 25916
rect 2872 25288 2924 25294
rect 2976 25276 3004 29718
rect 3252 29322 3280 33798
rect 3344 29714 3372 37062
rect 3608 35692 3660 35698
rect 3608 35634 3660 35640
rect 3424 31680 3476 31686
rect 3424 31622 3476 31628
rect 3436 31346 3464 31622
rect 3620 31346 3648 35634
rect 4080 34202 4108 37402
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4712 36100 4764 36106
rect 4712 36042 4764 36048
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4724 35290 4752 36042
rect 4712 35284 4764 35290
rect 4712 35226 4764 35232
rect 4712 34604 4764 34610
rect 4712 34546 4764 34552
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 34196 4120 34202
rect 4068 34138 4120 34144
rect 4080 33998 4108 34138
rect 4068 33992 4120 33998
rect 4068 33934 4120 33940
rect 4344 33992 4396 33998
rect 4344 33934 4396 33940
rect 3792 33856 3844 33862
rect 3792 33798 3844 33804
rect 3804 33590 3832 33798
rect 4356 33658 4384 33934
rect 4344 33652 4396 33658
rect 4344 33594 4396 33600
rect 3792 33584 3844 33590
rect 3792 33526 3844 33532
rect 4724 33522 4752 34546
rect 4620 33516 4672 33522
rect 4620 33458 4672 33464
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3424 31340 3476 31346
rect 3424 31282 3476 31288
rect 3608 31340 3660 31346
rect 3608 31282 3660 31288
rect 3332 29708 3384 29714
rect 3332 29650 3384 29656
rect 3436 29646 3464 31282
rect 3424 29640 3476 29646
rect 3424 29582 3476 29588
rect 3252 29294 3372 29322
rect 3240 26852 3292 26858
rect 3240 26794 3292 26800
rect 3056 26784 3108 26790
rect 3056 26726 3108 26732
rect 3068 26382 3096 26726
rect 3148 26444 3200 26450
rect 3148 26386 3200 26392
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 3056 26240 3108 26246
rect 3056 26182 3108 26188
rect 3068 25294 3096 26182
rect 3160 25362 3188 26386
rect 3252 26382 3280 26794
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3148 25356 3200 25362
rect 3148 25298 3200 25304
rect 3252 25294 3280 26318
rect 2924 25248 3004 25276
rect 2872 25230 2924 25236
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2884 24886 2912 25094
rect 2872 24880 2924 24886
rect 2872 24822 2924 24828
rect 2792 24670 2912 24698
rect 2688 23112 2740 23118
rect 2686 23080 2688 23089
rect 2780 23112 2832 23118
rect 2740 23080 2742 23089
rect 2780 23054 2832 23060
rect 2686 23015 2742 23024
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2596 22704 2648 22710
rect 2596 22646 2648 22652
rect 2700 22642 2728 22918
rect 2792 22778 2820 23054
rect 2780 22772 2832 22778
rect 2780 22714 2832 22720
rect 2688 22636 2740 22642
rect 2688 22578 2740 22584
rect 2884 22094 2912 24670
rect 2976 23322 3004 25248
rect 3056 25288 3108 25294
rect 3056 25230 3108 25236
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3252 24410 3280 25230
rect 3344 24818 3372 29294
rect 3620 28490 3648 31282
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3700 30048 3752 30054
rect 3700 29990 3752 29996
rect 3712 29170 3740 29990
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 3700 29164 3752 29170
rect 3700 29106 3752 29112
rect 3712 28558 3740 29106
rect 3792 29096 3844 29102
rect 3792 29038 3844 29044
rect 3804 28762 3832 29038
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 3792 28756 3844 28762
rect 3792 28698 3844 28704
rect 3700 28552 3752 28558
rect 3700 28494 3752 28500
rect 3976 28552 4028 28558
rect 3976 28494 4028 28500
rect 3608 28484 3660 28490
rect 3608 28426 3660 28432
rect 3988 28218 4016 28494
rect 3976 28212 4028 28218
rect 3976 28154 4028 28160
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27396 4120 27402
rect 4068 27338 4120 27344
rect 3976 27056 4028 27062
rect 3976 26998 4028 27004
rect 3988 26042 4016 26998
rect 4080 26382 4108 27338
rect 4632 27130 4660 33458
rect 4908 32570 4936 40394
rect 5448 40384 5500 40390
rect 5448 40326 5500 40332
rect 5724 40384 5776 40390
rect 5724 40326 5776 40332
rect 4988 40112 5040 40118
rect 4988 40054 5040 40060
rect 4896 32564 4948 32570
rect 4896 32506 4948 32512
rect 4712 29504 4764 29510
rect 4712 29446 4764 29452
rect 4804 29504 4856 29510
rect 4804 29446 4856 29452
rect 4724 29170 4752 29446
rect 4712 29164 4764 29170
rect 4712 29106 4764 29112
rect 4724 28422 4752 29106
rect 4712 28416 4764 28422
rect 4712 28358 4764 28364
rect 4620 27124 4672 27130
rect 4620 27066 4672 27072
rect 4816 26994 4844 29446
rect 4896 29028 4948 29034
rect 4896 28970 4948 28976
rect 4908 27470 4936 28970
rect 5000 28558 5028 40054
rect 5460 40050 5488 40326
rect 5736 40050 5764 40326
rect 5828 40186 5856 40394
rect 5816 40180 5868 40186
rect 5816 40122 5868 40128
rect 5448 40044 5500 40050
rect 5448 39986 5500 39992
rect 5724 40044 5776 40050
rect 5724 39986 5776 39992
rect 5172 39364 5224 39370
rect 5172 39306 5224 39312
rect 5184 39098 5212 39306
rect 5172 39092 5224 39098
rect 5172 39034 5224 39040
rect 5264 39092 5316 39098
rect 5264 39034 5316 39040
rect 5276 38826 5304 39034
rect 5460 38826 5488 39986
rect 6104 39982 6132 40462
rect 7196 40452 7248 40458
rect 7196 40394 7248 40400
rect 6920 40384 6972 40390
rect 6920 40326 6972 40332
rect 6932 40118 6960 40326
rect 6920 40112 6972 40118
rect 6920 40054 6972 40060
rect 6736 40044 6788 40050
rect 6736 39986 6788 39992
rect 6092 39976 6144 39982
rect 6092 39918 6144 39924
rect 5816 39500 5868 39506
rect 5816 39442 5868 39448
rect 5828 38962 5856 39442
rect 6104 39438 6132 39918
rect 6092 39432 6144 39438
rect 6092 39374 6144 39380
rect 6104 39030 6132 39374
rect 6644 39296 6696 39302
rect 6644 39238 6696 39244
rect 6000 39024 6052 39030
rect 6000 38966 6052 38972
rect 6092 39024 6144 39030
rect 6092 38966 6144 38972
rect 5816 38956 5868 38962
rect 5816 38898 5868 38904
rect 5264 38820 5316 38826
rect 5264 38762 5316 38768
rect 5448 38820 5500 38826
rect 5448 38762 5500 38768
rect 5828 38758 5856 38898
rect 5816 38752 5868 38758
rect 5816 38694 5868 38700
rect 5080 38208 5132 38214
rect 5080 38150 5132 38156
rect 5092 37874 5120 38150
rect 5080 37868 5132 37874
rect 5080 37810 5132 37816
rect 5092 29238 5120 37810
rect 5172 36780 5224 36786
rect 5172 36722 5224 36728
rect 5184 36378 5212 36722
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 5184 35766 5212 36314
rect 5172 35760 5224 35766
rect 5172 35702 5224 35708
rect 5172 35488 5224 35494
rect 5172 35430 5224 35436
rect 5184 35086 5212 35430
rect 5172 35080 5224 35086
rect 5172 35022 5224 35028
rect 5264 35012 5316 35018
rect 5316 34972 5580 35000
rect 5264 34954 5316 34960
rect 5448 34672 5500 34678
rect 5448 34614 5500 34620
rect 5172 33992 5224 33998
rect 5172 33934 5224 33940
rect 5184 33862 5212 33934
rect 5264 33924 5316 33930
rect 5264 33866 5316 33872
rect 5172 33856 5224 33862
rect 5172 33798 5224 33804
rect 5184 33590 5212 33798
rect 5172 33584 5224 33590
rect 5172 33526 5224 33532
rect 5184 33114 5212 33526
rect 5276 33114 5304 33866
rect 5172 33108 5224 33114
rect 5172 33050 5224 33056
rect 5264 33108 5316 33114
rect 5264 33050 5316 33056
rect 5276 31958 5304 33050
rect 5356 32564 5408 32570
rect 5356 32506 5408 32512
rect 5264 31952 5316 31958
rect 5264 31894 5316 31900
rect 5368 31822 5396 32506
rect 5172 31816 5224 31822
rect 5172 31758 5224 31764
rect 5356 31816 5408 31822
rect 5356 31758 5408 31764
rect 5184 31482 5212 31758
rect 5172 31476 5224 31482
rect 5172 31418 5224 31424
rect 5172 29640 5224 29646
rect 5172 29582 5224 29588
rect 5080 29232 5132 29238
rect 5080 29174 5132 29180
rect 5184 29170 5212 29582
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 5184 28558 5212 29106
rect 4988 28552 5040 28558
rect 4988 28494 5040 28500
rect 5172 28552 5224 28558
rect 5172 28494 5224 28500
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 5080 27396 5132 27402
rect 5080 27338 5132 27344
rect 5092 27062 5120 27338
rect 5080 27056 5132 27062
rect 5080 26998 5132 27004
rect 4804 26988 4856 26994
rect 5368 26976 5396 31758
rect 5460 27606 5488 34614
rect 5552 34542 5580 34972
rect 5540 34536 5592 34542
rect 5540 34478 5592 34484
rect 5724 34536 5776 34542
rect 5724 34478 5776 34484
rect 5540 34196 5592 34202
rect 5540 34138 5592 34144
rect 5552 33998 5580 34138
rect 5540 33992 5592 33998
rect 5538 33960 5540 33969
rect 5592 33960 5594 33969
rect 5538 33895 5594 33904
rect 5632 31680 5684 31686
rect 5632 31622 5684 31628
rect 5644 30734 5672 31622
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5448 27600 5500 27606
rect 5448 27542 5500 27548
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 4804 26930 4856 26936
rect 5276 26948 5396 26976
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4068 26376 4120 26382
rect 4068 26318 4120 26324
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3332 24812 3384 24818
rect 3332 24754 3384 24760
rect 4080 24682 4108 26318
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 5276 23866 5304 26948
rect 5460 26926 5488 26998
rect 5552 26994 5580 27406
rect 5540 26988 5592 26994
rect 5540 26930 5592 26936
rect 5448 26920 5500 26926
rect 5368 26868 5448 26874
rect 5368 26862 5500 26868
rect 5368 26846 5488 26862
rect 5368 26314 5396 26846
rect 5448 26784 5500 26790
rect 5448 26726 5500 26732
rect 5356 26308 5408 26314
rect 5356 26250 5408 26256
rect 5368 25974 5396 26250
rect 5356 25968 5408 25974
rect 5356 25910 5408 25916
rect 5460 24410 5488 26726
rect 5736 26586 5764 34478
rect 5814 33960 5870 33969
rect 5814 33895 5870 33904
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5736 26314 5764 26522
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5448 24404 5500 24410
rect 5448 24346 5500 24352
rect 5264 23860 5316 23866
rect 5264 23802 5316 23808
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 2964 23316 3016 23322
rect 2964 23258 3016 23264
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 3054 23080 3110 23089
rect 2516 22066 2636 22094
rect 2136 21956 2188 21962
rect 2136 21898 2188 21904
rect 2148 21690 2176 21898
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2608 21554 2636 22066
rect 2792 22066 2912 22094
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2596 21548 2648 21554
rect 2596 21490 2648 21496
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2240 19378 2268 19654
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 1964 17134 1992 19314
rect 2516 18970 2544 19790
rect 2700 19446 2728 21966
rect 2792 21418 2820 22066
rect 2976 21486 3004 23054
rect 3054 23015 3110 23024
rect 3068 21622 3096 23015
rect 3252 22234 3280 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 3792 22772 3844 22778
rect 3792 22714 3844 22720
rect 3804 22438 3832 22714
rect 3792 22432 3844 22438
rect 3792 22374 3844 22380
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3608 21956 3660 21962
rect 3608 21898 3660 21904
rect 3620 21690 3648 21898
rect 3608 21684 3660 21690
rect 3608 21626 3660 21632
rect 3056 21616 3108 21622
rect 3056 21558 3108 21564
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 2964 21480 3016 21486
rect 2964 21422 3016 21428
rect 2780 21412 2832 21418
rect 2780 21354 2832 21360
rect 2792 20874 2820 21354
rect 2780 20868 2832 20874
rect 2780 20810 2832 20816
rect 3896 20806 3924 21490
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 2688 19440 2740 19446
rect 2688 19382 2740 19388
rect 3988 18970 4016 23258
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4632 22642 4660 22986
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4712 22568 4764 22574
rect 4712 22510 4764 22516
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 21622 4660 22374
rect 4724 21894 4752 22510
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 5184 21554 5212 21966
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 5172 21548 5224 21554
rect 5172 21490 5224 21496
rect 5276 21418 5304 21830
rect 5736 21554 5764 26250
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5264 21412 5316 21418
rect 5264 21354 5316 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 5736 21146 5764 21490
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4632 19922 4660 20810
rect 5632 20800 5684 20806
rect 5632 20742 5684 20748
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 4620 19508 4672 19514
rect 4620 19450 4672 19456
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2792 18358 2820 18702
rect 4632 18698 4660 19450
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4620 18692 4672 18698
rect 4672 18652 4752 18680
rect 4620 18634 4672 18640
rect 2780 18352 2832 18358
rect 2780 18294 2832 18300
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1964 16046 1992 17070
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2240 16182 2268 16390
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 1952 16040 2004 16046
rect 1952 15982 2004 15988
rect 1964 15026 1992 15982
rect 2516 15706 2544 16526
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2792 15570 2820 18294
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4620 18284 4672 18290
rect 4620 18226 4672 18232
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2976 17270 3004 18022
rect 4080 17542 4108 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 3884 17060 3936 17066
rect 3884 17002 3936 17008
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 2780 15564 2832 15570
rect 2780 15506 2832 15512
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2792 14618 2820 15506
rect 3804 15502 3832 15846
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3712 14618 3740 14962
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 1584 14544 1636 14550
rect 1584 14486 1636 14492
rect 1400 9920 1452 9926
rect 1400 9862 1452 9868
rect 1412 9586 1440 9862
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 3058 1532 8298
rect 1596 8090 1624 14486
rect 2792 13938 2820 14554
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13394 2820 13874
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 2056 12850 2084 13126
rect 2332 12986 2360 13262
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 3804 12306 3832 12854
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2608 11694 2636 12174
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2884 11762 2912 12038
rect 3068 11898 3096 12106
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 10062 2636 11630
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1596 7993 1624 8026
rect 1582 7984 1638 7993
rect 1582 7919 1638 7928
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5642 1716 6054
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1780 4146 1808 7142
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1768 4140 1820 4146
rect 1768 4082 1820 4088
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 1596 2281 1624 3878
rect 1872 3534 1900 5646
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1964 3126 1992 8570
rect 2056 8498 2084 9454
rect 2332 9178 2360 9998
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2044 8356 2096 8362
rect 2044 8298 2096 8304
rect 1952 3120 2004 3126
rect 1952 3062 2004 3068
rect 2056 2938 2084 8298
rect 2516 7954 2544 8434
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2516 7002 2544 7890
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 2148 6322 2176 6598
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2240 5302 2268 6054
rect 2332 5370 2360 6734
rect 2516 5710 2544 6938
rect 2608 6866 2636 9998
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2780 8832 2832 8838
rect 2778 8800 2780 8809
rect 2832 8800 2834 8809
rect 2778 8735 2834 8744
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2700 6914 2728 7686
rect 2700 6886 2820 6914
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3505 2176 3878
rect 2412 3528 2464 3534
rect 2134 3496 2190 3505
rect 2412 3470 2464 3476
rect 2134 3431 2190 3440
rect 2424 3058 2452 3470
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2226 2952 2282 2961
rect 2056 2910 2226 2938
rect 2226 2887 2282 2896
rect 2240 2446 2268 2887
rect 2608 2854 2636 4082
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2700 2582 2728 6054
rect 2792 5273 2820 6886
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2884 5370 2912 5714
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2778 5264 2834 5273
rect 2778 5199 2780 5208
rect 2832 5199 2834 5208
rect 2780 5170 2832 5176
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 3126 2820 4422
rect 2976 3670 3004 9114
rect 3436 8906 3464 9318
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3436 8566 3464 8842
rect 3424 8560 3476 8566
rect 3424 8502 3476 8508
rect 3056 7812 3108 7818
rect 3056 7754 3108 7760
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2962 2680 3018 2689
rect 2962 2615 3018 2624
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2976 2446 3004 2615
rect 3068 2446 3096 7754
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 4049 3188 7142
rect 3240 6996 3292 7002
rect 3240 6938 3292 6944
rect 3252 6390 3280 6938
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3344 6390 3372 6598
rect 3240 6384 3292 6390
rect 3240 6326 3292 6332
rect 3332 6384 3384 6390
rect 3332 6326 3384 6332
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3146 4040 3202 4049
rect 3146 3975 3202 3984
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3252 3126 3280 3878
rect 3344 3398 3372 5646
rect 3436 3466 3464 6598
rect 3528 5166 3556 9522
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3804 8090 3832 8434
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3608 6724 3660 6730
rect 3608 6666 3660 6672
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 3528 3398 3556 4966
rect 3620 4282 3648 6666
rect 3712 5234 3740 7686
rect 3896 7546 3924 17002
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 14074 4016 14350
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4080 10130 4108 17478
rect 4632 16998 4660 18226
rect 4724 17746 4752 18652
rect 4816 18222 4844 18770
rect 5092 18358 5120 19722
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5184 19446 5212 19654
rect 5172 19440 5224 19446
rect 5172 19382 5224 19388
rect 5368 18698 5396 19722
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 5080 18352 5132 18358
rect 5080 18294 5132 18300
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16658 4660 16934
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15366 4660 15846
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13184 4672 13190
rect 4724 13172 4752 16934
rect 4816 15978 4844 18158
rect 5368 16998 5396 18634
rect 5460 17338 5488 19858
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5552 17882 5580 18090
rect 5644 18086 5672 20742
rect 5828 20534 5856 33895
rect 6012 32502 6040 38966
rect 6104 38554 6132 38966
rect 6656 38962 6684 39238
rect 6748 39001 6776 39986
rect 6734 38992 6790 39001
rect 6644 38956 6696 38962
rect 6734 38927 6736 38936
rect 6644 38898 6696 38904
rect 6788 38927 6790 38936
rect 6736 38898 6788 38904
rect 6092 38548 6144 38554
rect 6092 38490 6144 38496
rect 6104 37262 6132 38490
rect 6092 37256 6144 37262
rect 6092 37198 6144 37204
rect 6656 36854 6684 38898
rect 6748 38554 6776 38898
rect 6736 38548 6788 38554
rect 6736 38490 6788 38496
rect 6736 38276 6788 38282
rect 6736 38218 6788 38224
rect 6748 37670 6776 38218
rect 6736 37664 6788 37670
rect 6736 37606 6788 37612
rect 6644 36848 6696 36854
rect 6644 36790 6696 36796
rect 6748 33658 6776 37606
rect 7104 37188 7156 37194
rect 7104 37130 7156 37136
rect 6920 36576 6972 36582
rect 6920 36518 6972 36524
rect 6828 35080 6880 35086
rect 6828 35022 6880 35028
rect 6736 33652 6788 33658
rect 6736 33594 6788 33600
rect 6460 33584 6512 33590
rect 6460 33526 6512 33532
rect 6472 32570 6500 33526
rect 6748 32910 6776 33594
rect 6736 32904 6788 32910
rect 6736 32846 6788 32852
rect 6840 32842 6868 35022
rect 6828 32836 6880 32842
rect 6828 32778 6880 32784
rect 6460 32564 6512 32570
rect 6460 32506 6512 32512
rect 6736 32564 6788 32570
rect 6736 32506 6788 32512
rect 6000 32496 6052 32502
rect 6000 32438 6052 32444
rect 6012 31822 6040 32438
rect 6748 32026 6776 32506
rect 6840 32366 6868 32778
rect 6828 32360 6880 32366
rect 6828 32302 6880 32308
rect 6736 32020 6788 32026
rect 6736 31962 6788 31968
rect 6184 31952 6236 31958
rect 6184 31894 6236 31900
rect 6000 31816 6052 31822
rect 6000 31758 6052 31764
rect 6196 31754 6224 31894
rect 6748 31822 6776 31962
rect 6840 31958 6868 32302
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6736 31816 6788 31822
rect 6736 31758 6788 31764
rect 6196 31726 6408 31754
rect 6184 31680 6236 31686
rect 6184 31622 6236 31628
rect 6196 31414 6224 31622
rect 6184 31408 6236 31414
rect 6184 31350 6236 31356
rect 6380 31278 6408 31726
rect 6736 31476 6788 31482
rect 6736 31418 6788 31424
rect 6368 31272 6420 31278
rect 6368 31214 6420 31220
rect 6380 30938 6408 31214
rect 6368 30932 6420 30938
rect 6368 30874 6420 30880
rect 6748 30598 6776 31418
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 6368 28416 6420 28422
rect 6368 28358 6420 28364
rect 6380 28082 6408 28358
rect 6748 28150 6776 30534
rect 6736 28144 6788 28150
rect 6736 28086 6788 28092
rect 6368 28076 6420 28082
rect 6368 28018 6420 28024
rect 6460 28076 6512 28082
rect 6460 28018 6512 28024
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6472 27470 6500 28018
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6472 27130 6500 27406
rect 6656 27402 6684 28018
rect 6840 27606 6868 28018
rect 6828 27600 6880 27606
rect 6828 27542 6880 27548
rect 6644 27396 6696 27402
rect 6644 27338 6696 27344
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6460 27124 6512 27130
rect 6460 27066 6512 27072
rect 6092 26784 6144 26790
rect 6092 26726 6144 26732
rect 6104 26518 6132 26726
rect 6092 26512 6144 26518
rect 6092 26454 6144 26460
rect 6104 26382 6132 26454
rect 6092 26376 6144 26382
rect 6092 26318 6144 26324
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6288 26042 6316 26318
rect 6552 26308 6604 26314
rect 6552 26250 6604 26256
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 6184 25696 6236 25702
rect 6184 25638 6236 25644
rect 6092 23656 6144 23662
rect 6092 23598 6144 23604
rect 6104 22030 6132 23598
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 5908 21888 5960 21894
rect 5908 21830 5960 21836
rect 5920 21486 5948 21830
rect 6012 21690 6040 21898
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5908 21480 5960 21486
rect 5908 21422 5960 21428
rect 6000 21140 6052 21146
rect 6000 21082 6052 21088
rect 5816 20528 5868 20534
rect 5816 20470 5868 20476
rect 5908 18692 5960 18698
rect 5908 18634 5960 18640
rect 5920 18290 5948 18634
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 4804 15360 4856 15366
rect 4802 15328 4804 15337
rect 4856 15328 4858 15337
rect 4802 15263 4858 15272
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4816 14006 4844 14282
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4672 13144 4752 13172
rect 4620 13126 4672 13132
rect 4632 12850 4660 13126
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 11642 4660 12786
rect 4816 12594 4844 13942
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4724 12566 4844 12594
rect 4724 11762 4752 12566
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4632 11614 4752 11642
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4356 9586 4384 9930
rect 4540 9674 4568 10066
rect 4540 9646 4660 9674
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 9042 4016 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3988 7886 4016 8774
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3896 6934 3924 7482
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 5710 3924 6734
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3332 3392 3384 3398
rect 3330 3360 3332 3369
rect 3516 3392 3568 3398
rect 3384 3360 3386 3369
rect 3516 3334 3568 3340
rect 3330 3295 3386 3304
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3620 2774 3648 3606
rect 3712 2990 3740 5170
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4214 3924 4966
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3804 3194 3832 4082
rect 3988 3641 4016 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 4080 5914 4108 6802
rect 4632 6118 4660 9646
rect 4724 6186 4752 11614
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4724 5794 4752 6122
rect 4632 5766 4752 5794
rect 4632 5658 4660 5766
rect 4540 5630 4660 5658
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4540 5114 4568 5630
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4632 5370 4660 5510
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4540 5086 4660 5114
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4342 4720 4398 4729
rect 4342 4655 4344 4664
rect 4396 4655 4398 4664
rect 4344 4626 4396 4632
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4080 4146 4108 4218
rect 4632 4146 4660 5086
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3974 3632 4030 3641
rect 3974 3567 4030 3576
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3620 2746 3740 2774
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3712 2378 3740 2746
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4250 2408 4306 2417
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 1582 2272 1638 2281
rect 1582 2207 1638 2216
rect 4080 2038 4108 2382
rect 4250 2343 4306 2352
rect 4264 2310 4292 2343
rect 4252 2304 4304 2310
rect 4252 2246 4304 2252
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 4264 1902 4292 2246
rect 4252 1896 4304 1902
rect 4252 1838 4304 1844
rect 4632 1426 4660 3878
rect 4724 3194 4752 5646
rect 4816 4060 4844 11018
rect 4908 4321 4936 13670
rect 4894 4312 4950 4321
rect 4894 4247 4950 4256
rect 5000 4128 5028 15098
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5184 13530 5212 13874
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 5368 12782 5396 15914
rect 5460 15094 5488 16594
rect 5552 16590 5580 17614
rect 5920 17542 5948 18226
rect 6012 17882 6040 21082
rect 6196 20874 6224 25638
rect 6564 25242 6592 26250
rect 6736 26240 6788 26246
rect 6736 26182 6788 26188
rect 6472 25226 6592 25242
rect 6748 25226 6776 26182
rect 6460 25220 6592 25226
rect 6512 25214 6592 25220
rect 6460 25162 6512 25168
rect 6564 24954 6592 25214
rect 6736 25220 6788 25226
rect 6736 25162 6788 25168
rect 6552 24948 6604 24954
rect 6552 24890 6604 24896
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6288 24614 6316 24754
rect 6840 24698 6868 27270
rect 6932 25906 6960 36518
rect 7116 36378 7144 37130
rect 7104 36372 7156 36378
rect 7104 36314 7156 36320
rect 7012 35012 7064 35018
rect 7012 34954 7064 34960
rect 7024 34746 7052 34954
rect 7012 34740 7064 34746
rect 7012 34682 7064 34688
rect 7208 34678 7236 40394
rect 8116 40384 8168 40390
rect 8116 40326 8168 40332
rect 7656 38888 7708 38894
rect 7708 38836 7788 38842
rect 7656 38830 7788 38836
rect 7668 38814 7788 38830
rect 7564 37120 7616 37126
rect 7564 37062 7616 37068
rect 7576 36854 7604 37062
rect 7564 36848 7616 36854
rect 7564 36790 7616 36796
rect 7288 36780 7340 36786
rect 7288 36722 7340 36728
rect 7300 35698 7328 36722
rect 7656 36576 7708 36582
rect 7656 36518 7708 36524
rect 7668 36174 7696 36518
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 7656 36168 7708 36174
rect 7656 36110 7708 36116
rect 7288 35692 7340 35698
rect 7288 35634 7340 35640
rect 7196 34672 7248 34678
rect 7248 34620 7328 34626
rect 7196 34614 7328 34620
rect 7208 34598 7328 34614
rect 7196 34536 7248 34542
rect 7196 34478 7248 34484
rect 7208 33114 7236 34478
rect 7300 34134 7328 34598
rect 7288 34128 7340 34134
rect 7288 34070 7340 34076
rect 7196 33108 7248 33114
rect 7196 33050 7248 33056
rect 7208 32858 7236 33050
rect 7392 32910 7420 36110
rect 7564 34944 7616 34950
rect 7564 34886 7616 34892
rect 7472 34604 7524 34610
rect 7472 34546 7524 34552
rect 7484 34202 7512 34546
rect 7472 34196 7524 34202
rect 7472 34138 7524 34144
rect 7576 34066 7604 34886
rect 7564 34060 7616 34066
rect 7564 34002 7616 34008
rect 7564 33924 7616 33930
rect 7564 33866 7616 33872
rect 7576 33522 7604 33866
rect 7564 33516 7616 33522
rect 7564 33458 7616 33464
rect 7380 32904 7432 32910
rect 7208 32830 7328 32858
rect 7380 32846 7432 32852
rect 7196 32768 7248 32774
rect 7196 32710 7248 32716
rect 7208 32434 7236 32710
rect 7196 32428 7248 32434
rect 7196 32370 7248 32376
rect 7300 31890 7328 32830
rect 7472 32768 7524 32774
rect 7472 32710 7524 32716
rect 7196 31884 7248 31890
rect 7196 31826 7248 31832
rect 7288 31884 7340 31890
rect 7288 31826 7340 31832
rect 7208 30938 7236 31826
rect 7288 31136 7340 31142
rect 7288 31078 7340 31084
rect 7196 30932 7248 30938
rect 7196 30874 7248 30880
rect 7300 30666 7328 31078
rect 7288 30660 7340 30666
rect 7288 30602 7340 30608
rect 7012 27872 7064 27878
rect 7012 27814 7064 27820
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 7024 24818 7052 27814
rect 7104 27532 7156 27538
rect 7104 27474 7156 27480
rect 7116 27402 7144 27474
rect 7104 27396 7156 27402
rect 7104 27338 7156 27344
rect 7116 27062 7144 27338
rect 7104 27056 7156 27062
rect 7104 26998 7156 27004
rect 7300 25974 7328 30602
rect 7484 29866 7512 32710
rect 7576 32230 7604 33458
rect 7656 32904 7708 32910
rect 7656 32846 7708 32852
rect 7668 32570 7696 32846
rect 7656 32564 7708 32570
rect 7656 32506 7708 32512
rect 7564 32224 7616 32230
rect 7564 32166 7616 32172
rect 7576 31346 7604 32166
rect 7564 31340 7616 31346
rect 7564 31282 7616 31288
rect 7576 30734 7604 31282
rect 7564 30728 7616 30734
rect 7564 30670 7616 30676
rect 7484 29838 7604 29866
rect 7472 29776 7524 29782
rect 7472 29718 7524 29724
rect 7484 29034 7512 29718
rect 7472 29028 7524 29034
rect 7472 28970 7524 28976
rect 7380 28960 7432 28966
rect 7380 28902 7432 28908
rect 7392 26466 7420 28902
rect 7576 28762 7604 29838
rect 7760 29782 7788 38814
rect 8128 37262 8156 40326
rect 8956 40050 8984 40870
rect 8944 40044 8996 40050
rect 8944 39986 8996 39992
rect 8576 39840 8628 39846
rect 8576 39782 8628 39788
rect 8588 38350 8616 39782
rect 9036 39432 9088 39438
rect 9036 39374 9088 39380
rect 9048 39030 9076 39374
rect 9036 39024 9088 39030
rect 9036 38966 9088 38972
rect 9416 38554 9444 41074
rect 9692 41070 9720 41414
rect 9956 41268 10008 41274
rect 9956 41210 10008 41216
rect 9864 41200 9916 41206
rect 9864 41142 9916 41148
rect 9680 41064 9732 41070
rect 9680 41006 9732 41012
rect 9692 40662 9720 41006
rect 9680 40656 9732 40662
rect 9680 40598 9732 40604
rect 9876 40458 9904 41142
rect 9968 40526 9996 41210
rect 10324 41132 10376 41138
rect 10324 41074 10376 41080
rect 10876 41132 10928 41138
rect 10876 41074 10928 41080
rect 10140 40928 10192 40934
rect 10140 40870 10192 40876
rect 10152 40526 10180 40870
rect 9956 40520 10008 40526
rect 9956 40462 10008 40468
rect 10140 40520 10192 40526
rect 10140 40462 10192 40468
rect 9864 40452 9916 40458
rect 9864 40394 9916 40400
rect 9680 40384 9732 40390
rect 9680 40326 9732 40332
rect 9692 39030 9720 40326
rect 9876 40118 9904 40394
rect 9864 40112 9916 40118
rect 9864 40054 9916 40060
rect 9772 39840 9824 39846
rect 9772 39782 9824 39788
rect 9784 39438 9812 39782
rect 9772 39432 9824 39438
rect 9772 39374 9824 39380
rect 9680 39024 9732 39030
rect 9680 38966 9732 38972
rect 9404 38548 9456 38554
rect 9404 38490 9456 38496
rect 8576 38344 8628 38350
rect 8576 38286 8628 38292
rect 9312 38344 9364 38350
rect 9312 38286 9364 38292
rect 9324 37874 9352 38286
rect 9680 38276 9732 38282
rect 9680 38218 9732 38224
rect 9312 37868 9364 37874
rect 9312 37810 9364 37816
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 8024 37188 8076 37194
rect 8024 37130 8076 37136
rect 8036 36718 8064 37130
rect 8220 36922 8248 37198
rect 8944 37120 8996 37126
rect 8944 37062 8996 37068
rect 8208 36916 8260 36922
rect 8208 36858 8260 36864
rect 8024 36712 8076 36718
rect 8024 36654 8076 36660
rect 8116 36304 8168 36310
rect 8116 36246 8168 36252
rect 8128 35222 8156 36246
rect 8208 36168 8260 36174
rect 8208 36110 8260 36116
rect 8220 35630 8248 36110
rect 8208 35624 8260 35630
rect 8208 35566 8260 35572
rect 8116 35216 8168 35222
rect 8116 35158 8168 35164
rect 7932 34128 7984 34134
rect 7932 34070 7984 34076
rect 7748 29776 7800 29782
rect 7748 29718 7800 29724
rect 7748 29504 7800 29510
rect 7748 29446 7800 29452
rect 7760 29170 7788 29446
rect 7748 29164 7800 29170
rect 7748 29106 7800 29112
rect 7564 28756 7616 28762
rect 7564 28698 7616 28704
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 7484 26586 7512 26930
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7576 26518 7604 28698
rect 7656 28484 7708 28490
rect 7656 28426 7708 28432
rect 7668 27674 7696 28426
rect 7656 27668 7708 27674
rect 7656 27610 7708 27616
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7668 26518 7696 27270
rect 7760 27062 7788 29106
rect 7748 27056 7800 27062
rect 7748 26998 7800 27004
rect 7748 26920 7800 26926
rect 7748 26862 7800 26868
rect 7564 26512 7616 26518
rect 7392 26438 7512 26466
rect 7564 26454 7616 26460
rect 7656 26512 7708 26518
rect 7656 26454 7708 26460
rect 7484 26382 7512 26438
rect 7472 26376 7524 26382
rect 7472 26318 7524 26324
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 7104 25900 7156 25906
rect 7104 25842 7156 25848
rect 7116 25498 7144 25842
rect 7484 25702 7512 26318
rect 7472 25696 7524 25702
rect 7472 25638 7524 25644
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 7760 25294 7788 26862
rect 7748 25288 7800 25294
rect 7748 25230 7800 25236
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7944 24750 7972 34070
rect 8116 33312 8168 33318
rect 8116 33254 8168 33260
rect 8128 32978 8156 33254
rect 8116 32972 8168 32978
rect 8116 32914 8168 32920
rect 7932 24744 7984 24750
rect 6840 24670 7144 24698
rect 7932 24686 7984 24692
rect 6276 24608 6328 24614
rect 6276 24550 6328 24556
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6288 20058 6316 24550
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6380 22030 6408 22374
rect 6840 22234 6868 22578
rect 6828 22228 6880 22234
rect 6828 22170 6880 22176
rect 6363 22024 6415 22030
rect 6363 21966 6415 21972
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6380 19310 6408 21422
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6564 20466 6592 20742
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6564 19854 6592 20402
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6840 19718 6868 20334
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6552 19440 6604 19446
rect 6552 19382 6604 19388
rect 6368 19304 6420 19310
rect 6368 19246 6420 19252
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 6276 17536 6328 17542
rect 6276 17478 6328 17484
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5552 16046 5580 16526
rect 5736 16454 5764 17478
rect 5920 16998 5948 17478
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 16182 5764 16390
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 13938 5672 14758
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5644 13394 5672 13874
rect 5736 13870 5764 16118
rect 5724 13864 5776 13870
rect 5724 13806 5776 13812
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5540 13184 5592 13190
rect 5540 13126 5592 13132
rect 5552 12986 5580 13126
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5368 10266 5396 12718
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 12102 5580 12242
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5552 11762 5580 12038
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5736 11626 5764 13806
rect 5920 12434 5948 16934
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 5920 12406 6040 12434
rect 5540 11620 5592 11626
rect 5540 11562 5592 11568
rect 5724 11620 5776 11626
rect 5724 11562 5776 11568
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5080 6724 5132 6730
rect 5080 6666 5132 6672
rect 5092 5370 5120 6666
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5000 4100 5120 4128
rect 4816 4032 5028 4060
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4816 3738 4844 3878
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4620 1420 4672 1426
rect 4620 1362 4672 1368
rect 4816 1358 4844 2994
rect 5000 2446 5028 4032
rect 5092 3942 5120 4100
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5184 3482 5212 9046
rect 5368 9042 5396 10202
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5276 8362 5304 8774
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5460 8242 5488 10950
rect 5552 9586 5580 11562
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5276 8214 5488 8242
rect 5276 4622 5304 8214
rect 5552 6866 5580 8910
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5644 8634 5672 8842
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5736 8480 5764 9454
rect 6012 9042 6040 12406
rect 6196 12306 6224 13330
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 6196 10538 6224 12242
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6196 9382 6224 10474
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5828 8634 5856 8842
rect 5920 8634 5948 8910
rect 6196 8838 6224 8978
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 8492 5868 8498
rect 5736 8452 5816 8480
rect 5816 8434 5868 8440
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5632 7336 5684 7342
rect 5630 7304 5632 7313
rect 5684 7304 5686 7313
rect 5630 7239 5686 7248
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5368 5574 5396 6190
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5370 5580 5510
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5264 4480 5316 4486
rect 5262 4448 5264 4457
rect 5316 4448 5318 4457
rect 5262 4383 5318 4392
rect 5262 4312 5318 4321
rect 5262 4247 5318 4256
rect 5092 3466 5212 3482
rect 5080 3460 5212 3466
rect 5132 3454 5212 3460
rect 5080 3402 5132 3408
rect 5276 3058 5304 4247
rect 5368 4162 5396 5170
rect 5460 4434 5488 5170
rect 5552 4622 5580 5306
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5460 4406 5580 4434
rect 5368 4134 5488 4162
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5368 1630 5396 2858
rect 5460 2774 5488 4134
rect 5552 3942 5580 4406
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5644 2854 5672 6054
rect 5736 5778 5764 7346
rect 5828 7342 5856 8434
rect 6104 7886 6132 8774
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5828 6730 5856 7278
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 6288 6474 6316 17478
rect 6564 14074 6592 19382
rect 6840 18834 6868 19654
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6840 17542 6868 18770
rect 6932 18426 6960 19314
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 7024 17626 7052 18702
rect 6932 17598 7052 17626
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6564 13326 6592 14010
rect 6840 13870 6868 15982
rect 6932 15910 6960 17598
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 7024 16454 7052 17138
rect 7012 16448 7064 16454
rect 7012 16390 7064 16396
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6932 15162 6960 15302
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6932 14278 6960 14758
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6380 6798 6408 7754
rect 6460 7336 6512 7342
rect 6460 7278 6512 7284
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6196 6446 6316 6474
rect 6196 5846 6224 6446
rect 6276 6316 6328 6322
rect 6276 6258 6328 6264
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 5724 5772 5776 5778
rect 5724 5714 5776 5720
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5736 4690 5764 5034
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5828 3534 5856 5646
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6012 4842 6040 5238
rect 6104 5234 6132 5646
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6012 4826 6132 4842
rect 6012 4820 6144 4826
rect 6012 4814 6092 4820
rect 6092 4762 6144 4768
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5460 2746 5580 2774
rect 5552 2666 5580 2746
rect 5552 2638 5672 2666
rect 5538 2408 5594 2417
rect 5538 2343 5594 2352
rect 5356 1624 5408 1630
rect 5356 1566 5408 1572
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 5552 800 5580 2343
rect 5644 800 5672 2638
rect 5814 2544 5870 2553
rect 5814 2479 5870 2488
rect 5828 2446 5856 2479
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 2106 5856 2246
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 5920 1834 5948 4694
rect 6196 4622 6224 5510
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6288 4434 6316 6258
rect 6012 4406 6316 4434
rect 5908 1828 5960 1834
rect 5908 1770 5960 1776
rect 6012 1714 6040 4406
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6288 3670 6316 4218
rect 6276 3664 6328 3670
rect 6182 3632 6238 3641
rect 6276 3606 6328 3612
rect 6182 3567 6184 3576
rect 6236 3567 6238 3576
rect 6184 3538 6236 3544
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 5828 1686 6040 1714
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 5736 800 5764 1362
rect 5828 800 5856 1686
rect 5908 1624 5960 1630
rect 6104 1578 6132 2926
rect 5908 1566 5960 1572
rect 5920 800 5948 1566
rect 6012 1550 6132 1578
rect 6012 800 6040 1550
rect 6196 1442 6224 3538
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6104 1414 6224 1442
rect 6104 800 6132 1414
rect 6184 1352 6236 1358
rect 6184 1294 6236 1300
rect 6196 800 6224 1294
rect 6288 800 6316 2586
rect 6380 800 6408 6734
rect 6472 6458 6500 7278
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6564 6390 6592 13262
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6656 10674 6684 11698
rect 6748 11694 6776 12786
rect 6840 11830 6868 13806
rect 7024 13734 7052 16390
rect 7116 15910 7144 24670
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7392 21690 7420 23054
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7668 22574 7696 22918
rect 7656 22568 7708 22574
rect 7656 22510 7708 22516
rect 7668 22030 7696 22510
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7380 21684 7432 21690
rect 7380 21626 7432 21632
rect 7760 21418 7788 21898
rect 7748 21412 7800 21418
rect 7748 21354 7800 21360
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 18290 7420 18566
rect 7668 18358 7696 19110
rect 7760 18970 7788 19178
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7208 17134 7236 18158
rect 7668 17542 7696 18294
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7208 14958 7236 17070
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16590 7420 16934
rect 7380 16584 7432 16590
rect 7380 16526 7432 16532
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7300 15162 7328 15370
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7012 12640 7064 12646
rect 7012 12582 7064 12588
rect 7024 12238 7052 12582
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 9586 6776 10542
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6748 8294 6776 9522
rect 6840 8401 6868 9862
rect 6932 9382 6960 11494
rect 7024 11082 7052 12174
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 7116 10849 7144 12038
rect 7208 11286 7236 14894
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7102 10840 7158 10849
rect 7102 10775 7158 10784
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6826 8392 6882 8401
rect 6826 8327 6882 8336
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7478 6960 8230
rect 7024 7886 7052 9454
rect 7208 9042 7236 11222
rect 7300 11150 7328 14214
rect 7484 11150 7512 15846
rect 7668 14550 7696 17478
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7852 16250 7880 17070
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7944 14822 7972 24346
rect 8024 22568 8076 22574
rect 8024 22510 8076 22516
rect 8036 22438 8064 22510
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8128 22234 8156 32914
rect 8220 31346 8248 35566
rect 8956 33998 8984 37062
rect 9692 36038 9720 38218
rect 9772 36712 9824 36718
rect 9772 36654 9824 36660
rect 9784 36242 9812 36654
rect 9772 36236 9824 36242
rect 9772 36178 9824 36184
rect 9680 36032 9732 36038
rect 9680 35974 9732 35980
rect 9692 35766 9720 35974
rect 9680 35760 9732 35766
rect 9680 35702 9732 35708
rect 9220 35624 9272 35630
rect 9220 35566 9272 35572
rect 9232 35086 9260 35566
rect 9496 35556 9548 35562
rect 9496 35498 9548 35504
rect 9508 35086 9536 35498
rect 9784 35154 9812 36178
rect 9876 35698 9904 40054
rect 10336 38758 10364 41074
rect 10416 40996 10468 41002
rect 10416 40938 10468 40944
rect 10428 40526 10456 40938
rect 10888 40526 10916 41074
rect 10416 40520 10468 40526
rect 10416 40462 10468 40468
rect 10876 40520 10928 40526
rect 10876 40462 10928 40468
rect 10428 40050 10456 40462
rect 10508 40452 10560 40458
rect 10508 40394 10560 40400
rect 10416 40044 10468 40050
rect 10416 39986 10468 39992
rect 10324 38752 10376 38758
rect 10324 38694 10376 38700
rect 10336 38350 10364 38694
rect 10324 38344 10376 38350
rect 10324 38286 10376 38292
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 9864 35692 9916 35698
rect 9864 35634 9916 35640
rect 9772 35148 9824 35154
rect 9772 35090 9824 35096
rect 9220 35080 9272 35086
rect 9496 35080 9548 35086
rect 9272 35040 9352 35068
rect 9220 35022 9272 35028
rect 8944 33992 8996 33998
rect 8944 33934 8996 33940
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 8852 33856 8904 33862
rect 8852 33798 8904 33804
rect 8484 31816 8536 31822
rect 8484 31758 8536 31764
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8220 29850 8248 31282
rect 8392 31136 8444 31142
rect 8392 31078 8444 31084
rect 8208 29844 8260 29850
rect 8208 29786 8260 29792
rect 8220 29238 8248 29786
rect 8208 29232 8260 29238
rect 8208 29174 8260 29180
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8220 25702 8248 26318
rect 8300 25764 8352 25770
rect 8300 25706 8352 25712
rect 8208 25696 8260 25702
rect 8208 25638 8260 25644
rect 8220 24954 8248 25638
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 8208 24744 8260 24750
rect 8208 24686 8260 24692
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 8128 21894 8156 22170
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8128 19242 8156 21830
rect 8220 21146 8248 24686
rect 8208 21140 8260 21146
rect 8208 21082 8260 21088
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8208 19168 8260 19174
rect 8208 19110 8260 19116
rect 8116 18896 8168 18902
rect 8116 18838 8168 18844
rect 8128 18630 8156 18838
rect 8220 18766 8248 19110
rect 8312 18970 8340 25706
rect 8404 20602 8432 31078
rect 8496 30394 8524 31758
rect 8484 30388 8536 30394
rect 8484 30330 8536 30336
rect 8496 26858 8524 30330
rect 8576 29232 8628 29238
rect 8574 29200 8576 29209
rect 8628 29200 8630 29209
rect 8574 29135 8630 29144
rect 8484 26852 8536 26858
rect 8484 26794 8536 26800
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8392 20596 8444 20602
rect 8392 20538 8444 20544
rect 8496 19174 8524 20742
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8298 18864 8354 18873
rect 8298 18799 8300 18808
rect 8352 18799 8354 18808
rect 8300 18770 8352 18776
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 8312 18426 8340 18770
rect 8404 18766 8432 18906
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8588 18698 8616 23802
rect 8668 22704 8720 22710
rect 8668 22646 8720 22652
rect 8576 18692 8628 18698
rect 8576 18634 8628 18640
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8128 17202 8156 18226
rect 8116 17196 8168 17202
rect 8168 17156 8248 17184
rect 8116 17138 8168 17144
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 8128 15910 8156 16050
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 7932 14816 7984 14822
rect 7932 14758 7984 14764
rect 7656 14544 7708 14550
rect 7656 14486 7708 14492
rect 8024 13864 8076 13870
rect 8128 13841 8156 15846
rect 8024 13806 8076 13812
rect 8114 13832 8170 13841
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7576 12442 7604 12786
rect 7564 12436 7616 12442
rect 7564 12378 7616 12384
rect 8036 12306 8064 13806
rect 8114 13767 8170 13776
rect 8220 13326 8248 17156
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8312 13394 8340 15438
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8312 12850 8340 13330
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 12374 8340 12786
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8404 12238 8432 13262
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8024 11756 8076 11762
rect 8024 11698 8076 11704
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7576 11218 7604 11494
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7852 11150 7880 11494
rect 8036 11354 8064 11698
rect 8208 11552 8260 11558
rect 8260 11500 8340 11506
rect 8208 11494 8340 11500
rect 8220 11478 8340 11494
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7852 11014 7880 11086
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 8128 9450 8156 11018
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7300 8974 7328 9386
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7288 8968 7340 8974
rect 7288 8910 7340 8916
rect 7668 8362 7696 9318
rect 8220 8430 8248 9590
rect 8312 8906 8340 11478
rect 8496 9110 8524 15302
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8300 8900 8352 8906
rect 8300 8842 8352 8848
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6748 6866 6776 7278
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6552 6384 6604 6390
rect 6552 6326 6604 6332
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6564 5574 6592 5782
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 6564 4554 6592 5034
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6564 4214 6592 4490
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6458 4040 6514 4049
rect 6458 3975 6514 3984
rect 6472 3058 6500 3975
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6472 800 6500 2994
rect 6564 2854 6592 4150
rect 6656 3942 6684 6598
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6748 5234 6776 5646
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 5030 6776 5170
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4622 6776 4966
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6840 4554 6868 6598
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6840 4078 6868 4490
rect 6932 4486 6960 7414
rect 7024 6202 7052 7822
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 6798 7236 7686
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7024 6174 7144 6202
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6644 3936 6696 3942
rect 7024 3890 7052 4694
rect 7116 4282 7144 6174
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7102 4040 7158 4049
rect 7102 3975 7158 3984
rect 6644 3878 6696 3884
rect 6932 3862 7052 3890
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6748 1986 6776 3606
rect 6826 3224 6882 3233
rect 6932 3194 6960 3862
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6826 3159 6828 3168
rect 6880 3159 6882 3168
rect 6920 3188 6972 3194
rect 6828 3130 6880 3136
rect 6920 3130 6972 3136
rect 6918 2952 6974 2961
rect 6918 2887 6974 2896
rect 6564 1958 6776 1986
rect 6828 1964 6880 1970
rect 6564 800 6592 1958
rect 6828 1906 6880 1912
rect 6644 1828 6696 1834
rect 6644 1770 6696 1776
rect 6656 800 6684 1770
rect 6840 800 6868 1906
rect 6932 800 6960 2887
rect 7024 800 7052 3674
rect 7116 2446 7144 3975
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7116 1970 7144 2382
rect 7104 1964 7156 1970
rect 7104 1906 7156 1912
rect 7208 800 7236 6734
rect 7300 6322 7328 7754
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7300 2961 7328 6258
rect 7484 4978 7512 8026
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 5234 7604 6054
rect 7668 5914 7696 8298
rect 8036 8090 8064 8366
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8036 7410 8064 8026
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7760 5710 7788 7142
rect 7852 6798 7880 7210
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7392 4950 7512 4978
rect 7392 4078 7420 4950
rect 7576 4842 7604 5170
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7484 4826 7604 4842
rect 7472 4820 7604 4826
rect 7524 4814 7604 4820
rect 7472 4762 7524 4768
rect 7484 4146 7512 4762
rect 7668 4706 7696 5102
rect 7576 4678 7696 4706
rect 7576 4622 7604 4678
rect 7564 4616 7616 4622
rect 7760 4604 7788 5646
rect 7564 4558 7616 4564
rect 7668 4576 7788 4604
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7380 4072 7432 4078
rect 7576 4026 7604 4558
rect 7380 4014 7432 4020
rect 7484 4010 7604 4026
rect 7472 4004 7604 4010
rect 7524 3998 7604 4004
rect 7472 3946 7524 3952
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3126 7420 3878
rect 7484 3670 7512 3946
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7576 3058 7604 3878
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7286 2952 7342 2961
rect 7668 2938 7696 4576
rect 7286 2887 7342 2896
rect 7484 2910 7696 2938
rect 7748 2916 7800 2922
rect 7484 2774 7512 2910
rect 7748 2858 7800 2864
rect 7300 2746 7512 2774
rect 7654 2816 7710 2825
rect 7654 2751 7710 2760
rect 7300 800 7328 2746
rect 7562 2680 7618 2689
rect 7562 2615 7618 2624
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7392 800 7420 2518
rect 7576 800 7604 2615
rect 7668 2514 7696 2751
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 7656 2032 7708 2038
rect 7656 1974 7708 1980
rect 7668 800 7696 1974
rect 7760 800 7788 2858
rect 7852 800 7880 6734
rect 8312 6730 8340 8842
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 7750 8432 8434
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7410 8432 7686
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 7313 8432 7346
rect 8390 7304 8446 7313
rect 8390 7239 8446 7248
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6322 8064 6598
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7944 2961 7972 5578
rect 8036 3602 8064 6258
rect 8404 6186 8432 6258
rect 8392 6180 8444 6186
rect 8392 6122 8444 6128
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8128 5574 8156 5850
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8128 4826 8156 5102
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8220 4706 8248 5782
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8128 4678 8248 4706
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 7930 2952 7986 2961
rect 8036 2922 8064 3130
rect 7930 2887 7986 2896
rect 8024 2916 8076 2922
rect 8024 2858 8076 2864
rect 8036 2802 8064 2858
rect 7944 2774 8064 2802
rect 7944 800 7972 2774
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8036 800 8064 2246
rect 8128 800 8156 4678
rect 8312 4010 8340 5646
rect 8404 4078 8432 6122
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5234 8524 5510
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8496 4690 8524 5170
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8588 4078 8616 13806
rect 8680 8634 8708 22646
rect 8864 20058 8892 33798
rect 9048 32502 9076 33934
rect 9220 33924 9272 33930
rect 9220 33866 9272 33872
rect 9232 33658 9260 33866
rect 9220 33652 9272 33658
rect 9220 33594 9272 33600
rect 9128 32564 9180 32570
rect 9128 32506 9180 32512
rect 9036 32496 9088 32502
rect 9036 32438 9088 32444
rect 9140 31142 9168 32506
rect 9128 31136 9180 31142
rect 9128 31078 9180 31084
rect 9324 30190 9352 35040
rect 9496 35022 9548 35028
rect 9876 35018 9904 35634
rect 9864 35012 9916 35018
rect 9864 34954 9916 34960
rect 9876 34542 9904 34954
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9956 33108 10008 33114
rect 9956 33050 10008 33056
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9692 31278 9720 32370
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9680 31272 9732 31278
rect 9680 31214 9732 31220
rect 9312 30184 9364 30190
rect 9364 30144 9444 30172
rect 9312 30126 9364 30132
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9324 29714 9352 29990
rect 9312 29708 9364 29714
rect 9312 29650 9364 29656
rect 9128 29164 9180 29170
rect 9128 29106 9180 29112
rect 9220 29164 9272 29170
rect 9272 29124 9352 29152
rect 9220 29106 9272 29112
rect 9036 28960 9088 28966
rect 9036 28902 9088 28908
rect 9048 28490 9076 28902
rect 9140 28762 9168 29106
rect 9220 29028 9272 29034
rect 9220 28970 9272 28976
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 9036 28484 9088 28490
rect 9036 28426 9088 28432
rect 9232 28150 9260 28970
rect 9324 28966 9352 29124
rect 9416 29034 9444 30144
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 9404 29028 9456 29034
rect 9404 28970 9456 28976
rect 9312 28960 9364 28966
rect 9312 28902 9364 28908
rect 9416 28218 9444 28970
rect 9508 28422 9536 29582
rect 9586 29200 9642 29209
rect 9586 29135 9588 29144
rect 9640 29135 9642 29144
rect 9588 29106 9640 29112
rect 9496 28416 9548 28422
rect 9496 28358 9548 28364
rect 9404 28212 9456 28218
rect 9404 28154 9456 28160
rect 9220 28144 9272 28150
rect 9220 28086 9272 28092
rect 9508 28082 9536 28358
rect 8944 28076 8996 28082
rect 8944 28018 8996 28024
rect 9496 28076 9548 28082
rect 9496 28018 9548 28024
rect 8956 27878 8984 28018
rect 8944 27872 8996 27878
rect 8944 27814 8996 27820
rect 8956 27470 8984 27814
rect 9312 27600 9364 27606
rect 9312 27542 9364 27548
rect 8944 27464 8996 27470
rect 8944 27406 8996 27412
rect 8956 22574 8984 27406
rect 9324 26994 9352 27542
rect 9508 27470 9536 28018
rect 9692 27606 9720 31214
rect 9876 30326 9904 31758
rect 9864 30320 9916 30326
rect 9864 30262 9916 30268
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9784 29170 9812 29446
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9404 27464 9456 27470
rect 9404 27406 9456 27412
rect 9496 27464 9548 27470
rect 9496 27406 9548 27412
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9324 25974 9352 26930
rect 9416 25974 9444 27406
rect 9784 26926 9812 28494
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9772 26920 9824 26926
rect 9772 26862 9824 26868
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 9312 25968 9364 25974
rect 9312 25910 9364 25916
rect 9404 25968 9456 25974
rect 9404 25910 9456 25916
rect 9508 25906 9536 25978
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9036 24744 9088 24750
rect 9508 24698 9536 25842
rect 9876 25838 9904 26930
rect 9968 26790 9996 33050
rect 10244 32910 10272 36722
rect 10428 36718 10456 39986
rect 10520 39302 10548 40394
rect 10784 40384 10836 40390
rect 10784 40326 10836 40332
rect 10796 40118 10824 40326
rect 10784 40112 10836 40118
rect 10784 40054 10836 40060
rect 10508 39296 10560 39302
rect 10508 39238 10560 39244
rect 10520 37806 10548 39238
rect 10888 38282 10916 40462
rect 11060 40384 11112 40390
rect 11060 40326 11112 40332
rect 10968 39840 11020 39846
rect 10968 39782 11020 39788
rect 10980 38758 11008 39782
rect 11072 39642 11100 40326
rect 11716 39642 11744 41482
rect 12452 41478 12480 42026
rect 12348 41472 12400 41478
rect 12348 41414 12400 41420
rect 12440 41472 12492 41478
rect 12440 41414 12492 41420
rect 11796 40928 11848 40934
rect 11796 40870 11848 40876
rect 11808 40118 11836 40870
rect 11796 40112 11848 40118
rect 11796 40054 11848 40060
rect 11060 39636 11112 39642
rect 11060 39578 11112 39584
rect 11704 39636 11756 39642
rect 11704 39578 11756 39584
rect 10968 38752 11020 38758
rect 10968 38694 11020 38700
rect 10876 38276 10928 38282
rect 10876 38218 10928 38224
rect 11716 38010 11744 39578
rect 12360 39438 12388 41414
rect 12348 39432 12400 39438
rect 12348 39374 12400 39380
rect 12452 39098 12480 41414
rect 12544 40186 12572 42162
rect 12716 42152 12768 42158
rect 12716 42094 12768 42100
rect 12728 41750 12756 42094
rect 12808 42016 12860 42022
rect 12808 41958 12860 41964
rect 12716 41744 12768 41750
rect 12716 41686 12768 41692
rect 12728 41018 12756 41686
rect 12820 41138 12848 41958
rect 12898 41712 12954 41721
rect 12898 41647 12900 41656
rect 12952 41647 12954 41656
rect 12900 41618 12952 41624
rect 15028 41614 15056 42162
rect 12992 41608 13044 41614
rect 12992 41550 13044 41556
rect 14740 41608 14792 41614
rect 14740 41550 14792 41556
rect 15016 41608 15068 41614
rect 15016 41550 15068 41556
rect 13004 41138 13032 41550
rect 13820 41540 13872 41546
rect 13820 41482 13872 41488
rect 12808 41132 12860 41138
rect 12808 41074 12860 41080
rect 12992 41132 13044 41138
rect 12992 41074 13044 41080
rect 12900 41064 12952 41070
rect 12728 41012 12900 41018
rect 12728 41006 12952 41012
rect 12728 40990 12940 41006
rect 13004 40594 13032 41074
rect 12992 40588 13044 40594
rect 12992 40530 13044 40536
rect 13176 40452 13228 40458
rect 13176 40394 13228 40400
rect 12532 40180 12584 40186
rect 12532 40122 12584 40128
rect 12900 40180 12952 40186
rect 12900 40122 12952 40128
rect 12624 39840 12676 39846
rect 12624 39782 12676 39788
rect 12636 39438 12664 39782
rect 12624 39432 12676 39438
rect 12624 39374 12676 39380
rect 12440 39092 12492 39098
rect 12440 39034 12492 39040
rect 12532 38956 12584 38962
rect 12532 38898 12584 38904
rect 12544 38418 12572 38898
rect 12532 38412 12584 38418
rect 12532 38354 12584 38360
rect 11704 38004 11756 38010
rect 11704 37946 11756 37952
rect 11704 37868 11756 37874
rect 11704 37810 11756 37816
rect 12256 37868 12308 37874
rect 12256 37810 12308 37816
rect 10508 37800 10560 37806
rect 10508 37742 10560 37748
rect 11336 37664 11388 37670
rect 11336 37606 11388 37612
rect 11348 37194 11376 37606
rect 11716 37262 11744 37810
rect 12268 37738 12296 37810
rect 12256 37732 12308 37738
rect 12256 37674 12308 37680
rect 11704 37256 11756 37262
rect 11704 37198 11756 37204
rect 11336 37188 11388 37194
rect 11336 37130 11388 37136
rect 11716 36854 11744 37198
rect 12268 36922 12296 37674
rect 12348 37460 12400 37466
rect 12348 37402 12400 37408
rect 12360 37194 12388 37402
rect 12348 37188 12400 37194
rect 12348 37130 12400 37136
rect 12256 36916 12308 36922
rect 12256 36858 12308 36864
rect 11704 36848 11756 36854
rect 11704 36790 11756 36796
rect 10416 36712 10468 36718
rect 10416 36654 10468 36660
rect 10324 36100 10376 36106
rect 10324 36042 10376 36048
rect 10416 36100 10468 36106
rect 10416 36042 10468 36048
rect 10336 34746 10364 36042
rect 10428 35154 10456 36042
rect 11428 36032 11480 36038
rect 11428 35974 11480 35980
rect 11440 35834 11468 35974
rect 11428 35828 11480 35834
rect 11428 35770 11480 35776
rect 12256 35828 12308 35834
rect 12256 35770 12308 35776
rect 11796 35692 11848 35698
rect 11796 35634 11848 35640
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10784 35488 10836 35494
rect 10784 35430 10836 35436
rect 10416 35148 10468 35154
rect 10416 35090 10468 35096
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10428 33114 10456 34682
rect 10508 34672 10560 34678
rect 10508 34614 10560 34620
rect 10520 34202 10548 34614
rect 10796 34610 10824 35430
rect 10980 35086 11008 35566
rect 11808 35290 11836 35634
rect 11796 35284 11848 35290
rect 11796 35226 11848 35232
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 12268 34610 12296 35770
rect 10600 34604 10652 34610
rect 10600 34546 10652 34552
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 11152 34604 11204 34610
rect 11152 34546 11204 34552
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 10612 34406 10640 34546
rect 10600 34400 10652 34406
rect 10600 34342 10652 34348
rect 10508 34196 10560 34202
rect 10508 34138 10560 34144
rect 11164 33862 11192 34546
rect 11152 33856 11204 33862
rect 11152 33798 11204 33804
rect 10416 33108 10468 33114
rect 10416 33050 10468 33056
rect 10416 32972 10468 32978
rect 10416 32914 10468 32920
rect 10232 32904 10284 32910
rect 10232 32846 10284 32852
rect 10140 32768 10192 32774
rect 10140 32710 10192 32716
rect 10152 29306 10180 32710
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 10336 30258 10364 31078
rect 10324 30252 10376 30258
rect 10324 30194 10376 30200
rect 10428 29306 10456 32914
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10140 29300 10192 29306
rect 10140 29242 10192 29248
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 10152 29170 10180 29242
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 10048 28212 10100 28218
rect 10048 28154 10100 28160
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 25832 9916 25838
rect 9864 25774 9916 25780
rect 9680 24880 9732 24886
rect 9732 24840 9812 24868
rect 9680 24822 9732 24828
rect 9036 24686 9088 24692
rect 9048 24614 9076 24686
rect 9416 24670 9536 24698
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 8944 22568 8996 22574
rect 8944 22510 8996 22516
rect 9048 21894 9076 22578
rect 9232 22030 9260 22714
rect 9416 22094 9444 24670
rect 9588 24608 9640 24614
rect 9588 24550 9640 24556
rect 9600 24138 9628 24550
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9588 24132 9640 24138
rect 9588 24074 9640 24080
rect 9588 23724 9640 23730
rect 9588 23666 9640 23672
rect 9600 23526 9628 23666
rect 9496 23520 9548 23526
rect 9496 23462 9548 23468
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9508 23050 9536 23462
rect 9692 23118 9720 24142
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9416 22066 9536 22094
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9036 21888 9088 21894
rect 9036 21830 9088 21836
rect 9048 21486 9076 21830
rect 9036 21480 9088 21486
rect 9036 21422 9088 21428
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8956 17270 8984 19654
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 9508 16726 9536 22066
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9600 18290 9628 19382
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9600 16658 9628 18226
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 8864 15910 8892 16390
rect 9508 16182 9536 16390
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9692 16114 9720 16934
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 5778 8708 7686
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8300 4004 8352 4010
rect 8300 3946 8352 3952
rect 8312 3738 8340 3946
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8300 3732 8352 3738
rect 8300 3674 8352 3680
rect 8496 3670 8524 3878
rect 8484 3664 8536 3670
rect 8484 3606 8536 3612
rect 8680 3516 8708 5714
rect 8772 3602 8800 14758
rect 8864 5302 8892 15846
rect 8944 14340 8996 14346
rect 8944 14282 8996 14288
rect 8956 14006 8984 14282
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8956 13394 8984 13942
rect 8944 13388 8996 13394
rect 8944 13330 8996 13336
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9140 11762 9168 12310
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9232 9926 9260 15846
rect 9692 15416 9720 16050
rect 9784 15706 9812 24840
rect 9876 22094 9904 25774
rect 9968 25430 9996 26726
rect 9956 25424 10008 25430
rect 9956 25366 10008 25372
rect 9937 24812 9989 24818
rect 9989 24760 9996 24800
rect 9937 24754 9996 24760
rect 9968 23866 9996 24754
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 10060 22642 10088 28154
rect 10428 27674 10456 29242
rect 10520 28558 10548 29582
rect 10784 29572 10836 29578
rect 10784 29514 10836 29520
rect 10796 29306 10824 29514
rect 10784 29300 10836 29306
rect 10784 29242 10836 29248
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10796 28966 10824 29106
rect 10784 28960 10836 28966
rect 10784 28902 10836 28908
rect 10796 28762 10824 28902
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10796 28218 10824 28698
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10416 27668 10468 27674
rect 10416 27610 10468 27616
rect 10600 27532 10652 27538
rect 10600 27474 10652 27480
rect 10612 26926 10640 27474
rect 10692 27464 10744 27470
rect 10692 27406 10744 27412
rect 10600 26920 10652 26926
rect 10600 26862 10652 26868
rect 10612 26246 10640 26862
rect 10600 26240 10652 26246
rect 10600 26182 10652 26188
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10232 24064 10284 24070
rect 10232 24006 10284 24012
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 9876 22066 9996 22094
rect 9862 19816 9918 19825
rect 9862 19751 9864 19760
rect 9916 19751 9918 19760
rect 9864 19722 9916 19728
rect 9968 16794 9996 22066
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10060 21690 10088 21898
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10060 21554 10088 21626
rect 10152 21622 10180 22918
rect 10244 21894 10272 24006
rect 10336 23730 10364 24754
rect 10612 24206 10640 26182
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 10140 21616 10192 21622
rect 10140 21558 10192 21564
rect 10336 21554 10364 21966
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10428 18970 10456 19314
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 10046 15600 10102 15609
rect 10046 15535 10048 15544
rect 10100 15535 10102 15544
rect 10048 15506 10100 15512
rect 9692 15388 9996 15416
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9416 10441 9444 12922
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9600 12170 9628 12650
rect 9588 12164 9640 12170
rect 9588 12106 9640 12112
rect 9692 12102 9720 12854
rect 9784 12238 9812 12854
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9680 12096 9732 12102
rect 9680 12038 9732 12044
rect 9692 11121 9720 12038
rect 9876 11898 9904 12650
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9678 11112 9734 11121
rect 9678 11047 9734 11056
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9772 10464 9824 10470
rect 9402 10432 9458 10441
rect 9772 10406 9824 10412
rect 9402 10367 9458 10376
rect 9416 10033 9444 10367
rect 9784 10062 9812 10406
rect 9772 10056 9824 10062
rect 9402 10024 9458 10033
rect 9772 9998 9824 10004
rect 9402 9959 9458 9968
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9416 9382 9444 9862
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9404 9376 9456 9382
rect 9404 9318 9456 9324
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 6866 9260 7142
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 9312 6792 9364 6798
rect 8956 6740 9312 6746
rect 8956 6734 9364 6740
rect 8956 6718 9352 6734
rect 8956 6662 8984 6718
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 9036 6112 9088 6118
rect 9088 6060 9168 6066
rect 9036 6054 9168 6060
rect 9048 6038 9168 6054
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8956 5574 8984 5646
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 9048 5234 9076 5510
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8850 4448 8906 4457
rect 8850 4383 8906 4392
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8404 3488 8708 3516
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8220 800 8248 2994
rect 8300 2100 8352 2106
rect 8300 2042 8352 2048
rect 8312 800 8340 2042
rect 8404 800 8432 3488
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8576 3392 8628 3398
rect 8864 3346 8892 4383
rect 9048 3942 9076 5170
rect 9140 4622 9168 6038
rect 9416 4826 9444 9318
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9600 8129 9628 8570
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9692 7546 9720 8570
rect 9784 8498 9812 9658
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9784 7478 9812 8434
rect 9876 7546 9904 11018
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6322 9720 6598
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9784 5302 9812 7414
rect 9876 6934 9904 7482
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9772 5296 9824 5302
rect 9586 5264 9642 5273
rect 9508 5222 9586 5250
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9416 4049 9444 4218
rect 9402 4040 9458 4049
rect 9402 3975 9458 3984
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9310 3904 9366 3913
rect 8576 3334 8628 3340
rect 8496 3058 8524 3334
rect 8588 3194 8616 3334
rect 8680 3318 8892 3346
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8482 2272 8538 2281
rect 8482 2207 8538 2216
rect 8496 800 8524 2207
rect 8588 800 8616 2586
rect 8680 2378 8708 3318
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8772 800 8800 2994
rect 8864 800 8892 3130
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 9048 800 9076 2314
rect 9140 800 9168 3878
rect 9310 3839 9366 3848
rect 9324 3738 9352 3839
rect 9312 3732 9364 3738
rect 9312 3674 9364 3680
rect 9220 3528 9272 3534
rect 9218 3496 9220 3505
rect 9272 3496 9274 3505
rect 9274 3454 9352 3482
rect 9218 3431 9274 3440
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9232 2281 9260 2314
rect 9218 2272 9274 2281
rect 9218 2207 9274 2216
rect 9324 800 9352 3454
rect 9416 3398 9444 3975
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 9416 800 9444 2858
rect 9508 2854 9536 5222
rect 9772 5238 9824 5244
rect 9586 5199 9642 5208
rect 9784 4826 9812 5238
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9600 800 9628 3470
rect 9692 2854 9720 3975
rect 9770 3768 9826 3777
rect 9770 3703 9772 3712
rect 9824 3703 9826 3712
rect 9772 3674 9824 3680
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9876 2774 9904 4694
rect 9968 4146 9996 15388
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10244 14822 10272 14962
rect 10336 14958 10364 16662
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10520 15473 10548 16050
rect 10612 15638 10640 21286
rect 10704 16250 10732 27406
rect 10888 25838 10916 32846
rect 11164 31754 11192 33798
rect 11888 32496 11940 32502
rect 11888 32438 11940 32444
rect 11900 31958 11928 32438
rect 12072 32292 12124 32298
rect 12072 32234 12124 32240
rect 11888 31952 11940 31958
rect 11888 31894 11940 31900
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11072 31726 11192 31754
rect 10968 31680 11020 31686
rect 10968 31622 11020 31628
rect 10980 31346 11008 31622
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10968 30252 11020 30258
rect 10968 30194 11020 30200
rect 10980 27062 11008 30194
rect 11072 30190 11100 31726
rect 11532 30938 11560 31758
rect 11900 31414 11928 31894
rect 12084 31754 12112 32234
rect 12360 31754 12388 37130
rect 12440 36168 12492 36174
rect 12440 36110 12492 36116
rect 12452 35018 12480 36110
rect 12440 35012 12492 35018
rect 12440 34954 12492 34960
rect 12452 34610 12480 34954
rect 12440 34604 12492 34610
rect 12440 34546 12492 34552
rect 11992 31726 12112 31754
rect 12348 31748 12400 31754
rect 11888 31408 11940 31414
rect 11888 31350 11940 31356
rect 11992 31278 12020 31726
rect 12348 31690 12400 31696
rect 11980 31272 12032 31278
rect 11980 31214 12032 31220
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 11072 29510 11100 30126
rect 11060 29504 11112 29510
rect 11060 29446 11112 29452
rect 11072 27878 11100 29446
rect 11060 27872 11112 27878
rect 11060 27814 11112 27820
rect 10968 27056 11020 27062
rect 10968 26998 11020 27004
rect 10876 25832 10928 25838
rect 10876 25774 10928 25780
rect 10888 25294 10916 25774
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 10796 24410 10824 24686
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 10784 23724 10836 23730
rect 10784 23666 10836 23672
rect 10796 22982 10824 23666
rect 11072 23610 11100 27814
rect 11532 27130 11560 30874
rect 11992 30326 12020 31214
rect 12452 31142 12480 34546
rect 12544 32434 12572 38354
rect 12716 36848 12768 36854
rect 12716 36790 12768 36796
rect 12624 36576 12676 36582
rect 12624 36518 12676 36524
rect 12636 36122 12664 36518
rect 12728 36242 12756 36790
rect 12808 36780 12860 36786
rect 12808 36722 12860 36728
rect 12716 36236 12768 36242
rect 12716 36178 12768 36184
rect 12636 36094 12756 36122
rect 12624 35556 12676 35562
rect 12624 35498 12676 35504
rect 12636 34746 12664 35498
rect 12624 34740 12676 34746
rect 12624 34682 12676 34688
rect 12622 34640 12678 34649
rect 12622 34575 12678 34584
rect 12636 33658 12664 34575
rect 12624 33652 12676 33658
rect 12624 33594 12676 33600
rect 12728 33046 12756 36094
rect 12820 34950 12848 36722
rect 12808 34944 12860 34950
rect 12808 34886 12860 34892
rect 12820 34610 12848 34886
rect 12912 34678 12940 40122
rect 13188 35698 13216 40394
rect 13544 40180 13596 40186
rect 13544 40122 13596 40128
rect 13268 39432 13320 39438
rect 13268 39374 13320 39380
rect 13280 37126 13308 39374
rect 13360 37936 13412 37942
rect 13360 37878 13412 37884
rect 13268 37120 13320 37126
rect 13268 37062 13320 37068
rect 13280 36718 13308 37062
rect 13372 36854 13400 37878
rect 13360 36848 13412 36854
rect 13360 36790 13412 36796
rect 13268 36712 13320 36718
rect 13268 36654 13320 36660
rect 13280 36106 13308 36654
rect 13268 36100 13320 36106
rect 13268 36042 13320 36048
rect 13176 35692 13228 35698
rect 13176 35634 13228 35640
rect 12900 34672 12952 34678
rect 12900 34614 12952 34620
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 12716 33040 12768 33046
rect 12716 32982 12768 32988
rect 12728 32910 12756 32982
rect 12716 32904 12768 32910
rect 12716 32846 12768 32852
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 12820 31754 12848 34546
rect 13188 33153 13216 35634
rect 13280 33522 13308 36042
rect 13556 35154 13584 40122
rect 13832 38758 13860 41482
rect 14556 41472 14608 41478
rect 14556 41414 14608 41420
rect 14476 41386 14596 41414
rect 14280 40656 14332 40662
rect 14280 40598 14332 40604
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13636 38276 13688 38282
rect 13636 38218 13688 38224
rect 13648 37738 13676 38218
rect 13728 38208 13780 38214
rect 13728 38150 13780 38156
rect 13740 37942 13768 38150
rect 13728 37936 13780 37942
rect 13728 37878 13780 37884
rect 13636 37732 13688 37738
rect 13636 37674 13688 37680
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 13740 37126 13768 37606
rect 13728 37120 13780 37126
rect 13728 37062 13780 37068
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 14108 36378 14136 36722
rect 14096 36372 14148 36378
rect 14096 36314 14148 36320
rect 14292 36174 14320 40598
rect 14476 40526 14504 41386
rect 14648 41200 14700 41206
rect 14648 41142 14700 41148
rect 14660 40730 14688 41142
rect 14752 41138 14780 41550
rect 14740 41132 14792 41138
rect 14740 41074 14792 41080
rect 14752 41002 15056 41018
rect 14740 40996 15068 41002
rect 14792 40990 15016 40996
rect 14740 40938 14792 40944
rect 15016 40938 15068 40944
rect 14648 40724 14700 40730
rect 14648 40666 14700 40672
rect 14464 40520 14516 40526
rect 14464 40462 14516 40468
rect 14740 40452 14792 40458
rect 14740 40394 14792 40400
rect 14752 40186 14780 40394
rect 14740 40180 14792 40186
rect 14740 40122 14792 40128
rect 14648 37324 14700 37330
rect 14648 37266 14700 37272
rect 14372 37188 14424 37194
rect 14372 37130 14424 37136
rect 14556 37188 14608 37194
rect 14556 37130 14608 37136
rect 14384 36922 14412 37130
rect 14372 36916 14424 36922
rect 14372 36858 14424 36864
rect 14568 36650 14596 37130
rect 14556 36644 14608 36650
rect 14556 36586 14608 36592
rect 14660 36174 14688 37266
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14648 36168 14700 36174
rect 14648 36110 14700 36116
rect 14740 36168 14792 36174
rect 14740 36110 14792 36116
rect 13728 35828 13780 35834
rect 13728 35770 13780 35776
rect 13544 35148 13596 35154
rect 13544 35090 13596 35096
rect 13636 33992 13688 33998
rect 13636 33934 13688 33940
rect 13648 33658 13676 33934
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13174 33144 13230 33153
rect 13556 33114 13584 33458
rect 13174 33079 13230 33088
rect 13544 33108 13596 33114
rect 13544 33050 13596 33056
rect 13084 32904 13136 32910
rect 13084 32846 13136 32852
rect 12900 32768 12952 32774
rect 12900 32710 12952 32716
rect 12636 31726 12848 31754
rect 12636 31346 12664 31726
rect 12912 31414 12940 32710
rect 13096 32570 13124 32846
rect 13084 32564 13136 32570
rect 13084 32506 13136 32512
rect 13268 32428 13320 32434
rect 13268 32370 13320 32376
rect 12992 31748 13044 31754
rect 12992 31690 13044 31696
rect 13004 31482 13032 31690
rect 12992 31476 13044 31482
rect 12992 31418 13044 31424
rect 12900 31408 12952 31414
rect 12900 31350 12952 31356
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 11704 30320 11756 30326
rect 11704 30262 11756 30268
rect 11980 30320 12032 30326
rect 11980 30262 12032 30268
rect 11716 30054 11744 30262
rect 11704 30048 11756 30054
rect 11704 29990 11756 29996
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11716 29238 11744 29446
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11992 29170 12020 30262
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11900 28082 11928 28358
rect 12452 28218 12480 31078
rect 12532 28688 12584 28694
rect 12532 28630 12584 28636
rect 12440 28212 12492 28218
rect 12440 28154 12492 28160
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 11520 27124 11572 27130
rect 11520 27066 11572 27072
rect 11532 26382 11560 27066
rect 11716 26586 11744 28018
rect 12452 27334 12480 28154
rect 12544 28082 12572 28630
rect 12636 28082 12664 31282
rect 12912 30054 12940 31350
rect 12992 31272 13044 31278
rect 12992 31214 13044 31220
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 13004 29850 13032 31214
rect 13176 30048 13228 30054
rect 13176 29990 13228 29996
rect 12992 29844 13044 29850
rect 12992 29786 13044 29792
rect 13004 28694 13032 29786
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 12992 28688 13044 28694
rect 12992 28630 13044 28636
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12532 28076 12584 28082
rect 12532 28018 12584 28024
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12440 27328 12492 27334
rect 12440 27270 12492 27276
rect 12636 26994 12664 28018
rect 12912 27470 12940 28358
rect 13096 28218 13124 28698
rect 13084 28212 13136 28218
rect 13084 28154 13136 28160
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11704 26580 11756 26586
rect 11704 26522 11756 26528
rect 11520 26376 11572 26382
rect 11520 26318 11572 26324
rect 11428 25152 11480 25158
rect 11428 25094 11480 25100
rect 11440 24954 11468 25094
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11152 24132 11204 24138
rect 11152 24074 11204 24080
rect 11336 24132 11388 24138
rect 11336 24074 11388 24080
rect 11164 23798 11192 24074
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11152 23792 11204 23798
rect 11152 23734 11204 23740
rect 11072 23582 11192 23610
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10796 19378 10824 19450
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10796 16114 10824 19314
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10888 18766 10916 19110
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10704 15570 10732 16050
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10784 15496 10836 15502
rect 10506 15464 10562 15473
rect 10506 15399 10562 15408
rect 10782 15464 10784 15473
rect 10836 15464 10838 15473
rect 10782 15399 10838 15408
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10416 14884 10468 14890
rect 10416 14826 10468 14832
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10244 14278 10272 14758
rect 10428 14550 10456 14826
rect 10416 14544 10468 14550
rect 10416 14486 10468 14492
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10060 12850 10088 13262
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 10060 12714 10088 12786
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10244 9722 10272 14214
rect 10888 12986 10916 17002
rect 10980 16114 11008 21830
rect 11072 21418 11100 22714
rect 11060 21412 11112 21418
rect 11060 21354 11112 21360
rect 11164 21078 11192 23582
rect 11256 23118 11284 24006
rect 11348 23866 11376 24074
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11532 23118 11560 26318
rect 11992 26314 12020 26862
rect 11980 26308 12032 26314
rect 11980 26250 12032 26256
rect 12440 26308 12492 26314
rect 12440 26250 12492 26256
rect 11796 25356 11848 25362
rect 11796 25298 11848 25304
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11624 24206 11652 24550
rect 11612 24200 11664 24206
rect 11612 24142 11664 24148
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11520 23112 11572 23118
rect 11520 23054 11572 23060
rect 11624 22094 11652 24142
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11716 22982 11744 23598
rect 11808 23594 11836 25298
rect 11796 23588 11848 23594
rect 11796 23530 11848 23536
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11532 22066 11652 22094
rect 11152 21072 11204 21078
rect 11152 21014 11204 21020
rect 11164 20058 11192 21014
rect 11532 20534 11560 22066
rect 11716 22030 11744 22918
rect 11900 22438 11928 22986
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 22166 11928 22374
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11704 22024 11756 22030
rect 11704 21966 11756 21972
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 11624 21690 11652 21898
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11164 19242 11192 19994
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11164 18766 11192 19178
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 11532 18358 11560 18566
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11072 17542 11100 18226
rect 11624 18204 11652 20742
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11532 18176 11652 18204
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11072 14074 11100 17478
rect 11164 15502 11192 18022
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 16454 11284 16594
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10612 10577 10640 10610
rect 10692 10600 10744 10606
rect 10598 10568 10654 10577
rect 10692 10542 10744 10548
rect 10598 10503 10654 10512
rect 10704 10130 10732 10542
rect 11072 10266 11100 14010
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12434 11468 13262
rect 11348 12406 11468 12434
rect 11348 11694 11376 12406
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11348 11150 11376 11630
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10692 10124 10744 10130
rect 10692 10066 10744 10072
rect 10704 9722 10732 10066
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 11348 7342 11376 11086
rect 11440 9654 11468 12174
rect 11532 11370 11560 18176
rect 11808 18154 11836 18702
rect 11796 18148 11848 18154
rect 11796 18090 11848 18096
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11808 15502 11836 17478
rect 11900 17338 11928 17478
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11992 16250 12020 26250
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12360 25906 12388 26182
rect 12452 26042 12480 26250
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12360 25294 12388 25842
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12268 23866 12296 24142
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12176 21962 12204 22578
rect 12164 21956 12216 21962
rect 12164 21898 12216 21904
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 11980 16244 12032 16250
rect 11980 16186 12032 16192
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 12084 15026 12112 21830
rect 12256 21072 12308 21078
rect 12256 21014 12308 21020
rect 12268 19854 12296 21014
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12176 18766 12204 19178
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12268 18086 12296 18702
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 12360 17762 12388 25230
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 12912 24206 12940 24550
rect 12992 24404 13044 24410
rect 12992 24346 13044 24352
rect 12900 24200 12952 24206
rect 12898 24168 12900 24177
rect 12952 24168 12954 24177
rect 12898 24103 12954 24112
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12452 23526 12480 23802
rect 13004 23798 13032 24346
rect 12992 23792 13044 23798
rect 12992 23734 13044 23740
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12440 22024 12492 22030
rect 12440 21966 12492 21972
rect 12452 21554 12480 21966
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12544 20602 12572 23462
rect 13188 21876 13216 29990
rect 13280 28082 13308 32370
rect 13452 32360 13504 32366
rect 13452 32302 13504 32308
rect 13464 32026 13492 32302
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13452 32020 13504 32026
rect 13452 31962 13504 31968
rect 13360 31680 13412 31686
rect 13360 31622 13412 31628
rect 13372 31346 13400 31622
rect 13648 31346 13676 32166
rect 13740 31346 13768 35770
rect 14752 35562 14780 36110
rect 14740 35556 14792 35562
rect 14740 35498 14792 35504
rect 13820 33992 13872 33998
rect 13820 33934 13872 33940
rect 13832 32978 13860 33934
rect 14464 33584 14516 33590
rect 14462 33552 14464 33561
rect 14516 33552 14518 33561
rect 14462 33487 14518 33496
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 14648 33312 14700 33318
rect 14648 33254 14700 33260
rect 13820 32972 13872 32978
rect 13820 32914 13872 32920
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 14108 32434 14136 32846
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 13636 31340 13688 31346
rect 13636 31282 13688 31288
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13740 30870 13768 31282
rect 14384 31278 14412 33254
rect 14660 32502 14688 33254
rect 14740 32904 14792 32910
rect 14740 32846 14792 32852
rect 14648 32496 14700 32502
rect 14648 32438 14700 32444
rect 14660 31346 14688 32438
rect 14752 31822 14780 32846
rect 14740 31816 14792 31822
rect 14740 31758 14792 31764
rect 14648 31340 14700 31346
rect 14648 31282 14700 31288
rect 14372 31272 14424 31278
rect 14372 31214 14424 31220
rect 13728 30864 13780 30870
rect 13728 30806 13780 30812
rect 13740 29306 13768 30806
rect 14752 30802 14780 31758
rect 15016 31680 15068 31686
rect 15016 31622 15068 31628
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 14740 30796 14792 30802
rect 14740 30738 14792 30744
rect 14740 30660 14792 30666
rect 14740 30602 14792 30608
rect 14752 30394 14780 30602
rect 14740 30388 14792 30394
rect 14740 30330 14792 30336
rect 14648 30320 14700 30326
rect 14648 30262 14700 30268
rect 13728 29300 13780 29306
rect 13728 29242 13780 29248
rect 13636 28960 13688 28966
rect 13636 28902 13688 28908
rect 13360 28552 13412 28558
rect 13360 28494 13412 28500
rect 13372 28218 13400 28494
rect 13648 28422 13676 28902
rect 13740 28558 13768 29242
rect 14188 29232 14240 29238
rect 14188 29174 14240 29180
rect 14200 28558 14228 29174
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 14188 28552 14240 28558
rect 14188 28494 14240 28500
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 13636 28416 13688 28422
rect 13636 28358 13688 28364
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 13268 28076 13320 28082
rect 13268 28018 13320 28024
rect 13280 27878 13308 28018
rect 13268 27872 13320 27878
rect 13268 27814 13320 27820
rect 13464 27674 13492 28086
rect 13648 28014 13676 28358
rect 13636 28008 13688 28014
rect 13636 27950 13688 27956
rect 13452 27668 13504 27674
rect 13452 27610 13504 27616
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13280 25158 13308 25842
rect 13268 25152 13320 25158
rect 13268 25094 13320 25100
rect 13280 22710 13308 25094
rect 13268 22704 13320 22710
rect 13268 22646 13320 22652
rect 13372 22030 13400 26862
rect 13648 26042 13676 27950
rect 14568 26518 14596 28494
rect 14660 28150 14688 30262
rect 14844 30258 14872 31282
rect 15028 30258 15056 31622
rect 14832 30252 14884 30258
rect 14832 30194 14884 30200
rect 15016 30252 15068 30258
rect 15016 30194 15068 30200
rect 14844 28490 14872 30194
rect 15028 30054 15056 30194
rect 15016 30048 15068 30054
rect 14936 30008 15016 30036
rect 14832 28484 14884 28490
rect 14832 28426 14884 28432
rect 14648 28144 14700 28150
rect 14648 28086 14700 28092
rect 14556 26512 14608 26518
rect 14556 26454 14608 26460
rect 13636 26036 13688 26042
rect 13636 25978 13688 25984
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13636 24676 13688 24682
rect 13636 24618 13688 24624
rect 13648 24206 13676 24618
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 23730 13492 24006
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13556 23526 13584 24142
rect 13740 24138 13768 25774
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 14108 24410 14136 24754
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 14200 23798 14228 24550
rect 14660 24206 14688 25094
rect 14936 24410 14964 30008
rect 15016 29990 15068 29996
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 15028 25226 15056 25638
rect 15016 25220 15068 25226
rect 15016 25162 15068 25168
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 15028 24342 15056 25162
rect 15016 24336 15068 24342
rect 15016 24278 15068 24284
rect 14648 24200 14700 24206
rect 14832 24200 14884 24206
rect 14648 24142 14700 24148
rect 14830 24168 14832 24177
rect 14884 24168 14886 24177
rect 14830 24103 14886 24112
rect 14924 24132 14976 24138
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 14844 23662 14872 24103
rect 14924 24074 14976 24080
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14936 23594 14964 24074
rect 14464 23588 14516 23594
rect 14464 23530 14516 23536
rect 14924 23588 14976 23594
rect 14924 23530 14976 23536
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 14372 23044 14424 23050
rect 14372 22986 14424 22992
rect 14384 22642 14412 22986
rect 14476 22710 14504 23530
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13544 21888 13596 21894
rect 13188 21848 13544 21876
rect 13544 21830 13596 21836
rect 13556 21486 13584 21830
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12716 20868 12768 20874
rect 12716 20810 12768 20816
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 12440 20256 12492 20262
rect 12440 20198 12492 20204
rect 12452 19446 12480 20198
rect 12544 20058 12572 20402
rect 12532 20052 12584 20058
rect 12532 19994 12584 20000
rect 12728 19718 12756 20810
rect 12992 20800 13044 20806
rect 12992 20742 13044 20748
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12820 19990 12848 20402
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12544 19310 12572 19654
rect 12728 19378 12756 19654
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12728 18698 12756 19314
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12728 18222 12756 18634
rect 12820 18630 12848 19926
rect 13004 19854 13032 20742
rect 13096 19854 13124 21082
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13648 20602 13676 20946
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 14096 20392 14148 20398
rect 14096 20334 14148 20340
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12716 18216 12768 18222
rect 12716 18158 12768 18164
rect 12268 17734 12388 17762
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12176 16114 12204 16390
rect 12164 16108 12216 16114
rect 12164 16050 12216 16056
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11624 12238 11652 12582
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11716 12102 11744 12786
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11808 11762 11836 14350
rect 12072 13796 12124 13802
rect 12072 13738 12124 13744
rect 12084 12850 12112 13738
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11888 12776 11940 12782
rect 11888 12718 11940 12724
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11532 11342 11652 11370
rect 11624 11286 11652 11342
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 11428 9648 11480 9654
rect 11428 9590 11480 9596
rect 11440 9110 11468 9590
rect 11428 9104 11480 9110
rect 11428 9046 11480 9052
rect 11440 7886 11468 9046
rect 11520 8288 11572 8294
rect 11520 8230 11572 8236
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11336 7336 11388 7342
rect 11336 7278 11388 7284
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10152 3942 10180 4694
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3602 10180 3878
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 9876 2746 9996 2774
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9692 800 9720 2518
rect 9968 800 9996 2746
rect 10048 2304 10100 2310
rect 10048 2246 10100 2252
rect 10060 2038 10088 2246
rect 10048 2032 10100 2038
rect 10048 1974 10100 1980
rect 10244 800 10272 4966
rect 10336 3534 10364 7142
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6118 11100 6734
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6458 11284 6598
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11440 6390 11468 7822
rect 11532 7818 11560 8230
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11624 7410 11652 11222
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9586 11744 9862
rect 11808 9586 11836 9930
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11900 8906 11928 12718
rect 11992 10198 12020 12718
rect 12176 12434 12204 16050
rect 12268 13530 12296 17734
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12360 17338 12388 17614
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12728 17202 12756 18158
rect 12820 17746 12848 18566
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12268 13297 12296 13466
rect 12254 13288 12310 13297
rect 12254 13223 12310 13232
rect 12084 12406 12204 12434
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11980 9512 12032 9518
rect 11980 9454 12032 9460
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 11900 8498 11928 8842
rect 11992 8838 12020 9454
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11612 7404 11664 7410
rect 11612 7346 11664 7352
rect 11716 6662 11744 7822
rect 11808 7750 11836 8434
rect 11900 7954 11928 8434
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10428 4078 10456 4626
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10428 3602 10456 4014
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10428 2990 10456 3538
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10414 2408 10470 2417
rect 10414 2343 10470 2352
rect 10428 2310 10456 2343
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10428 1902 10456 2246
rect 10416 1896 10468 1902
rect 10416 1838 10468 1844
rect 10520 800 10548 5646
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10600 4548 10652 4554
rect 10600 4490 10652 4496
rect 10612 4010 10640 4490
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10612 3534 10640 3946
rect 10704 3602 10732 3946
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10690 3360 10746 3369
rect 10690 3295 10746 3304
rect 10704 3058 10732 3295
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 10796 800 10824 4966
rect 10888 4554 10916 5578
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10980 4078 11008 4558
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10980 3670 11008 4014
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 11072 800 11100 5646
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 800 11376 4966
rect 11440 2774 11468 6054
rect 11532 4146 11560 6598
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11440 2746 11560 2774
rect 11532 2446 11560 2746
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11624 800 11652 5646
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11716 3534 11744 4082
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11808 3058 11836 7686
rect 11886 7576 11942 7585
rect 11886 7511 11888 7520
rect 11940 7511 11942 7520
rect 11888 7482 11940 7488
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11900 800 11928 4966
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11992 3602 12020 3878
rect 12084 3738 12112 12406
rect 12360 12170 12388 16118
rect 12544 16046 12572 16118
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12544 14074 12572 14826
rect 12636 14822 12664 15370
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12728 14890 12756 15098
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12820 14618 12848 14962
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 12912 14278 12940 18702
rect 12992 17672 13044 17678
rect 13096 17660 13124 19790
rect 14108 19514 14136 20334
rect 14200 19786 14228 22510
rect 14384 21690 14412 22578
rect 14844 22506 14872 23054
rect 14924 22976 14976 22982
rect 14924 22918 14976 22924
rect 14936 22574 14964 22918
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14464 21616 14516 21622
rect 14464 21558 14516 21564
rect 14476 20942 14504 21558
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14188 19780 14240 19786
rect 14188 19722 14240 19728
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13188 18086 13216 19382
rect 14200 19378 14228 19722
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 13728 19304 13780 19310
rect 13728 19246 13780 19252
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13176 18080 13228 18086
rect 13176 18022 13228 18028
rect 13188 17814 13216 18022
rect 13268 17876 13320 17882
rect 13268 17818 13320 17824
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13044 17632 13124 17660
rect 12992 17614 13044 17620
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 13096 15638 13124 17206
rect 13188 15706 13216 17750
rect 13280 17678 13308 17818
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 17338 13308 17614
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 12990 15464 13046 15473
rect 12990 15399 13046 15408
rect 13004 15026 13032 15399
rect 13096 15094 13124 15574
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12176 9722 12204 9930
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 7818 12204 8774
rect 12268 8362 12296 11494
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12544 9042 12572 9998
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12544 8922 12572 8978
rect 12452 8894 12572 8922
rect 12452 8650 12480 8894
rect 12360 8622 12480 8650
rect 12360 8566 12388 8622
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12256 8356 12308 8362
rect 12256 8298 12308 8304
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12452 7546 12480 8298
rect 12636 7750 12664 8434
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12544 6798 12572 7686
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12636 6730 12664 7686
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12624 6724 12676 6730
rect 12624 6666 12676 6672
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12072 3732 12124 3738
rect 12072 3674 12124 3680
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 12176 800 12204 4558
rect 12268 4146 12296 6666
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12452 800 12480 5646
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12636 1306 12664 2450
rect 12728 2446 12756 12038
rect 12808 10192 12860 10198
rect 12808 10134 12860 10140
rect 12820 9926 12848 10134
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 8974 13032 9862
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 13004 8634 13032 8910
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13096 8566 13124 9318
rect 13084 8560 13136 8566
rect 13084 8502 13136 8508
rect 12992 8356 13044 8362
rect 12992 8298 13044 8304
rect 12806 6352 12862 6361
rect 12806 6287 12862 6296
rect 12820 2774 12848 6287
rect 12900 6248 12952 6254
rect 13004 6202 13032 8298
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6390 13124 6734
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 12952 6196 13032 6202
rect 12900 6190 13032 6196
rect 12912 6174 13032 6190
rect 13004 6118 13032 6174
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12912 5846 12940 6054
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12820 2746 12940 2774
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12912 2038 12940 2746
rect 12900 2032 12952 2038
rect 12900 1974 12952 1980
rect 12636 1278 12756 1306
rect 12728 800 12756 1278
rect 13004 800 13032 4558
rect 13188 3942 13216 15438
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 8430 13308 10542
rect 13360 9580 13412 9586
rect 13360 9522 13412 9528
rect 13372 8634 13400 9522
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13464 7954 13492 18838
rect 13740 18358 13768 19246
rect 14200 18970 14228 19314
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 13728 18352 13780 18358
rect 13728 18294 13780 18300
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17746 13860 18022
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13924 17338 13952 18906
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14292 17202 14320 19314
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 17882 14412 18226
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14384 17202 14412 17818
rect 14568 17202 14596 22374
rect 14936 22234 14964 22510
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14016 14958 14044 17138
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14200 15638 14228 16050
rect 14292 15978 14320 17138
rect 14556 16516 14608 16522
rect 14556 16458 14608 16464
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14188 15632 14240 15638
rect 14188 15574 14240 15580
rect 14188 15428 14240 15434
rect 14292 15416 14320 15914
rect 14476 15706 14504 16050
rect 14568 15706 14596 16458
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14568 15502 14596 15642
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14240 15388 14320 15416
rect 14188 15370 14240 15376
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14004 14952 14056 14958
rect 14004 14894 14056 14900
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13924 12918 13952 13874
rect 14108 12918 14136 15302
rect 14568 15162 14596 15438
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14550 14412 14758
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14476 14006 14504 14554
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14844 13462 14872 21966
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14832 13456 14884 13462
rect 14832 13398 14884 13404
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 14096 12912 14148 12918
rect 14096 12854 14148 12860
rect 13924 12238 13952 12854
rect 14108 12442 14136 12854
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13740 11898 13768 12106
rect 14752 11898 14780 13262
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14844 11830 14872 12038
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14936 11082 14964 19654
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 15028 17610 15056 18770
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 15028 16114 15056 17070
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13394 15056 13670
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13556 9722 13584 10202
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13556 9178 13584 9658
rect 14752 9586 14780 10134
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14016 8634 14044 8978
rect 14476 8974 14504 9318
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13924 7750 13952 8434
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13556 6361 13584 7686
rect 14752 7206 14780 9522
rect 15028 9382 15056 11834
rect 15016 9376 15068 9382
rect 15016 9318 15068 9324
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 13542 6352 13598 6361
rect 13542 6287 13598 6296
rect 13740 6186 13952 6202
rect 13728 6180 13952 6186
rect 13780 6174 13952 6180
rect 13728 6122 13780 6128
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 13280 800 13308 5646
rect 13464 5166 13492 6054
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13464 2774 13492 4626
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13556 3466 13584 3878
rect 13544 3460 13596 3466
rect 13544 3402 13596 3408
rect 13728 3120 13780 3126
rect 13726 3088 13728 3097
rect 13780 3088 13782 3097
rect 13726 3023 13782 3032
rect 13464 2746 13584 2774
rect 13556 800 13584 2746
rect 13832 800 13860 4966
rect 13924 4622 13952 6174
rect 14292 5234 14320 7142
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14476 5914 14504 6258
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14660 5778 14688 6258
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14752 5710 14780 7142
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 13912 4616 13964 4622
rect 13912 4558 13964 4564
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 14016 3534 14044 4422
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 14004 3528 14056 3534
rect 14004 3470 14056 3476
rect 13924 2774 13952 3470
rect 13924 2746 14044 2774
rect 14016 1494 14044 2746
rect 14004 1488 14056 1494
rect 14004 1430 14056 1436
rect 14108 800 14136 4966
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14200 800 14228 4558
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14292 1426 14320 4082
rect 14462 4040 14518 4049
rect 14462 3975 14518 3984
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14280 1420 14332 1426
rect 14280 1362 14332 1368
rect 14384 800 14412 3538
rect 14476 3194 14504 3975
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14568 2774 14596 5170
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14476 2746 14596 2774
rect 14476 800 14504 2746
rect 14554 2680 14610 2689
rect 14554 2615 14610 2624
rect 14568 2582 14596 2615
rect 14556 2576 14608 2582
rect 14556 2518 14608 2524
rect 14660 800 14688 3674
rect 14752 3602 14780 4966
rect 14740 3596 14792 3602
rect 14740 3538 14792 3544
rect 14844 3466 14872 6394
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 3534 14964 6054
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 3058 14872 3402
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14936 3233 14964 3334
rect 14922 3224 14978 3233
rect 14922 3159 14978 3168
rect 15028 3058 15056 7210
rect 15120 3126 15148 55558
rect 15200 42220 15252 42226
rect 15200 42162 15252 42168
rect 15212 41818 15240 42162
rect 15568 42152 15620 42158
rect 15568 42094 15620 42100
rect 15200 41812 15252 41818
rect 15200 41754 15252 41760
rect 15580 41546 15608 42094
rect 15660 42016 15712 42022
rect 15660 41958 15712 41964
rect 15200 41540 15252 41546
rect 15200 41482 15252 41488
rect 15568 41540 15620 41546
rect 15568 41482 15620 41488
rect 15212 41414 15240 41482
rect 15212 41386 15516 41414
rect 15384 40928 15436 40934
rect 15384 40870 15436 40876
rect 15396 40118 15424 40870
rect 15384 40112 15436 40118
rect 15384 40054 15436 40060
rect 15488 39642 15516 41386
rect 15580 41070 15608 41482
rect 15568 41064 15620 41070
rect 15568 41006 15620 41012
rect 15476 39636 15528 39642
rect 15476 39578 15528 39584
rect 15488 38282 15516 39578
rect 15580 38962 15608 41006
rect 15672 40458 15700 41958
rect 16120 40520 16172 40526
rect 16120 40462 16172 40468
rect 15660 40452 15712 40458
rect 15660 40394 15712 40400
rect 16132 40050 16160 40462
rect 16120 40044 16172 40050
rect 16120 39986 16172 39992
rect 16132 39438 16160 39986
rect 16120 39432 16172 39438
rect 16120 39374 16172 39380
rect 15568 38956 15620 38962
rect 15568 38898 15620 38904
rect 16304 38820 16356 38826
rect 16304 38762 16356 38768
rect 15476 38276 15528 38282
rect 15476 38218 15528 38224
rect 15200 37188 15252 37194
rect 15200 37130 15252 37136
rect 15568 37188 15620 37194
rect 15568 37130 15620 37136
rect 15212 36718 15240 37130
rect 15580 36922 15608 37130
rect 16120 37120 16172 37126
rect 16120 37062 16172 37068
rect 15568 36916 15620 36922
rect 15568 36858 15620 36864
rect 16132 36786 16160 37062
rect 15752 36780 15804 36786
rect 15752 36722 15804 36728
rect 16120 36780 16172 36786
rect 16120 36722 16172 36728
rect 15200 36712 15252 36718
rect 15200 36654 15252 36660
rect 15212 36106 15240 36654
rect 15764 36378 15792 36722
rect 15752 36372 15804 36378
rect 15752 36314 15804 36320
rect 15200 36100 15252 36106
rect 15200 36042 15252 36048
rect 15212 35562 15240 36042
rect 16132 35766 16160 36722
rect 16316 36378 16344 38762
rect 16304 36372 16356 36378
rect 16304 36314 16356 36320
rect 16120 35760 16172 35766
rect 16120 35702 16172 35708
rect 15200 35556 15252 35562
rect 15200 35498 15252 35504
rect 15212 34066 15240 35498
rect 15936 34400 15988 34406
rect 15936 34342 15988 34348
rect 15200 34060 15252 34066
rect 15200 34002 15252 34008
rect 15948 33998 15976 34342
rect 15936 33992 15988 33998
rect 15936 33934 15988 33940
rect 15476 33924 15528 33930
rect 15476 33866 15528 33872
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15212 33386 15240 33458
rect 15200 33380 15252 33386
rect 15200 33322 15252 33328
rect 15212 31346 15240 33322
rect 15488 32978 15516 33866
rect 16132 33862 16160 35702
rect 15660 33856 15712 33862
rect 15660 33798 15712 33804
rect 16120 33856 16172 33862
rect 16120 33798 16172 33804
rect 15476 32972 15528 32978
rect 15476 32914 15528 32920
rect 15672 32842 15700 33798
rect 15660 32836 15712 32842
rect 15660 32778 15712 32784
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 16040 31414 16068 31962
rect 15844 31408 15896 31414
rect 15844 31350 15896 31356
rect 16028 31408 16080 31414
rect 16028 31350 16080 31356
rect 15200 31340 15252 31346
rect 15200 31282 15252 31288
rect 15212 30394 15240 31282
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15200 30388 15252 30394
rect 15200 30330 15252 30336
rect 15212 28558 15240 30330
rect 15304 30258 15332 31078
rect 15292 30252 15344 30258
rect 15292 30194 15344 30200
rect 15384 30252 15436 30258
rect 15384 30194 15436 30200
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15212 20058 15240 28358
rect 15396 28082 15424 30194
rect 15384 28076 15436 28082
rect 15384 28018 15436 28024
rect 15396 24886 15424 28018
rect 15384 24880 15436 24886
rect 15384 24822 15436 24828
rect 15384 23520 15436 23526
rect 15384 23462 15436 23468
rect 15292 22976 15344 22982
rect 15292 22918 15344 22924
rect 15304 20942 15332 22918
rect 15396 22030 15424 23462
rect 15384 22024 15436 22030
rect 15384 21966 15436 21972
rect 15384 21888 15436 21894
rect 15384 21830 15436 21836
rect 15396 21418 15424 21830
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15292 20936 15344 20942
rect 15292 20878 15344 20884
rect 15292 20460 15344 20466
rect 15292 20402 15344 20408
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15198 19952 15254 19961
rect 15198 19887 15200 19896
rect 15252 19887 15254 19896
rect 15200 19858 15252 19864
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15212 17202 15240 19450
rect 15304 17202 15332 20402
rect 15488 19174 15516 31146
rect 15856 30870 15884 31350
rect 15844 30864 15896 30870
rect 15844 30806 15896 30812
rect 15844 30184 15896 30190
rect 15844 30126 15896 30132
rect 15752 29572 15804 29578
rect 15752 29514 15804 29520
rect 15660 29164 15712 29170
rect 15660 29106 15712 29112
rect 15568 28960 15620 28966
rect 15568 28902 15620 28908
rect 15580 28082 15608 28902
rect 15672 28762 15700 29106
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15568 25152 15620 25158
rect 15568 25094 15620 25100
rect 15580 24614 15608 25094
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15580 23050 15608 24550
rect 15568 23044 15620 23050
rect 15568 22986 15620 22992
rect 15764 22522 15792 29514
rect 15856 22658 15884 30126
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15948 29782 15976 29990
rect 15936 29776 15988 29782
rect 15936 29718 15988 29724
rect 16028 28484 16080 28490
rect 16028 28426 16080 28432
rect 16040 28218 16068 28426
rect 16028 28212 16080 28218
rect 16028 28154 16080 28160
rect 16028 27532 16080 27538
rect 16028 27474 16080 27480
rect 16040 27130 16068 27474
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 16028 27124 16080 27130
rect 16028 27066 16080 27072
rect 16040 25906 16068 27066
rect 16224 26926 16252 27270
rect 16212 26920 16264 26926
rect 16212 26862 16264 26868
rect 16028 25900 16080 25906
rect 16028 25842 16080 25848
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15948 22778 15976 23054
rect 15936 22772 15988 22778
rect 15936 22714 15988 22720
rect 15856 22630 15976 22658
rect 15764 22494 15884 22522
rect 15752 22432 15804 22438
rect 15752 22374 15804 22380
rect 15764 22098 15792 22374
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15764 21706 15792 22034
rect 15856 21894 15884 22494
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15568 21684 15620 21690
rect 15764 21678 15884 21706
rect 15568 21626 15620 21632
rect 15580 20942 15608 21626
rect 15752 21548 15804 21554
rect 15752 21490 15804 21496
rect 15568 20936 15620 20942
rect 15568 20878 15620 20884
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15292 17196 15344 17202
rect 15292 17138 15344 17144
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15212 13530 15240 14282
rect 15580 13802 15608 18022
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15672 13326 15700 20810
rect 15764 20466 15792 21490
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15764 20058 15792 20402
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15856 14006 15884 21678
rect 15948 20398 15976 22630
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15948 19718 15976 20334
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15304 12782 15332 13126
rect 15396 12850 15424 13262
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15212 12238 15240 12582
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15488 11762 15516 12174
rect 15580 11898 15608 13194
rect 15672 12646 15700 13262
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15396 9518 15424 9862
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15212 6866 15240 9454
rect 15488 9330 15516 9862
rect 15304 9302 15516 9330
rect 15304 7886 15332 9302
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15488 8634 15516 9114
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15304 7478 15332 7822
rect 15384 7812 15436 7818
rect 15384 7754 15436 7760
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 15396 7002 15424 7754
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15580 6390 15608 7822
rect 15672 7546 15700 10746
rect 15764 9654 15792 12650
rect 15856 10266 15884 13942
rect 15948 10810 15976 19654
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16040 16998 16068 17274
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16028 15428 16080 15434
rect 16028 15370 16080 15376
rect 16040 15094 16068 15370
rect 16028 15088 16080 15094
rect 16028 15030 16080 15036
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 12306 16160 12718
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11558 16068 12174
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15304 5234 15332 5646
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5234 15516 5510
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 15016 3052 15068 3058
rect 15016 2994 15068 3000
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14752 2650 14780 2790
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14740 1420 14792 1426
rect 14740 1362 14792 1368
rect 14752 800 14780 1362
rect 14936 800 14964 2858
rect 15212 2836 15240 3946
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 15028 2808 15240 2836
rect 15028 2428 15056 2808
rect 15304 2774 15332 3402
rect 15120 2746 15332 2774
rect 15120 2666 15148 2746
rect 15120 2638 15332 2666
rect 15028 2400 15240 2428
rect 15016 1488 15068 1494
rect 15016 1430 15068 1436
rect 15028 800 15056 1430
rect 15212 800 15240 2400
rect 15304 800 15332 2638
rect 15396 800 15424 4558
rect 15580 4146 15608 6326
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5778 15792 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15474 3088 15530 3097
rect 15474 3023 15530 3032
rect 15568 3052 15620 3058
rect 15488 2378 15516 3023
rect 15568 2994 15620 3000
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 15488 1766 15516 2314
rect 15476 1760 15528 1766
rect 15476 1702 15528 1708
rect 15580 800 15608 2994
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 15672 800 15700 2926
rect 15764 1170 15792 3470
rect 15856 2650 15884 9998
rect 15948 9926 15976 10610
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 16040 9178 16068 11494
rect 16224 10606 16252 26862
rect 16304 25492 16356 25498
rect 16304 25434 16356 25440
rect 16316 24954 16344 25434
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16316 23526 16344 24142
rect 16304 23520 16356 23526
rect 16304 23462 16356 23468
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16316 16794 16344 18090
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16316 16590 16344 16730
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16316 14958 16344 15302
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16316 13870 16344 14894
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16408 12434 16436 55626
rect 16316 12406 16436 12434
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 16040 8294 16068 8434
rect 16028 8288 16080 8294
rect 16026 8256 16028 8265
rect 16080 8256 16082 8265
rect 16026 8191 16082 8200
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 5642 15976 6666
rect 16040 5778 16068 6734
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 16132 5642 16160 6258
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15948 5302 15976 5578
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 15936 3936 15988 3942
rect 15936 3878 15988 3884
rect 15948 3602 15976 3878
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 16040 2530 16068 4558
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 15948 2502 16068 2530
rect 15764 1142 15884 1170
rect 15856 800 15884 1142
rect 15948 800 15976 2502
rect 16026 2408 16082 2417
rect 16026 2343 16082 2352
rect 16040 2310 16068 2343
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16132 800 16160 2586
rect 16224 800 16252 4014
rect 16316 3126 16344 12406
rect 16500 4706 16528 56306
rect 16592 55622 16620 56306
rect 17236 55622 17264 56306
rect 17880 55962 17908 56306
rect 17868 55956 17920 55962
rect 17868 55898 17920 55904
rect 16580 55616 16632 55622
rect 16578 55584 16580 55593
rect 17224 55616 17276 55622
rect 16632 55584 16634 55593
rect 16578 55519 16634 55528
rect 17222 55584 17224 55593
rect 17276 55584 17278 55593
rect 17222 55519 17278 55528
rect 16948 42764 17000 42770
rect 16948 42706 17000 42712
rect 16580 41676 16632 41682
rect 16580 41618 16632 41624
rect 16592 39370 16620 41618
rect 16764 41540 16816 41546
rect 16764 41482 16816 41488
rect 16776 40390 16804 41482
rect 16764 40384 16816 40390
rect 16764 40326 16816 40332
rect 16580 39364 16632 39370
rect 16580 39306 16632 39312
rect 16776 37942 16804 40326
rect 16764 37936 16816 37942
rect 16764 37878 16816 37884
rect 16856 37392 16908 37398
rect 16856 37334 16908 37340
rect 16868 36854 16896 37334
rect 16856 36848 16908 36854
rect 16856 36790 16908 36796
rect 16672 34740 16724 34746
rect 16672 34682 16724 34688
rect 16580 33992 16632 33998
rect 16580 33934 16632 33940
rect 16592 33114 16620 33934
rect 16684 33522 16712 34682
rect 16856 33924 16908 33930
rect 16856 33866 16908 33872
rect 16868 33522 16896 33866
rect 16672 33516 16724 33522
rect 16672 33458 16724 33464
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16868 33114 16896 33458
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16856 33108 16908 33114
rect 16856 33050 16908 33056
rect 16672 32972 16724 32978
rect 16672 32914 16724 32920
rect 16684 30258 16712 32914
rect 16856 32428 16908 32434
rect 16856 32370 16908 32376
rect 16868 30326 16896 32370
rect 16960 31754 16988 42706
rect 17224 42560 17276 42566
rect 17224 42502 17276 42508
rect 17236 42226 17264 42502
rect 17224 42220 17276 42226
rect 17224 42162 17276 42168
rect 17236 41614 17264 42162
rect 17224 41608 17276 41614
rect 17224 41550 17276 41556
rect 17776 41200 17828 41206
rect 17776 41142 17828 41148
rect 17408 40112 17460 40118
rect 17408 40054 17460 40060
rect 17420 39846 17448 40054
rect 17408 39840 17460 39846
rect 17408 39782 17460 39788
rect 17420 37466 17448 39782
rect 17592 38344 17644 38350
rect 17592 38286 17644 38292
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 17604 38010 17632 38286
rect 17592 38004 17644 38010
rect 17592 37946 17644 37952
rect 17408 37460 17460 37466
rect 17408 37402 17460 37408
rect 17696 37398 17724 38286
rect 17788 38010 17816 41142
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 17776 37664 17828 37670
rect 17776 37606 17828 37612
rect 17684 37392 17736 37398
rect 17684 37334 17736 37340
rect 17408 37256 17460 37262
rect 17408 37198 17460 37204
rect 17592 37256 17644 37262
rect 17592 37198 17644 37204
rect 17420 37126 17448 37198
rect 17408 37120 17460 37126
rect 17408 37062 17460 37068
rect 17604 36922 17632 37198
rect 17592 36916 17644 36922
rect 17592 36858 17644 36864
rect 17788 36854 17816 37606
rect 17776 36848 17828 36854
rect 17776 36790 17828 36796
rect 17684 36780 17736 36786
rect 17684 36722 17736 36728
rect 17132 35692 17184 35698
rect 17132 35634 17184 35640
rect 17408 35692 17460 35698
rect 17408 35634 17460 35640
rect 17144 35562 17172 35634
rect 17132 35556 17184 35562
rect 17132 35498 17184 35504
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17236 35086 17264 35430
rect 17316 35284 17368 35290
rect 17316 35226 17368 35232
rect 17132 35080 17184 35086
rect 17132 35022 17184 35028
rect 17224 35080 17276 35086
rect 17224 35022 17276 35028
rect 17144 32910 17172 35022
rect 17328 34932 17356 35226
rect 17236 34904 17356 34932
rect 17236 34406 17264 34904
rect 17420 34746 17448 35634
rect 17408 34740 17460 34746
rect 17408 34682 17460 34688
rect 17696 34610 17724 36722
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17224 34400 17276 34406
rect 17224 34342 17276 34348
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 17052 32502 17080 32710
rect 17040 32496 17092 32502
rect 17040 32438 17092 32444
rect 17132 32360 17184 32366
rect 17132 32302 17184 32308
rect 17144 32026 17172 32302
rect 17132 32020 17184 32026
rect 17132 31962 17184 31968
rect 16960 31726 17080 31754
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16856 30320 16908 30326
rect 16856 30262 16908 30268
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16592 29714 16620 30126
rect 16580 29708 16632 29714
rect 16580 29650 16632 29656
rect 16592 29510 16620 29650
rect 16960 29510 16988 30534
rect 16580 29504 16632 29510
rect 16580 29446 16632 29452
rect 16948 29504 17000 29510
rect 16948 29446 17000 29452
rect 16592 27334 16620 29446
rect 16580 27328 16632 27334
rect 16580 27270 16632 27276
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16868 25906 16896 27066
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16868 21468 16896 24210
rect 16960 22166 16988 29446
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 16948 21480 17000 21486
rect 16868 21440 16948 21468
rect 16948 21422 17000 21428
rect 16764 21344 16816 21350
rect 16764 21286 16816 21292
rect 16776 20874 16804 21286
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16592 19990 16620 20402
rect 16960 20330 16988 21422
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 16592 17882 16620 18702
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16592 12152 16620 17206
rect 16960 17202 16988 17478
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 16684 15026 16712 15302
rect 16776 15094 16804 17138
rect 17052 17082 17080 31726
rect 17144 30054 17172 31962
rect 17132 30048 17184 30054
rect 17132 29990 17184 29996
rect 17144 29238 17172 29990
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 17132 28960 17184 28966
rect 17132 28902 17184 28908
rect 17236 28914 17264 34342
rect 17696 33998 17724 34546
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17408 33584 17460 33590
rect 17406 33552 17408 33561
rect 17460 33552 17462 33561
rect 17406 33487 17462 33496
rect 17316 33312 17368 33318
rect 17316 33254 17368 33260
rect 17328 29034 17356 33254
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17316 29028 17368 29034
rect 17316 28970 17368 28976
rect 17144 28558 17172 28902
rect 17236 28886 17356 28914
rect 17224 28756 17276 28762
rect 17224 28698 17276 28704
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17144 28218 17172 28494
rect 17132 28212 17184 28218
rect 17132 28154 17184 28160
rect 17236 28082 17264 28698
rect 17328 28422 17356 28886
rect 17316 28416 17368 28422
rect 17316 28358 17368 28364
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17236 27674 17264 28018
rect 17224 27668 17276 27674
rect 17224 27610 17276 27616
rect 17420 27130 17448 29038
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17408 27124 17460 27130
rect 17408 27066 17460 27072
rect 17408 26376 17460 26382
rect 17408 26318 17460 26324
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17328 26042 17356 26250
rect 17316 26036 17368 26042
rect 17316 25978 17368 25984
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17144 25158 17172 25842
rect 17316 25764 17368 25770
rect 17316 25706 17368 25712
rect 17224 25696 17276 25702
rect 17224 25638 17276 25644
rect 17132 25152 17184 25158
rect 17132 25094 17184 25100
rect 17144 24342 17172 25094
rect 17132 24336 17184 24342
rect 17132 24278 17184 24284
rect 17132 24132 17184 24138
rect 17132 24074 17184 24080
rect 17144 23798 17172 24074
rect 17236 24070 17264 25638
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 17236 23633 17264 23666
rect 17222 23624 17278 23633
rect 17222 23559 17278 23568
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 16960 17054 17080 17082
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16672 14408 16724 14414
rect 16776 14396 16804 15030
rect 16868 14414 16896 16390
rect 16724 14368 16804 14396
rect 16672 14350 16724 14356
rect 16776 12918 16804 14368
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16776 12238 16804 12718
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16672 12164 16724 12170
rect 16592 12124 16672 12152
rect 16672 12106 16724 12112
rect 16684 11898 16712 12106
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16776 11558 16804 12174
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16408 4678 16528 4706
rect 16408 3670 16436 4678
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16396 3664 16448 3670
rect 16396 3606 16448 3612
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16302 2680 16358 2689
rect 16302 2615 16358 2624
rect 16316 2582 16344 2615
rect 16304 2576 16356 2582
rect 16304 2518 16356 2524
rect 16396 1760 16448 1766
rect 16396 1702 16448 1708
rect 16408 800 16436 1702
rect 16500 800 16528 4558
rect 16592 3058 16620 8774
rect 16764 8560 16816 8566
rect 16762 8528 16764 8537
rect 16816 8528 16818 8537
rect 16762 8463 16818 8472
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16868 7478 16896 7958
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 6866 16712 7142
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16776 6712 16804 7210
rect 16684 6684 16804 6712
rect 16684 5846 16712 6684
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16684 5710 16712 5782
rect 16672 5704 16724 5710
rect 16672 5646 16724 5652
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16684 3194 16712 3946
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16592 2774 16620 2994
rect 16592 2746 16712 2774
rect 16684 800 16712 2746
rect 16776 800 16804 4966
rect 16868 3534 16896 6598
rect 16960 6202 16988 17054
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 10742 17080 15846
rect 17144 14890 17172 21966
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17236 20602 17264 21490
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17328 18850 17356 25706
rect 17420 24682 17448 26318
rect 17512 25906 17540 28358
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17592 26988 17644 26994
rect 17592 26930 17644 26936
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17604 25362 17632 26930
rect 17592 25356 17644 25362
rect 17592 25298 17644 25304
rect 17408 24676 17460 24682
rect 17408 24618 17460 24624
rect 17420 22982 17448 24618
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17408 22976 17460 22982
rect 17408 22918 17460 22924
rect 17420 22642 17448 22918
rect 17408 22636 17460 22642
rect 17408 22578 17460 22584
rect 17420 20942 17448 22578
rect 17512 22094 17540 24074
rect 17604 23186 17632 25298
rect 17592 23180 17644 23186
rect 17592 23122 17644 23128
rect 17512 22066 17632 22094
rect 17500 21072 17552 21078
rect 17500 21014 17552 21020
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17420 19378 17448 20878
rect 17512 19854 17540 21014
rect 17604 20466 17632 22066
rect 17696 22030 17724 27950
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 17788 26042 17816 26386
rect 17776 26036 17828 26042
rect 17776 25978 17828 25984
rect 17788 24750 17816 25978
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 17788 24206 17816 24686
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17776 24064 17828 24070
rect 17776 24006 17828 24012
rect 17788 23730 17816 24006
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17788 21554 17816 23666
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17776 20800 17828 20806
rect 17776 20742 17828 20748
rect 17788 20534 17816 20742
rect 17776 20528 17828 20534
rect 17776 20470 17828 20476
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17512 18970 17540 19314
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17328 18822 17632 18850
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17328 16794 17356 17614
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17420 16250 17448 16526
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17512 13258 17540 13806
rect 17500 13252 17552 13258
rect 17500 13194 17552 13200
rect 17512 12238 17540 13194
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17040 10736 17092 10742
rect 17040 10678 17092 10684
rect 17052 10266 17080 10678
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17052 9722 17080 10202
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 17052 6866 17080 9658
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17052 6390 17080 6802
rect 17040 6384 17092 6390
rect 17040 6326 17092 6332
rect 16960 6174 17080 6202
rect 16948 5092 17000 5098
rect 16948 5034 17000 5040
rect 16960 4146 16988 5034
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 17052 3738 17080 6174
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 2774 16896 3470
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16868 2746 16988 2774
rect 16960 800 16988 2746
rect 17052 800 17080 3130
rect 17144 2650 17172 10474
rect 17408 8900 17460 8906
rect 17408 8842 17460 8848
rect 17420 8634 17448 8842
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17316 7472 17368 7478
rect 17316 7414 17368 7420
rect 17328 6458 17356 7414
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17420 3602 17448 4558
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17132 2644 17184 2650
rect 17132 2586 17184 2592
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17236 800 17264 2450
rect 17328 800 17356 3062
rect 17512 800 17540 3470
rect 17604 3126 17632 18822
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17788 17610 17816 18566
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17788 17270 17816 17546
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17788 16658 17816 17206
rect 17776 16652 17828 16658
rect 17776 16594 17828 16600
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17788 14006 17816 15302
rect 17776 14000 17828 14006
rect 17776 13942 17828 13948
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17696 8129 17724 8230
rect 17682 8120 17738 8129
rect 17682 8055 17684 8064
rect 17736 8055 17738 8064
rect 17684 8026 17736 8032
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 17696 2774 17724 3878
rect 17880 3670 17908 55898
rect 18616 55690 18644 56306
rect 18604 55684 18656 55690
rect 18604 55626 18656 55632
rect 19076 55622 19104 56306
rect 19260 56234 19288 57394
rect 19340 57384 19392 57390
rect 19340 57326 19392 57332
rect 19352 56438 19380 57326
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 20640 56506 20668 57394
rect 20628 56500 20680 56506
rect 20628 56442 20680 56448
rect 19340 56432 19392 56438
rect 19340 56374 19392 56380
rect 20352 56364 20404 56370
rect 20352 56306 20404 56312
rect 20168 56296 20220 56302
rect 20168 56238 20220 56244
rect 19248 56228 19300 56234
rect 19248 56170 19300 56176
rect 19064 55616 19116 55622
rect 19064 55558 19116 55564
rect 18512 41268 18564 41274
rect 18512 41210 18564 41216
rect 17960 40928 18012 40934
rect 17960 40870 18012 40876
rect 17972 40526 18000 40870
rect 17960 40520 18012 40526
rect 17960 40462 18012 40468
rect 17972 38350 18000 40462
rect 18144 39432 18196 39438
rect 18144 39374 18196 39380
rect 17960 38344 18012 38350
rect 17960 38286 18012 38292
rect 18156 37874 18184 39374
rect 18144 37868 18196 37874
rect 18144 37810 18196 37816
rect 18236 37868 18288 37874
rect 18236 37810 18288 37816
rect 18248 37466 18276 37810
rect 18524 37466 18552 41210
rect 18604 38208 18656 38214
rect 18604 38150 18656 38156
rect 18236 37460 18288 37466
rect 18236 37402 18288 37408
rect 18512 37460 18564 37466
rect 18512 37402 18564 37408
rect 18524 37262 18552 37402
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 18328 34944 18380 34950
rect 18328 34886 18380 34892
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18340 34610 18368 34886
rect 18524 34678 18552 34886
rect 18512 34672 18564 34678
rect 18512 34614 18564 34620
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 18512 33924 18564 33930
rect 18512 33866 18564 33872
rect 18236 33312 18288 33318
rect 18236 33254 18288 33260
rect 18144 32972 18196 32978
rect 18144 32914 18196 32920
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 17972 31686 18000 32846
rect 18156 32570 18184 32914
rect 18248 32910 18276 33254
rect 18236 32904 18288 32910
rect 18236 32846 18288 32852
rect 18144 32564 18196 32570
rect 18144 32506 18196 32512
rect 18524 32502 18552 33866
rect 18512 32496 18564 32502
rect 18512 32438 18564 32444
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17972 30802 18000 31622
rect 18328 31476 18380 31482
rect 18328 31418 18380 31424
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 17972 30190 18000 30738
rect 18340 30734 18368 31418
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18512 30728 18564 30734
rect 18512 30670 18564 30676
rect 18052 30592 18104 30598
rect 18052 30534 18104 30540
rect 18064 30326 18092 30534
rect 18052 30320 18104 30326
rect 18052 30262 18104 30268
rect 17960 30184 18012 30190
rect 17960 30126 18012 30132
rect 17972 28626 18000 30126
rect 18524 29850 18552 30670
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18512 29232 18564 29238
rect 18512 29174 18564 29180
rect 18144 29164 18196 29170
rect 18144 29106 18196 29112
rect 18052 29028 18104 29034
rect 18052 28970 18104 28976
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17972 27470 18000 27882
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17972 24818 18000 26318
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17972 21146 18000 24754
rect 18064 22094 18092 28970
rect 18156 26994 18184 29106
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18432 27130 18460 27270
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18236 26920 18288 26926
rect 18236 26862 18288 26868
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18156 25702 18184 25842
rect 18144 25696 18196 25702
rect 18144 25638 18196 25644
rect 18248 25362 18276 26862
rect 18328 26852 18380 26858
rect 18328 26794 18380 26800
rect 18340 26586 18368 26794
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18236 25356 18288 25362
rect 18236 25298 18288 25304
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18156 24410 18184 24754
rect 18144 24404 18196 24410
rect 18144 24346 18196 24352
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18156 23594 18184 24142
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 18248 23730 18276 24006
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18144 23588 18196 23594
rect 18144 23530 18196 23536
rect 18248 23322 18276 23666
rect 18236 23316 18288 23322
rect 18236 23258 18288 23264
rect 18248 22166 18276 23258
rect 18236 22160 18288 22166
rect 18236 22102 18288 22108
rect 18064 22066 18184 22094
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 18156 20262 18184 22066
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 17972 18902 18000 20198
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18340 18766 18368 26522
rect 18420 25356 18472 25362
rect 18420 25298 18472 25304
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18064 18426 18092 18702
rect 18052 18420 18104 18426
rect 18052 18362 18104 18368
rect 18340 18222 18368 18702
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17972 16658 18000 17614
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 18064 16114 18092 16526
rect 18156 16522 18184 16934
rect 18248 16590 18276 18090
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18144 16516 18196 16522
rect 18144 16458 18196 16464
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17972 14618 18000 15914
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 18156 14550 18184 16458
rect 18340 15026 18368 16934
rect 18432 15706 18460 25298
rect 18524 24070 18552 29174
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18512 23656 18564 23662
rect 18510 23624 18512 23633
rect 18564 23624 18566 23633
rect 18510 23559 18566 23568
rect 18512 23520 18564 23526
rect 18512 23462 18564 23468
rect 18524 22710 18552 23462
rect 18512 22704 18564 22710
rect 18512 22646 18564 22652
rect 18616 22642 18644 38150
rect 18696 35012 18748 35018
rect 18696 34954 18748 34960
rect 18708 33522 18736 34954
rect 18972 34672 19024 34678
rect 18970 34640 18972 34649
rect 19024 34640 19026 34649
rect 18970 34575 19026 34584
rect 18696 33516 18748 33522
rect 18696 33458 18748 33464
rect 18708 32434 18736 33458
rect 18696 32428 18748 32434
rect 18696 32370 18748 32376
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18800 29170 18828 31758
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 18892 30326 18920 30670
rect 18880 30320 18932 30326
rect 18880 30262 18932 30268
rect 18788 29164 18840 29170
rect 18788 29106 18840 29112
rect 18892 29034 18920 30262
rect 18880 29028 18932 29034
rect 18880 28970 18932 28976
rect 18696 26784 18748 26790
rect 18696 26726 18748 26732
rect 18708 25906 18736 26726
rect 18788 25968 18840 25974
rect 18788 25910 18840 25916
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18708 25294 18736 25842
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18800 24342 18828 25910
rect 18892 25106 18920 28970
rect 19076 25770 19104 55558
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 20180 55214 20208 56238
rect 20364 56166 20392 56306
rect 20916 56234 20944 57462
rect 22192 57452 22244 57458
rect 22192 57394 22244 57400
rect 24400 57452 24452 57458
rect 24400 57394 24452 57400
rect 28448 57452 28500 57458
rect 28448 57394 28500 57400
rect 29000 57452 29052 57458
rect 29000 57394 29052 57400
rect 21088 57044 21140 57050
rect 21088 56986 21140 56992
rect 21100 56438 21128 56986
rect 21088 56432 21140 56438
rect 21088 56374 21140 56380
rect 21916 56364 21968 56370
rect 21916 56306 21968 56312
rect 20904 56228 20956 56234
rect 20904 56170 20956 56176
rect 20352 56160 20404 56166
rect 20350 56128 20352 56137
rect 20404 56128 20406 56137
rect 20350 56063 20406 56072
rect 21928 55622 21956 56306
rect 22204 55962 22232 57394
rect 22284 57248 22336 57254
rect 22284 57190 22336 57196
rect 22296 56506 22324 57190
rect 24412 56506 24440 57394
rect 28080 56704 28132 56710
rect 28080 56646 28132 56652
rect 22284 56500 22336 56506
rect 22284 56442 22336 56448
rect 24400 56500 24452 56506
rect 24400 56442 24452 56448
rect 28092 56438 28120 56646
rect 28460 56506 28488 57394
rect 28448 56500 28500 56506
rect 28448 56442 28500 56448
rect 28080 56432 28132 56438
rect 28080 56374 28132 56380
rect 23112 56364 23164 56370
rect 23112 56306 23164 56312
rect 23124 56273 23152 56306
rect 23110 56264 23166 56273
rect 29012 56234 29040 57394
rect 29184 56704 29236 56710
rect 29184 56646 29236 56652
rect 29196 56370 29224 56646
rect 29184 56364 29236 56370
rect 29184 56306 29236 56312
rect 30012 56364 30064 56370
rect 30012 56306 30064 56312
rect 30840 56364 30892 56370
rect 30840 56306 30892 56312
rect 23110 56199 23166 56208
rect 29000 56228 29052 56234
rect 29000 56170 29052 56176
rect 23572 56160 23624 56166
rect 23572 56102 23624 56108
rect 22192 55956 22244 55962
rect 22192 55898 22244 55904
rect 20444 55616 20496 55622
rect 20444 55558 20496 55564
rect 21916 55616 21968 55622
rect 21916 55558 21968 55564
rect 20180 55186 20300 55214
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19892 41744 19944 41750
rect 19892 41686 19944 41692
rect 19904 41614 19932 41686
rect 19892 41608 19944 41614
rect 19892 41550 19944 41556
rect 19340 41540 19392 41546
rect 19340 41482 19392 41488
rect 19352 41018 19380 41482
rect 19432 41472 19484 41478
rect 19904 41460 19932 41550
rect 20168 41540 20220 41546
rect 20168 41482 20220 41488
rect 19904 41432 20024 41460
rect 19432 41414 19484 41420
rect 19444 41206 19472 41414
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19432 41200 19484 41206
rect 19432 41142 19484 41148
rect 19996 41018 20024 41432
rect 20076 41132 20128 41138
rect 20076 41074 20128 41080
rect 19352 40990 19472 41018
rect 19340 40928 19392 40934
rect 19340 40870 19392 40876
rect 19248 40384 19300 40390
rect 19248 40326 19300 40332
rect 19260 40186 19288 40326
rect 19248 40180 19300 40186
rect 19248 40122 19300 40128
rect 19352 40032 19380 40870
rect 19444 40526 19472 40990
rect 19536 40990 20024 41018
rect 19536 40662 19564 40990
rect 19800 40928 19852 40934
rect 19800 40870 19852 40876
rect 19524 40656 19576 40662
rect 19524 40598 19576 40604
rect 19812 40526 19840 40870
rect 19904 40526 19932 40990
rect 19984 40656 20036 40662
rect 19984 40598 20036 40604
rect 19432 40520 19484 40526
rect 19432 40462 19484 40468
rect 19800 40520 19852 40526
rect 19800 40462 19852 40468
rect 19892 40520 19944 40526
rect 19892 40462 19944 40468
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19524 40180 19576 40186
rect 19524 40122 19576 40128
rect 19260 40004 19380 40032
rect 19260 39846 19288 40004
rect 19248 39840 19300 39846
rect 19248 39782 19300 39788
rect 19260 39438 19288 39782
rect 19536 39438 19564 40122
rect 19248 39432 19300 39438
rect 19248 39374 19300 39380
rect 19524 39432 19576 39438
rect 19524 39374 19576 39380
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 38752 19484 38758
rect 19432 38694 19484 38700
rect 19248 38480 19300 38486
rect 19248 38422 19300 38428
rect 19156 38412 19208 38418
rect 19156 38354 19208 38360
rect 19168 37874 19196 38354
rect 19260 38350 19288 38422
rect 19248 38344 19300 38350
rect 19248 38286 19300 38292
rect 19340 38344 19392 38350
rect 19340 38286 19392 38292
rect 19248 38208 19300 38214
rect 19248 38150 19300 38156
rect 19156 37868 19208 37874
rect 19156 37810 19208 37816
rect 19260 37482 19288 38150
rect 19352 37670 19380 38286
rect 19444 37942 19472 38694
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19432 37936 19484 37942
rect 19432 37878 19484 37884
rect 19708 37868 19760 37874
rect 19708 37810 19760 37816
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 19260 37454 19380 37482
rect 19352 37448 19380 37454
rect 19352 37420 19472 37448
rect 19340 37256 19392 37262
rect 19340 37198 19392 37204
rect 19156 37120 19208 37126
rect 19156 37062 19208 37068
rect 19168 34542 19196 37062
rect 19248 36916 19300 36922
rect 19248 36858 19300 36864
rect 19156 34536 19208 34542
rect 19156 34478 19208 34484
rect 19168 33658 19196 34478
rect 19260 34202 19288 36858
rect 19352 36650 19380 37198
rect 19444 37194 19472 37420
rect 19720 37262 19748 37810
rect 19996 37754 20024 40598
rect 20088 39302 20116 41074
rect 20180 40730 20208 41482
rect 20168 40724 20220 40730
rect 20168 40666 20220 40672
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 20088 38282 20116 39238
rect 20076 38276 20128 38282
rect 20076 38218 20128 38224
rect 20168 38208 20220 38214
rect 20168 38150 20220 38156
rect 20180 37874 20208 38150
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 19996 37738 20208 37754
rect 19996 37732 20220 37738
rect 19996 37726 20168 37732
rect 20168 37674 20220 37680
rect 20076 37664 20128 37670
rect 20076 37606 20128 37612
rect 19708 37256 19760 37262
rect 19708 37198 19760 37204
rect 19432 37188 19484 37194
rect 19432 37130 19484 37136
rect 19340 36644 19392 36650
rect 19340 36586 19392 36592
rect 19444 34649 19472 37130
rect 19720 37126 19748 37198
rect 19708 37120 19760 37126
rect 19708 37062 19760 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 20088 36922 20116 37606
rect 20076 36916 20128 36922
rect 20076 36858 20128 36864
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 20076 35080 20128 35086
rect 20076 35022 20128 35028
rect 19984 34944 20036 34950
rect 19984 34886 20036 34892
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19430 34640 19486 34649
rect 19430 34575 19486 34584
rect 19996 34490 20024 34886
rect 20088 34746 20116 35022
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 19904 34462 20024 34490
rect 19248 34196 19300 34202
rect 19248 34138 19300 34144
rect 19260 33998 19288 34138
rect 19904 33998 19932 34462
rect 20180 34354 20208 37674
rect 19996 34326 20208 34354
rect 19996 33998 20024 34326
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19892 33992 19944 33998
rect 19892 33934 19944 33940
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 19260 33658 19288 33934
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 19260 33114 19288 33254
rect 19248 33108 19300 33114
rect 19248 33050 19300 33056
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19156 31136 19208 31142
rect 19156 31078 19208 31084
rect 19168 30240 19196 31078
rect 19260 30802 19288 32846
rect 19996 32774 20024 33934
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 20272 31754 20300 55186
rect 20456 42770 20484 55558
rect 21928 55214 21956 55558
rect 21928 55186 22048 55214
rect 20444 42764 20496 42770
rect 20444 42706 20496 42712
rect 20352 41676 20404 41682
rect 20352 41618 20404 41624
rect 20364 40662 20392 41618
rect 20720 41132 20772 41138
rect 20720 41074 20772 41080
rect 20628 40996 20680 41002
rect 20628 40938 20680 40944
rect 20352 40656 20404 40662
rect 20352 40598 20404 40604
rect 20640 40594 20668 40938
rect 20628 40588 20680 40594
rect 20628 40530 20680 40536
rect 20444 40520 20496 40526
rect 20444 40462 20496 40468
rect 20352 40452 20404 40458
rect 20352 40394 20404 40400
rect 20364 39846 20392 40394
rect 20352 39840 20404 39846
rect 20352 39782 20404 39788
rect 20364 38350 20392 39782
rect 20352 38344 20404 38350
rect 20352 38286 20404 38292
rect 20352 38004 20404 38010
rect 20352 37946 20404 37952
rect 20364 33998 20392 37946
rect 20456 37670 20484 40462
rect 20732 40390 20760 41074
rect 21364 40452 21416 40458
rect 21364 40394 21416 40400
rect 21916 40452 21968 40458
rect 21916 40394 21968 40400
rect 20720 40384 20772 40390
rect 20720 40326 20772 40332
rect 20628 38820 20680 38826
rect 20628 38762 20680 38768
rect 20536 38276 20588 38282
rect 20536 38218 20588 38224
rect 20444 37664 20496 37670
rect 20444 37606 20496 37612
rect 20548 37466 20576 38218
rect 20640 37806 20668 38762
rect 20732 38282 20760 40326
rect 21376 39642 21404 40394
rect 21928 39982 21956 40394
rect 21916 39976 21968 39982
rect 21916 39918 21968 39924
rect 21824 39840 21876 39846
rect 21824 39782 21876 39788
rect 21364 39636 21416 39642
rect 21364 39578 21416 39584
rect 21836 39438 21864 39782
rect 21640 39432 21692 39438
rect 21640 39374 21692 39380
rect 21824 39432 21876 39438
rect 21824 39374 21876 39380
rect 21652 38758 21680 39374
rect 21928 39370 21956 39918
rect 21916 39364 21968 39370
rect 21916 39306 21968 39312
rect 21640 38752 21692 38758
rect 21640 38694 21692 38700
rect 21088 38480 21140 38486
rect 21088 38422 21140 38428
rect 20720 38276 20772 38282
rect 20720 38218 20772 38224
rect 20628 37800 20680 37806
rect 20628 37742 20680 37748
rect 20536 37460 20588 37466
rect 20536 37402 20588 37408
rect 20640 37346 20668 37742
rect 20548 37318 20668 37346
rect 20352 33992 20404 33998
rect 20352 33934 20404 33940
rect 20364 33386 20392 33934
rect 20352 33380 20404 33386
rect 20352 33322 20404 33328
rect 20180 31726 20300 31754
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 19996 31142 20024 31282
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 19248 30796 19300 30802
rect 19248 30738 19300 30744
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19444 30394 19472 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19248 30252 19300 30258
rect 19168 30212 19248 30240
rect 19248 30194 19300 30200
rect 19260 29238 19288 30194
rect 19340 30048 19392 30054
rect 19340 29990 19392 29996
rect 19352 29646 19380 29990
rect 19996 29646 20024 31078
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 19340 29640 19392 29646
rect 19340 29582 19392 29588
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19248 29232 19300 29238
rect 19248 29174 19300 29180
rect 19352 29170 19380 29582
rect 20088 29578 20116 30534
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19444 28694 19472 29174
rect 19984 29096 20036 29102
rect 19984 29038 20036 29044
rect 19432 28688 19484 28694
rect 19432 28630 19484 28636
rect 19444 28082 19472 28630
rect 19996 28558 20024 29038
rect 20088 28626 20116 29514
rect 20076 28620 20128 28626
rect 20076 28562 20128 28568
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19996 28082 20024 28494
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 19340 28008 19392 28014
rect 19340 27950 19392 27956
rect 19156 27872 19208 27878
rect 19156 27814 19208 27820
rect 19168 27470 19196 27814
rect 19156 27464 19208 27470
rect 19156 27406 19208 27412
rect 19064 25764 19116 25770
rect 19064 25706 19116 25712
rect 19168 25242 19196 27406
rect 19352 26602 19380 27950
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19616 27056 19668 27062
rect 19616 26998 19668 27004
rect 19260 26574 19380 26602
rect 19260 25362 19288 26574
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19352 25888 19380 26454
rect 19628 26382 19656 26998
rect 19892 26988 19944 26994
rect 19892 26930 19944 26936
rect 19904 26586 19932 26930
rect 19892 26580 19944 26586
rect 19892 26522 19944 26528
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19444 26042 19472 26318
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 19432 25900 19484 25906
rect 19352 25860 19432 25888
rect 19432 25842 19484 25848
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19168 25214 19288 25242
rect 18892 25078 19196 25106
rect 18788 24336 18840 24342
rect 18788 24278 18840 24284
rect 18800 24138 18828 24278
rect 18788 24132 18840 24138
rect 18788 24074 18840 24080
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18880 21140 18932 21146
rect 18880 21082 18932 21088
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18512 17332 18564 17338
rect 18512 17274 18564 17280
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18420 15496 18472 15502
rect 18420 15438 18472 15444
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18432 14822 18460 15438
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18144 14544 18196 14550
rect 18144 14486 18196 14492
rect 18432 14482 18460 14758
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18524 14362 18552 17274
rect 18800 17202 18828 17750
rect 18788 17196 18840 17202
rect 18788 17138 18840 17144
rect 18248 14334 18552 14362
rect 17960 13456 18012 13462
rect 17960 13398 18012 13404
rect 17972 8634 18000 13398
rect 18248 12442 18276 14334
rect 18236 12436 18288 12442
rect 18236 12378 18288 12384
rect 18144 12368 18196 12374
rect 18196 12316 18368 12322
rect 18144 12310 18368 12316
rect 18156 12294 18368 12310
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11762 18184 12038
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18248 11082 18276 12174
rect 18340 12102 18368 12294
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18340 10470 18368 11698
rect 18708 11354 18736 12174
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 8974 18368 10406
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 9382 18460 9522
rect 18800 9382 18828 11018
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17958 8528 18014 8537
rect 17958 8463 17960 8472
rect 18012 8463 18014 8472
rect 17960 8434 18012 8440
rect 17972 8090 18000 8434
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17788 3058 17816 3402
rect 17972 3058 18000 7142
rect 18340 6730 18368 7278
rect 18328 6724 18380 6730
rect 18328 6666 18380 6672
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18052 5704 18104 5710
rect 18052 5646 18104 5652
rect 18064 5234 18092 5646
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18156 4842 18184 5850
rect 18248 5710 18276 6054
rect 18340 5846 18368 6666
rect 18432 6662 18460 9318
rect 18800 8838 18828 9318
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18708 8362 18736 8434
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18708 7954 18736 8298
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18708 7410 18736 7890
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 6254 18460 6598
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18340 5166 18368 5782
rect 18524 5642 18552 6122
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18064 4814 18184 4842
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17604 2746 17724 2774
rect 17604 800 17632 2746
rect 17682 2680 17738 2689
rect 17682 2615 17684 2624
rect 17736 2615 17738 2624
rect 17684 2586 17736 2592
rect 17788 800 17816 2994
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 17960 2916 18012 2922
rect 17960 2858 18012 2864
rect 17880 800 17908 2858
rect 17972 2446 18000 2858
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18064 2378 18092 4814
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18064 800 18092 2314
rect 18156 800 18184 4694
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 3534 18368 4422
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18234 3224 18290 3233
rect 18234 3159 18236 3168
rect 18288 3159 18290 3168
rect 18236 3130 18288 3136
rect 18340 800 18368 3470
rect 18432 800 18460 4966
rect 18524 4010 18552 5578
rect 18616 5234 18644 6190
rect 18800 5710 18828 6734
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18512 2576 18564 2582
rect 18510 2544 18512 2553
rect 18564 2544 18566 2553
rect 18510 2479 18566 2488
rect 18616 800 18644 2994
rect 18708 800 18736 3538
rect 18800 2106 18828 5646
rect 18892 3738 18920 21082
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18984 19242 19012 19450
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 18984 18358 19012 19178
rect 18972 18352 19024 18358
rect 18972 18294 19024 18300
rect 19168 17678 19196 25078
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19168 17202 19196 17614
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 18984 16794 19012 17138
rect 18972 16788 19024 16794
rect 18972 16730 19024 16736
rect 19260 16266 19288 25214
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19352 24954 19380 25094
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19352 24614 19380 24754
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19352 22778 19380 23598
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19352 17066 19380 22374
rect 19444 20641 19472 25842
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19430 20632 19486 20641
rect 19574 20635 19882 20644
rect 19430 20567 19486 20576
rect 19616 20528 19668 20534
rect 19430 20496 19486 20505
rect 19616 20470 19668 20476
rect 19430 20431 19486 20440
rect 19524 20460 19576 20466
rect 19444 20330 19472 20431
rect 19524 20402 19576 20408
rect 19536 20330 19564 20402
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19628 20058 19656 20470
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19812 20369 19840 20402
rect 19798 20360 19854 20369
rect 19798 20295 19854 20304
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19996 19786 20024 27270
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 20088 25430 20116 26318
rect 20076 25424 20128 25430
rect 20076 25366 20128 25372
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 20088 20466 20116 21422
rect 20180 21146 20208 31726
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20272 29850 20300 30194
rect 20352 30184 20404 30190
rect 20352 30126 20404 30132
rect 20260 29844 20312 29850
rect 20260 29786 20312 29792
rect 20364 29510 20392 30126
rect 20352 29504 20404 29510
rect 20352 29446 20404 29452
rect 20352 29028 20404 29034
rect 20352 28970 20404 28976
rect 20260 26240 20312 26246
rect 20260 26182 20312 26188
rect 20272 25974 20300 26182
rect 20260 25968 20312 25974
rect 20260 25910 20312 25916
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20777 20208 20810
rect 20260 20800 20312 20806
rect 20166 20768 20222 20777
rect 20260 20742 20312 20748
rect 20166 20703 20222 20712
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20180 20262 20208 20538
rect 20272 20534 20300 20742
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 20272 20398 20300 20470
rect 20364 20466 20392 28970
rect 20548 28966 20576 37318
rect 20732 35018 20760 38218
rect 20996 37664 21048 37670
rect 20996 37606 21048 37612
rect 21008 37262 21036 37606
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 20904 37120 20956 37126
rect 20904 37062 20956 37068
rect 20812 35216 20864 35222
rect 20812 35158 20864 35164
rect 20720 35012 20772 35018
rect 20720 34954 20772 34960
rect 20720 34604 20772 34610
rect 20720 34546 20772 34552
rect 20732 34202 20760 34546
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 20640 33046 20668 33390
rect 20628 33040 20680 33046
rect 20628 32982 20680 32988
rect 20824 32366 20852 35158
rect 20812 32360 20864 32366
rect 20812 32302 20864 32308
rect 20916 31754 20944 37062
rect 21100 31754 21128 38422
rect 21652 36242 21680 38694
rect 21824 37256 21876 37262
rect 21824 37198 21876 37204
rect 21640 36236 21692 36242
rect 21640 36178 21692 36184
rect 21732 36032 21784 36038
rect 21732 35974 21784 35980
rect 21180 35556 21232 35562
rect 21180 35498 21232 35504
rect 21192 32570 21220 35498
rect 21640 34944 21692 34950
rect 21640 34886 21692 34892
rect 21652 34678 21680 34886
rect 21640 34672 21692 34678
rect 21640 34614 21692 34620
rect 21180 32564 21232 32570
rect 21180 32506 21232 32512
rect 21640 32564 21692 32570
rect 21640 32506 21692 32512
rect 21364 32292 21416 32298
rect 21364 32234 21416 32240
rect 20916 31726 21036 31754
rect 21100 31726 21312 31754
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20548 27062 20576 28902
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20536 27056 20588 27062
rect 20536 26998 20588 27004
rect 20536 26920 20588 26926
rect 20640 26908 20668 27338
rect 20588 26880 20668 26908
rect 20536 26862 20588 26868
rect 20444 26376 20496 26382
rect 20444 26318 20496 26324
rect 20456 25702 20484 26318
rect 20548 25838 20576 26862
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20812 26376 20864 26382
rect 20812 26318 20864 26324
rect 20640 26042 20668 26318
rect 20628 26036 20680 26042
rect 20628 25978 20680 25984
rect 20824 25974 20852 26318
rect 20812 25968 20864 25974
rect 20812 25910 20864 25916
rect 20536 25832 20588 25838
rect 20536 25774 20588 25780
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20548 24886 20576 25774
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 20536 24880 20588 24886
rect 20536 24822 20588 24828
rect 20442 23080 20498 23089
rect 20442 23015 20444 23024
rect 20496 23015 20498 23024
rect 20444 22986 20496 22992
rect 20536 22976 20588 22982
rect 20536 22918 20588 22924
rect 20548 22094 20576 22918
rect 20628 22772 20680 22778
rect 20628 22714 20680 22720
rect 20456 22066 20576 22094
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19340 17060 19392 17066
rect 19340 17002 19392 17008
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19340 16448 19392 16454
rect 19340 16390 19392 16396
rect 19168 16238 19288 16266
rect 19168 13734 19196 16238
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19260 15094 19288 16118
rect 19352 16114 19380 16390
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19352 15706 19380 16050
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19352 14414 19380 15302
rect 19444 14890 19472 16458
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 15706 19932 15846
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19904 15434 19932 15642
rect 19892 15428 19944 15434
rect 19892 15370 19944 15376
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 20180 14482 20208 14962
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19984 14408 20036 14414
rect 19984 14350 20036 14356
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19352 14006 19380 14350
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19168 12850 19196 13126
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18984 12306 19012 12650
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 19168 11626 19196 12582
rect 19260 12374 19288 12786
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19156 11620 19208 11626
rect 19156 11562 19208 11568
rect 19168 11082 19196 11562
rect 19156 11076 19208 11082
rect 19156 11018 19208 11024
rect 19352 10470 19380 11698
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 18984 8498 19012 9590
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 19076 8634 19104 8842
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18984 8294 19012 8434
rect 19248 8424 19300 8430
rect 19248 8366 19300 8372
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 19260 8090 19288 8366
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19352 7426 19380 10406
rect 19444 9722 19472 13262
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12434 20024 14350
rect 20088 13938 20116 14350
rect 20180 14278 20208 14418
rect 20272 14414 20300 20334
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20364 15706 20392 17614
rect 20352 15700 20404 15706
rect 20352 15642 20404 15648
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20364 15366 20392 15438
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 19996 12406 20116 12434
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11898 20024 12106
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 20088 9654 20116 12406
rect 20180 12238 20208 13806
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20456 11830 20484 22066
rect 20640 22012 20668 22714
rect 20824 22642 20852 25094
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 21008 22438 21036 31726
rect 21180 31272 21232 31278
rect 21180 31214 21232 31220
rect 21192 30326 21220 31214
rect 21180 30320 21232 30326
rect 21180 30262 21232 30268
rect 21088 28416 21140 28422
rect 21088 28358 21140 28364
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 20548 21984 20668 22012
rect 20548 21078 20576 21984
rect 20536 21072 20588 21078
rect 20536 21014 20588 21020
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20536 20528 20588 20534
rect 20534 20496 20536 20505
rect 20588 20496 20590 20505
rect 20640 20466 20668 20810
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20534 20431 20590 20440
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20640 20058 20668 20402
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20548 18698 20576 19314
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20548 18290 20576 18634
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20732 16674 20760 20470
rect 20916 18850 20944 22374
rect 21100 22094 21128 28358
rect 21180 27940 21232 27946
rect 21180 27882 21232 27888
rect 21192 27062 21220 27882
rect 21180 27056 21232 27062
rect 21180 26998 21232 27004
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 21192 22642 21220 24006
rect 21180 22636 21232 22642
rect 21180 22578 21232 22584
rect 21284 22234 21312 31726
rect 21376 25378 21404 32234
rect 21652 31346 21680 32506
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21548 30728 21600 30734
rect 21548 30670 21600 30676
rect 21456 29164 21508 29170
rect 21456 29106 21508 29112
rect 21468 28694 21496 29106
rect 21456 28688 21508 28694
rect 21456 28630 21508 28636
rect 21468 28490 21496 28630
rect 21456 28484 21508 28490
rect 21456 28426 21508 28432
rect 21560 27402 21588 30670
rect 21652 27946 21680 31282
rect 21744 28914 21772 35974
rect 21836 35766 21864 37198
rect 21824 35760 21876 35766
rect 21824 35702 21876 35708
rect 21836 34610 21864 35702
rect 21928 34950 21956 39306
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 21824 34604 21876 34610
rect 21824 34546 21876 34552
rect 21928 34490 21956 34886
rect 21836 34462 21956 34490
rect 21836 31278 21864 34462
rect 21916 32768 21968 32774
rect 21916 32710 21968 32716
rect 21928 32434 21956 32710
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 21824 31272 21876 31278
rect 21824 31214 21876 31220
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21928 30666 21956 31078
rect 21916 30660 21968 30666
rect 21916 30602 21968 30608
rect 21744 28886 21864 28914
rect 21640 27940 21692 27946
rect 21640 27882 21692 27888
rect 21548 27396 21600 27402
rect 21548 27338 21600 27344
rect 21732 26376 21784 26382
rect 21730 26344 21732 26353
rect 21784 26344 21786 26353
rect 21640 26308 21692 26314
rect 21730 26279 21786 26288
rect 21640 26250 21692 26256
rect 21456 26240 21508 26246
rect 21456 26182 21508 26188
rect 21468 25974 21496 26182
rect 21652 25974 21680 26250
rect 21456 25968 21508 25974
rect 21456 25910 21508 25916
rect 21640 25968 21692 25974
rect 21640 25910 21692 25916
rect 21548 25424 21600 25430
rect 21376 25350 21496 25378
rect 21548 25366 21600 25372
rect 21364 25288 21416 25294
rect 21364 25230 21416 25236
rect 21376 24818 21404 25230
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21376 24206 21404 24754
rect 21364 24200 21416 24206
rect 21364 24142 21416 24148
rect 21376 23662 21404 24142
rect 21364 23656 21416 23662
rect 21364 23598 21416 23604
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21008 22066 21128 22094
rect 21008 20942 21036 22066
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 21100 21690 21128 21966
rect 21180 21888 21232 21894
rect 21180 21830 21232 21836
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 21100 20466 21128 20810
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 21008 19446 21036 20198
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 20916 18822 21036 18850
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20824 17746 20852 18702
rect 20904 18692 20956 18698
rect 20904 18634 20956 18640
rect 20916 18426 20944 18634
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20812 17740 20864 17746
rect 20812 17682 20864 17688
rect 20640 16646 20760 16674
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 15502 20576 16050
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20640 12238 20668 16646
rect 20824 16250 20852 17682
rect 21008 17338 21036 18822
rect 21192 18086 21220 21830
rect 21376 21146 21404 23598
rect 21468 23594 21496 25350
rect 21560 23866 21588 25366
rect 21732 24608 21784 24614
rect 21732 24550 21784 24556
rect 21744 24206 21772 24550
rect 21732 24200 21784 24206
rect 21836 24188 21864 28886
rect 21916 27056 21968 27062
rect 21916 26998 21968 27004
rect 21928 26382 21956 26998
rect 21916 26376 21968 26382
rect 21916 26318 21968 26324
rect 21916 25220 21968 25226
rect 21916 25162 21968 25168
rect 21928 24886 21956 25162
rect 21916 24880 21968 24886
rect 21916 24822 21968 24828
rect 21916 24200 21968 24206
rect 21836 24160 21916 24188
rect 21732 24142 21784 24148
rect 21916 24142 21968 24148
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21652 23769 21680 24074
rect 21638 23760 21694 23769
rect 21638 23695 21694 23704
rect 21456 23588 21508 23594
rect 21456 23530 21508 23536
rect 21652 21622 21680 23695
rect 22020 22094 22048 55186
rect 23020 41268 23072 41274
rect 23020 41210 23072 41216
rect 22100 41132 22152 41138
rect 22100 41074 22152 41080
rect 22112 40186 22140 41074
rect 23032 40934 23060 41210
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 22652 40928 22704 40934
rect 22652 40870 22704 40876
rect 23020 40928 23072 40934
rect 23020 40870 23072 40876
rect 22284 40520 22336 40526
rect 22284 40462 22336 40468
rect 22100 40180 22152 40186
rect 22100 40122 22152 40128
rect 22192 40180 22244 40186
rect 22192 40122 22244 40128
rect 22112 39098 22140 40122
rect 22100 39092 22152 39098
rect 22100 39034 22152 39040
rect 22204 37806 22232 40122
rect 22296 40050 22324 40462
rect 22560 40384 22612 40390
rect 22560 40326 22612 40332
rect 22572 40118 22600 40326
rect 22560 40112 22612 40118
rect 22560 40054 22612 40060
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22296 39438 22324 39986
rect 22284 39432 22336 39438
rect 22284 39374 22336 39380
rect 22192 37800 22244 37806
rect 22192 37742 22244 37748
rect 22100 36236 22152 36242
rect 22100 36178 22152 36184
rect 22112 32570 22140 36178
rect 22192 36168 22244 36174
rect 22192 36110 22244 36116
rect 22204 36038 22232 36110
rect 22192 36032 22244 36038
rect 22192 35974 22244 35980
rect 22204 35698 22232 35974
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22112 30598 22140 32506
rect 22100 30592 22152 30598
rect 22100 30534 22152 30540
rect 22204 30410 22232 35634
rect 22296 35086 22324 39374
rect 22376 36576 22428 36582
rect 22376 36518 22428 36524
rect 22388 36106 22416 36518
rect 22572 36174 22600 40054
rect 22664 40050 22692 40870
rect 23032 40526 23060 40870
rect 22744 40520 22796 40526
rect 22744 40462 22796 40468
rect 23020 40520 23072 40526
rect 23020 40462 23072 40468
rect 22652 40044 22704 40050
rect 22652 39986 22704 39992
rect 22652 39296 22704 39302
rect 22652 39238 22704 39244
rect 22664 38962 22692 39238
rect 22756 39098 22784 40462
rect 23400 39846 23428 41074
rect 23480 40384 23532 40390
rect 23480 40326 23532 40332
rect 23388 39840 23440 39846
rect 23388 39782 23440 39788
rect 22744 39092 22796 39098
rect 22744 39034 22796 39040
rect 23020 39024 23072 39030
rect 23020 38966 23072 38972
rect 22652 38956 22704 38962
rect 22652 38898 22704 38904
rect 22836 37120 22888 37126
rect 22836 37062 22888 37068
rect 22848 36786 22876 37062
rect 22836 36780 22888 36786
rect 22836 36722 22888 36728
rect 22848 36174 22876 36722
rect 22928 36576 22980 36582
rect 22928 36518 22980 36524
rect 22560 36168 22612 36174
rect 22560 36110 22612 36116
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 22376 36100 22428 36106
rect 22376 36042 22428 36048
rect 22848 36038 22876 36110
rect 22836 36032 22888 36038
rect 22836 35974 22888 35980
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 22468 35488 22520 35494
rect 22848 35442 22876 35634
rect 22468 35430 22520 35436
rect 22284 35080 22336 35086
rect 22284 35022 22336 35028
rect 22284 31204 22336 31210
rect 22284 31146 22336 31152
rect 22296 30734 22324 31146
rect 22284 30728 22336 30734
rect 22284 30670 22336 30676
rect 22112 30382 22232 30410
rect 22112 28626 22140 30382
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22204 29646 22232 30194
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22204 28422 22232 29582
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 21928 22066 22048 22094
rect 21640 21616 21692 21622
rect 21640 21558 21692 21564
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21836 21146 21864 21354
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 21822 20768 21878 20777
rect 21822 20703 21878 20712
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21180 18080 21232 18086
rect 21180 18022 21232 18028
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20916 13462 20944 16662
rect 21008 16114 21036 17070
rect 21192 16794 21220 17546
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 21560 16726 21588 18634
rect 21836 17542 21864 20703
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21836 17270 21864 17478
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21732 16992 21784 16998
rect 21732 16934 21784 16940
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21272 16108 21324 16114
rect 21272 16050 21324 16056
rect 20996 15156 21048 15162
rect 20996 15098 21048 15104
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20732 12238 20760 13194
rect 21008 12850 21036 15098
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21192 13530 21220 14962
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21008 12238 21036 12786
rect 21192 12442 21220 13466
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 11830 20668 12038
rect 20444 11824 20496 11830
rect 20444 11766 20496 11772
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20732 11762 20760 12174
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20548 11354 20576 11698
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20076 9648 20128 9654
rect 20076 9590 20128 9596
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19444 7886 19472 9114
rect 20272 9110 20300 9522
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20364 9178 20392 9386
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20260 9104 20312 9110
rect 20260 9046 20312 9052
rect 20548 8974 20576 9590
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 20640 8566 20668 9114
rect 21284 8974 21312 16050
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21376 14822 21404 15302
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 14346 21404 14758
rect 21468 14482 21496 15370
rect 21560 15162 21588 16662
rect 21744 16658 21772 16934
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21652 15366 21680 16050
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21836 12986 21864 13670
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21732 12164 21784 12170
rect 21836 12152 21864 12922
rect 21784 12124 21864 12152
rect 21732 12106 21784 12112
rect 21548 11688 21600 11694
rect 21548 11630 21600 11636
rect 21560 11218 21588 11630
rect 21548 11212 21600 11218
rect 21548 11154 21600 11160
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21284 8634 21312 8910
rect 21272 8628 21324 8634
rect 21272 8570 21324 8576
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19996 7818 20024 8434
rect 19984 7812 20036 7818
rect 19984 7754 20036 7760
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19352 7398 19472 7426
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19352 6390 19380 7142
rect 19444 6866 19472 7398
rect 19996 7274 20024 7754
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19248 6248 19300 6254
rect 19248 6190 19300 6196
rect 19260 5710 19288 6190
rect 19444 5914 19472 6258
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19536 5794 19564 6258
rect 19444 5766 19564 5794
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18878 3224 18934 3233
rect 18878 3159 18880 3168
rect 18932 3159 18934 3168
rect 18880 3130 18932 3136
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18892 2922 18920 2994
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18892 800 18920 2858
rect 18984 800 19012 4626
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19168 3720 19196 4558
rect 19260 4146 19288 5646
rect 19340 5568 19392 5574
rect 19444 5556 19472 5766
rect 19392 5528 19472 5556
rect 19340 5510 19392 5516
rect 19444 5302 19472 5528
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19432 5092 19484 5098
rect 19432 5034 19484 5040
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19168 3692 19288 3720
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19076 3058 19104 3606
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19076 2774 19104 2994
rect 19076 2746 19196 2774
rect 19168 800 19196 2746
rect 19260 800 19288 3692
rect 19352 1494 19380 4558
rect 19444 4214 19472 5034
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19444 3108 19472 3878
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19536 3398 19564 3470
rect 19524 3392 19576 3398
rect 19505 3340 19524 3380
rect 19505 3334 19576 3340
rect 19505 3176 19533 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19505 3148 19748 3176
rect 19444 3080 19656 3108
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19340 1488 19392 1494
rect 19340 1430 19392 1436
rect 19444 1442 19472 2790
rect 19628 2650 19656 3080
rect 19616 2644 19668 2650
rect 19616 2586 19668 2592
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19720 2394 19748 3148
rect 19996 3058 20024 6598
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19996 2514 20024 2994
rect 19984 2508 20036 2514
rect 19984 2450 20036 2456
rect 19536 2292 19564 2382
rect 19720 2366 20024 2394
rect 19505 2264 19564 2292
rect 19505 2088 19533 2264
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19505 2060 19656 2088
rect 19444 1414 19564 1442
rect 19432 1352 19484 1358
rect 19432 1294 19484 1300
rect 19444 800 19472 1294
rect 19536 800 19564 1414
rect 19628 1358 19656 2060
rect 19800 1488 19852 1494
rect 19800 1430 19852 1436
rect 19708 1420 19760 1426
rect 19708 1362 19760 1368
rect 19616 1352 19668 1358
rect 19616 1294 19668 1300
rect 19720 800 19748 1362
rect 19812 800 19840 1430
rect 19996 800 20024 2366
rect 20088 800 20116 4966
rect 20180 2774 20208 6666
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20272 3126 20300 6054
rect 20442 5672 20498 5681
rect 20442 5607 20498 5616
rect 20350 4040 20406 4049
rect 20350 3975 20406 3984
rect 20364 3194 20392 3975
rect 20456 3738 20484 5607
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20548 3210 20576 6394
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20456 3182 20576 3210
rect 20260 3120 20312 3126
rect 20260 3062 20312 3068
rect 20456 2774 20484 3182
rect 20536 3120 20588 3126
rect 20536 3062 20588 3068
rect 20180 2746 20300 2774
rect 20168 2508 20220 2514
rect 20168 2450 20220 2456
rect 20180 1426 20208 2450
rect 20272 2378 20300 2746
rect 20364 2746 20484 2774
rect 20364 2582 20392 2746
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20352 2576 20404 2582
rect 20352 2518 20404 2524
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20168 1420 20220 1426
rect 20168 1362 20220 1368
rect 20272 800 20300 2314
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20364 2038 20392 2246
rect 20352 2032 20404 2038
rect 20352 1974 20404 1980
rect 20456 1442 20484 2586
rect 20364 1414 20484 1442
rect 20364 800 20392 1414
rect 20548 800 20576 3062
rect 20640 800 20668 4558
rect 20732 2446 20760 6598
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20824 3534 20852 6054
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20732 1766 20760 2382
rect 20720 1760 20772 1766
rect 20720 1702 20772 1708
rect 20824 800 20852 3470
rect 20916 800 20944 4966
rect 21008 2514 21036 6598
rect 21376 5234 21404 8910
rect 21744 7750 21772 12106
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 21836 11150 21864 11494
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21824 9512 21876 9518
rect 21824 9454 21876 9460
rect 21836 9042 21864 9454
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21836 6254 21864 6734
rect 21928 6458 21956 22066
rect 22112 22030 22140 24550
rect 22204 23866 22232 25434
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 22204 22030 22232 23802
rect 22296 22982 22324 30670
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22388 23730 22416 29990
rect 22480 28506 22508 35430
rect 22664 35414 22876 35442
rect 22560 35080 22612 35086
rect 22560 35022 22612 35028
rect 22572 31958 22600 35022
rect 22560 31952 22612 31958
rect 22560 31894 22612 31900
rect 22572 31346 22600 31894
rect 22664 31890 22692 35414
rect 22744 35012 22796 35018
rect 22744 34954 22796 34960
rect 22756 34746 22784 34954
rect 22744 34740 22796 34746
rect 22744 34682 22796 34688
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 22560 31340 22612 31346
rect 22560 31282 22612 31288
rect 22560 30252 22612 30258
rect 22560 30194 22612 30200
rect 22572 29646 22600 30194
rect 22756 29646 22784 34682
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 22848 32026 22876 32370
rect 22836 32020 22888 32026
rect 22836 31962 22888 31968
rect 22836 31884 22888 31890
rect 22836 31826 22888 31832
rect 22560 29640 22612 29646
rect 22560 29582 22612 29588
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 22572 29238 22600 29582
rect 22560 29232 22612 29238
rect 22560 29174 22612 29180
rect 22848 29034 22876 31826
rect 22836 29028 22888 29034
rect 22836 28970 22888 28976
rect 22744 28620 22796 28626
rect 22744 28562 22796 28568
rect 22480 28478 22692 28506
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22480 26586 22508 26930
rect 22560 26784 22612 26790
rect 22560 26726 22612 26732
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 22468 26444 22520 26450
rect 22468 26386 22520 26392
rect 22480 26353 22508 26386
rect 22572 26382 22600 26726
rect 22560 26376 22612 26382
rect 22466 26344 22522 26353
rect 22560 26318 22612 26324
rect 22466 26279 22522 26288
rect 22572 23730 22600 26318
rect 22664 25294 22692 28478
rect 22756 28422 22784 28562
rect 22744 28416 22796 28422
rect 22744 28358 22796 28364
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22664 23798 22692 24754
rect 22652 23792 22704 23798
rect 22650 23760 22652 23769
rect 22704 23760 22706 23769
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22560 23724 22612 23730
rect 22650 23695 22706 23704
rect 22560 23666 22612 23672
rect 22756 23118 22784 28358
rect 22836 25696 22888 25702
rect 22836 25638 22888 25644
rect 22848 24818 22876 25638
rect 22940 24818 22968 36518
rect 23032 35018 23060 38966
rect 23296 38956 23348 38962
rect 23296 38898 23348 38904
rect 23308 36786 23336 38898
rect 23296 36780 23348 36786
rect 23296 36722 23348 36728
rect 23296 36032 23348 36038
rect 23296 35974 23348 35980
rect 23308 35630 23336 35974
rect 23400 35698 23428 39782
rect 23492 39370 23520 40326
rect 23480 39364 23532 39370
rect 23480 39306 23532 39312
rect 23388 35692 23440 35698
rect 23388 35634 23440 35640
rect 23296 35624 23348 35630
rect 23296 35566 23348 35572
rect 23020 35012 23072 35018
rect 23020 34954 23072 34960
rect 23032 31414 23060 34954
rect 23112 34672 23164 34678
rect 23112 34614 23164 34620
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 23032 31142 23060 31350
rect 23020 31136 23072 31142
rect 23020 31078 23072 31084
rect 23020 29504 23072 29510
rect 23020 29446 23072 29452
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22928 24812 22980 24818
rect 22928 24754 22980 24760
rect 22744 23112 22796 23118
rect 22744 23054 22796 23060
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22204 21706 22232 21966
rect 22112 21678 22232 21706
rect 22112 21350 22140 21678
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22112 20942 22140 21286
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22112 20534 22140 20878
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22008 19712 22060 19718
rect 22008 19654 22060 19660
rect 22020 19310 22048 19654
rect 22112 19446 22140 19994
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22204 19378 22232 19790
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22008 19304 22060 19310
rect 22008 19246 22060 19252
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 22020 18358 22048 18906
rect 22008 18352 22060 18358
rect 22008 18294 22060 18300
rect 22204 18086 22232 19110
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22100 17264 22152 17270
rect 22100 17206 22152 17212
rect 22008 15632 22060 15638
rect 22008 15574 22060 15580
rect 22020 15434 22048 15574
rect 22008 15428 22060 15434
rect 22008 15370 22060 15376
rect 22112 13938 22140 17206
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22204 15026 22232 15438
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 22204 14822 22232 14962
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22204 13530 22232 14758
rect 22192 13524 22244 13530
rect 22192 13466 22244 13472
rect 22192 12436 22244 12442
rect 22192 12378 22244 12384
rect 22204 11558 22232 12378
rect 22192 11552 22244 11558
rect 22192 11494 22244 11500
rect 22296 10742 22324 22918
rect 22468 22160 22520 22166
rect 22468 22102 22520 22108
rect 22928 22160 22980 22166
rect 22928 22102 22980 22108
rect 22480 21962 22508 22102
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22652 21888 22704 21894
rect 22652 21830 22704 21836
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22572 20942 22600 21490
rect 22664 21486 22692 21830
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22756 21128 22784 21966
rect 22836 21140 22888 21146
rect 22756 21100 22836 21128
rect 22836 21082 22888 21088
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22940 20874 22968 22102
rect 23032 22094 23060 29446
rect 23124 23322 23152 34614
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 23216 30938 23244 31282
rect 23204 30932 23256 30938
rect 23204 30874 23256 30880
rect 23216 30258 23244 30874
rect 23204 30252 23256 30258
rect 23204 30194 23256 30200
rect 23480 30184 23532 30190
rect 23480 30126 23532 30132
rect 23492 29306 23520 30126
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23296 29232 23348 29238
rect 23296 29174 23348 29180
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23216 28370 23244 28970
rect 23308 28558 23336 29174
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 23216 28342 23336 28370
rect 23204 23520 23256 23526
rect 23204 23462 23256 23468
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 23124 22778 23152 23122
rect 23216 23118 23244 23462
rect 23204 23112 23256 23118
rect 23204 23054 23256 23060
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23308 22710 23336 28342
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23400 22166 23428 23054
rect 23388 22160 23440 22166
rect 23388 22102 23440 22108
rect 23032 22066 23152 22094
rect 23124 21894 23152 22066
rect 23112 21888 23164 21894
rect 23112 21830 23164 21836
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23112 21616 23164 21622
rect 23112 21558 23164 21564
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 23032 20942 23060 21286
rect 23124 21146 23152 21558
rect 23112 21140 23164 21146
rect 23112 21082 23164 21088
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 22940 20058 22968 20810
rect 23032 20466 23060 20878
rect 23308 20466 23336 21830
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 22928 20052 22980 20058
rect 22928 19994 22980 20000
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 22744 19372 22796 19378
rect 22744 19314 22796 19320
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 22376 18828 22428 18834
rect 22376 18770 22428 18776
rect 22388 17270 22416 18770
rect 22376 17264 22428 17270
rect 22376 17206 22428 17212
rect 22480 16454 22508 19110
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22388 14006 22416 15370
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22388 11762 22416 12378
rect 22480 12102 22508 16390
rect 22664 15910 22692 16390
rect 22756 16114 22784 19314
rect 23492 18290 23520 19450
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22940 16114 22968 17070
rect 22744 16108 22796 16114
rect 22744 16050 22796 16056
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 22652 15904 22704 15910
rect 22652 15846 22704 15852
rect 22664 15570 22692 15846
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22664 15026 22692 15506
rect 22756 15076 22784 16050
rect 22940 15706 22968 16050
rect 23296 16040 23348 16046
rect 23296 15982 23348 15988
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 22836 15088 22888 15094
rect 22756 15048 22836 15076
rect 22652 15020 22704 15026
rect 22652 14962 22704 14968
rect 22560 14816 22612 14822
rect 22560 14758 22612 14764
rect 22572 14414 22600 14758
rect 22756 14482 22784 15048
rect 22836 15030 22888 15036
rect 23112 15088 23164 15094
rect 23112 15030 23164 15036
rect 22744 14476 22796 14482
rect 22744 14418 22796 14424
rect 23124 14414 23152 15030
rect 23308 15026 23336 15982
rect 23492 15706 23520 16050
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23204 14952 23256 14958
rect 23204 14894 23256 14900
rect 23308 14906 23336 14962
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 23124 13734 23152 14214
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 22926 13288 22982 13297
rect 22926 13223 22982 13232
rect 22940 12850 22968 13223
rect 23112 12912 23164 12918
rect 23112 12854 23164 12860
rect 22928 12844 22980 12850
rect 22928 12786 22980 12792
rect 23124 12434 23152 12854
rect 23032 12406 23152 12434
rect 22742 12200 22798 12209
rect 22742 12135 22798 12144
rect 22468 12096 22520 12102
rect 22468 12038 22520 12044
rect 22756 11762 22784 12135
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22284 10736 22336 10742
rect 22284 10678 22336 10684
rect 22296 10062 22324 10678
rect 22480 10674 22508 10950
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22572 10606 22600 11698
rect 22756 11626 22784 11698
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22928 11008 22980 11014
rect 22928 10950 22980 10956
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22940 9654 22968 10950
rect 22928 9648 22980 9654
rect 22928 9590 22980 9596
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 22204 6866 22232 9454
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22940 7886 22968 8230
rect 22928 7880 22980 7886
rect 22928 7822 22980 7828
rect 22560 7812 22612 7818
rect 22560 7754 22612 7760
rect 22572 7410 22600 7754
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 21916 6452 21968 6458
rect 21916 6394 21968 6400
rect 22572 6390 22600 7346
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21364 5228 21416 5234
rect 21364 5170 21416 5176
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 21100 3738 21128 5102
rect 21180 4616 21232 4622
rect 21180 4558 21232 4564
rect 21088 3732 21140 3738
rect 21088 3674 21140 3680
rect 21086 3224 21142 3233
rect 21086 3159 21088 3168
rect 21140 3159 21142 3168
rect 21088 3130 21140 3136
rect 20996 2508 21048 2514
rect 20996 2450 21048 2456
rect 21088 1760 21140 1766
rect 21088 1702 21140 1708
rect 21100 800 21128 1702
rect 21192 800 21220 4558
rect 21376 4010 21404 5170
rect 21364 4004 21416 4010
rect 21364 3946 21416 3952
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 21284 2446 21312 3130
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21284 1766 21312 2382
rect 21272 1760 21324 1766
rect 21272 1702 21324 1708
rect 21376 800 21404 2994
rect 21468 800 21496 3538
rect 21652 3534 21680 5510
rect 21836 5370 21864 6190
rect 22192 5568 22244 5574
rect 22192 5510 22244 5516
rect 22652 5568 22704 5574
rect 22652 5510 22704 5516
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21652 800 21680 3470
rect 21744 800 21772 4966
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 21914 3768 21970 3777
rect 21914 3703 21916 3712
rect 21968 3703 21970 3712
rect 21916 3674 21968 3680
rect 21916 1760 21968 1766
rect 21916 1702 21968 1708
rect 21928 800 21956 1702
rect 22020 800 22048 4694
rect 22112 3058 22140 5034
rect 22204 3126 22232 5510
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22284 4616 22336 4622
rect 22284 4558 22336 4564
rect 22192 3120 22244 3126
rect 22192 3062 22244 3068
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22112 2774 22140 2994
rect 22112 2746 22232 2774
rect 22204 800 22232 2746
rect 22296 800 22324 4558
rect 22376 4548 22428 4554
rect 22376 4490 22428 4496
rect 22388 2854 22416 4490
rect 22468 4004 22520 4010
rect 22468 3946 22520 3952
rect 22376 2848 22428 2854
rect 22376 2790 22428 2796
rect 22480 2446 22508 3946
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22480 800 22508 2382
rect 22572 800 22600 4966
rect 22664 3194 22692 5510
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22652 3188 22704 3194
rect 22652 3130 22704 3136
rect 22848 3058 22876 3334
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22848 2774 22876 2994
rect 22756 2746 22876 2774
rect 22652 2576 22704 2582
rect 22652 2518 22704 2524
rect 22664 2106 22692 2518
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 22756 800 22784 2746
rect 22940 898 22968 3878
rect 23032 3194 23060 12406
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 23124 11558 23152 11698
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23124 9450 23152 11086
rect 23112 9444 23164 9450
rect 23112 9386 23164 9392
rect 23124 7970 23152 9386
rect 23216 8090 23244 14894
rect 23308 14878 23428 14906
rect 23308 14822 23336 14878
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23400 14414 23428 14878
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 23124 7942 23244 7970
rect 23216 7886 23244 7942
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23216 7410 23244 7822
rect 23308 7546 23336 13806
rect 23492 13734 23520 14758
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 23492 11762 23520 12038
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23400 11150 23428 11698
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23400 10674 23428 10950
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23584 10538 23612 56102
rect 27620 55752 27672 55758
rect 27618 55720 27620 55729
rect 27672 55720 27674 55729
rect 27618 55655 27674 55664
rect 23940 55412 23992 55418
rect 23940 55354 23992 55360
rect 23664 40384 23716 40390
rect 23664 40326 23716 40332
rect 23676 40186 23704 40326
rect 23664 40180 23716 40186
rect 23664 40122 23716 40128
rect 23664 37936 23716 37942
rect 23664 37878 23716 37884
rect 23676 34678 23704 37878
rect 23848 34944 23900 34950
rect 23848 34886 23900 34892
rect 23664 34672 23716 34678
rect 23664 34614 23716 34620
rect 23676 32026 23704 34614
rect 23860 33930 23888 34886
rect 23848 33924 23900 33930
rect 23848 33866 23900 33872
rect 23860 33318 23888 33866
rect 23848 33312 23900 33318
rect 23848 33254 23900 33260
rect 23756 32496 23808 32502
rect 23756 32438 23808 32444
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 23676 30258 23704 31282
rect 23768 30326 23796 32438
rect 23860 32298 23888 33254
rect 23848 32292 23900 32298
rect 23848 32234 23900 32240
rect 23848 32020 23900 32026
rect 23848 31962 23900 31968
rect 23860 30938 23888 31962
rect 23848 30932 23900 30938
rect 23848 30874 23900 30880
rect 23848 30592 23900 30598
rect 23848 30534 23900 30540
rect 23756 30320 23808 30326
rect 23756 30262 23808 30268
rect 23664 30252 23716 30258
rect 23664 30194 23716 30200
rect 23676 29170 23704 30194
rect 23754 29200 23810 29209
rect 23664 29164 23716 29170
rect 23754 29135 23810 29144
rect 23664 29106 23716 29112
rect 23768 29102 23796 29135
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23860 28994 23888 30534
rect 23676 28966 23888 28994
rect 23676 24954 23704 28966
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23768 28150 23796 28358
rect 23756 28144 23808 28150
rect 23756 28086 23808 28092
rect 23952 26908 23980 55354
rect 29196 45554 29224 56306
rect 30024 55622 30052 56306
rect 30852 56166 30880 56306
rect 31772 56166 31800 57462
rect 32128 57452 32180 57458
rect 32128 57394 32180 57400
rect 33140 57452 33192 57458
rect 33140 57394 33192 57400
rect 34704 57452 34756 57458
rect 34704 57394 34756 57400
rect 37832 57452 37884 57458
rect 37832 57394 37884 57400
rect 39856 57452 39908 57458
rect 39856 57394 39908 57400
rect 42524 57452 42576 57458
rect 42524 57394 42576 57400
rect 44088 57452 44140 57458
rect 44088 57394 44140 57400
rect 44180 57452 44232 57458
rect 44180 57394 44232 57400
rect 32140 56506 32168 57394
rect 33152 56506 33180 57394
rect 34716 56506 34744 57394
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 37844 56506 37872 57394
rect 32128 56500 32180 56506
rect 32128 56442 32180 56448
rect 33140 56500 33192 56506
rect 33140 56442 33192 56448
rect 34704 56500 34756 56506
rect 34704 56442 34756 56448
rect 37832 56500 37884 56506
rect 37832 56442 37884 56448
rect 32128 56364 32180 56370
rect 32128 56306 32180 56312
rect 33600 56364 33652 56370
rect 33600 56306 33652 56312
rect 35808 56364 35860 56370
rect 35808 56306 35860 56312
rect 30840 56160 30892 56166
rect 30840 56102 30892 56108
rect 31760 56160 31812 56166
rect 31760 56102 31812 56108
rect 30012 55616 30064 55622
rect 30012 55558 30064 55564
rect 29012 45526 29224 45554
rect 24400 41472 24452 41478
rect 24400 41414 24452 41420
rect 29012 41414 29040 45526
rect 30024 43761 30052 55558
rect 30010 43752 30066 43761
rect 30010 43687 30066 43696
rect 30852 41414 30880 56102
rect 32140 42401 32168 56306
rect 33612 44849 33640 56306
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 33598 44840 33654 44849
rect 33598 44775 33654 44784
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 32126 42392 32182 42401
rect 32126 42327 32182 42336
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 24216 37664 24268 37670
rect 24216 37606 24268 37612
rect 24228 37194 24256 37606
rect 24216 37188 24268 37194
rect 24216 37130 24268 37136
rect 24228 36854 24256 37130
rect 24216 36848 24268 36854
rect 24216 36790 24268 36796
rect 24216 35692 24268 35698
rect 24216 35634 24268 35640
rect 24308 35692 24360 35698
rect 24308 35634 24360 35640
rect 24228 35154 24256 35634
rect 24216 35148 24268 35154
rect 24216 35090 24268 35096
rect 24216 34944 24268 34950
rect 24216 34886 24268 34892
rect 24124 33992 24176 33998
rect 24124 33934 24176 33940
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 24044 32434 24072 32710
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 23768 26880 23980 26908
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23676 14074 23704 14486
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23480 9580 23532 9586
rect 23480 9522 23532 9528
rect 23492 8974 23520 9522
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23204 7404 23256 7410
rect 23204 7346 23256 7352
rect 23216 6322 23244 7346
rect 23480 7200 23532 7206
rect 23584 7188 23612 9590
rect 23532 7160 23612 7188
rect 23480 7142 23532 7148
rect 23492 6934 23520 7142
rect 23480 6928 23532 6934
rect 23480 6870 23532 6876
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 23020 3188 23072 3194
rect 23020 3130 23072 3136
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 22848 870 22968 898
rect 22848 800 22876 870
rect 23032 800 23060 2246
rect 23124 800 23152 3878
rect 23216 2990 23244 5510
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23204 2984 23256 2990
rect 23204 2926 23256 2932
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23308 800 23336 2382
rect 23400 800 23428 3878
rect 23492 3466 23520 4966
rect 23584 4622 23612 6598
rect 23676 6458 23704 13806
rect 23768 12918 23796 26880
rect 24044 22094 24072 32370
rect 24136 32026 24164 33934
rect 24228 32434 24256 34886
rect 24320 34202 24348 35634
rect 24412 34218 24440 41414
rect 29012 41386 29316 41414
rect 24768 41200 24820 41206
rect 24768 41142 24820 41148
rect 24584 38956 24636 38962
rect 24584 38898 24636 38904
rect 24596 38350 24624 38898
rect 24780 38758 24808 41142
rect 26608 40928 26660 40934
rect 26608 40870 26660 40876
rect 25044 39976 25096 39982
rect 25044 39918 25096 39924
rect 25056 39438 25084 39918
rect 25044 39432 25096 39438
rect 25044 39374 25096 39380
rect 24952 39024 25004 39030
rect 24952 38966 25004 38972
rect 24768 38752 24820 38758
rect 24768 38694 24820 38700
rect 24964 38486 24992 38966
rect 24952 38480 25004 38486
rect 24952 38422 25004 38428
rect 24584 38344 24636 38350
rect 24584 38286 24636 38292
rect 24768 38344 24820 38350
rect 24768 38286 24820 38292
rect 24492 35012 24544 35018
rect 24492 34954 24544 34960
rect 24504 34746 24532 34954
rect 24492 34740 24544 34746
rect 24492 34682 24544 34688
rect 24412 34202 24532 34218
rect 24308 34196 24360 34202
rect 24308 34138 24360 34144
rect 24412 34196 24544 34202
rect 24412 34190 24492 34196
rect 24412 33998 24440 34190
rect 24492 34138 24544 34144
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24596 33522 24624 38286
rect 24676 38208 24728 38214
rect 24676 38150 24728 38156
rect 24584 33516 24636 33522
rect 24584 33458 24636 33464
rect 24596 32978 24624 33458
rect 24584 32972 24636 32978
rect 24584 32914 24636 32920
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 24124 32020 24176 32026
rect 24124 31962 24176 31968
rect 24228 31482 24256 32370
rect 24216 31476 24268 31482
rect 24216 31418 24268 31424
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 24216 30252 24268 30258
rect 24216 30194 24268 30200
rect 24124 29708 24176 29714
rect 24124 29650 24176 29656
rect 24136 29034 24164 29650
rect 24228 29170 24256 30194
rect 24412 30122 24440 30670
rect 24596 30258 24624 32914
rect 24688 31686 24716 38150
rect 24780 37466 24808 38286
rect 24768 37460 24820 37466
rect 24768 37402 24820 37408
rect 24964 37346 24992 38422
rect 25056 37942 25084 39374
rect 25412 38956 25464 38962
rect 25412 38898 25464 38904
rect 25596 38956 25648 38962
rect 25596 38898 25648 38904
rect 25228 38752 25280 38758
rect 25228 38694 25280 38700
rect 25044 37936 25096 37942
rect 25044 37878 25096 37884
rect 24872 37318 24992 37346
rect 24768 36236 24820 36242
rect 24768 36178 24820 36184
rect 24780 35290 24808 36178
rect 24768 35284 24820 35290
rect 24768 35226 24820 35232
rect 24872 34610 24900 37318
rect 24952 37188 25004 37194
rect 24952 37130 25004 37136
rect 24964 34950 24992 37130
rect 25056 36582 25084 37878
rect 25044 36576 25096 36582
rect 25044 36518 25096 36524
rect 25056 35766 25084 36518
rect 25044 35760 25096 35766
rect 25044 35702 25096 35708
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 25136 34604 25188 34610
rect 25136 34546 25188 34552
rect 24872 34490 24900 34546
rect 24780 34462 24900 34490
rect 24780 33998 24808 34462
rect 25148 33998 25176 34546
rect 24768 33992 24820 33998
rect 24768 33934 24820 33940
rect 25136 33992 25188 33998
rect 25136 33934 25188 33940
rect 24780 33590 24808 33934
rect 24768 33584 24820 33590
rect 24768 33526 24820 33532
rect 24676 31680 24728 31686
rect 24676 31622 24728 31628
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24400 30116 24452 30122
rect 24400 30058 24452 30064
rect 24412 29209 24440 30058
rect 24688 29782 24716 31622
rect 24780 30802 24808 33526
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24872 32570 24900 33458
rect 25240 33114 25268 38694
rect 25320 38208 25372 38214
rect 25320 38150 25372 38156
rect 25332 37874 25360 38150
rect 25424 38010 25452 38898
rect 25608 38758 25636 38898
rect 25596 38752 25648 38758
rect 25596 38694 25648 38700
rect 25964 38752 26016 38758
rect 25964 38694 26016 38700
rect 25976 38350 26004 38694
rect 25688 38344 25740 38350
rect 25688 38286 25740 38292
rect 25964 38344 26016 38350
rect 25964 38286 26016 38292
rect 25412 38004 25464 38010
rect 25412 37946 25464 37952
rect 25700 37942 25728 38286
rect 26332 38208 26384 38214
rect 26332 38150 26384 38156
rect 25688 37936 25740 37942
rect 25688 37878 25740 37884
rect 26148 37936 26200 37942
rect 26148 37878 26200 37884
rect 25320 37868 25372 37874
rect 25320 37810 25372 37816
rect 26160 37194 26188 37878
rect 26344 37874 26372 38150
rect 26332 37868 26384 37874
rect 26332 37810 26384 37816
rect 26148 37188 26200 37194
rect 26148 37130 26200 37136
rect 25780 35284 25832 35290
rect 25780 35226 25832 35232
rect 25792 34678 25820 35226
rect 25964 34944 26016 34950
rect 25964 34886 26016 34892
rect 26240 34944 26292 34950
rect 26240 34886 26292 34892
rect 25976 34678 26004 34886
rect 25780 34672 25832 34678
rect 25780 34614 25832 34620
rect 25964 34672 26016 34678
rect 25964 34614 26016 34620
rect 26252 34066 26280 34886
rect 26240 34060 26292 34066
rect 26240 34002 26292 34008
rect 25504 33516 25556 33522
rect 25504 33458 25556 33464
rect 25516 33318 25544 33458
rect 25320 33312 25372 33318
rect 25320 33254 25372 33260
rect 25504 33312 25556 33318
rect 25504 33254 25556 33260
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 25332 32502 25360 33254
rect 25412 32564 25464 32570
rect 25412 32506 25464 32512
rect 25320 32496 25372 32502
rect 25320 32438 25372 32444
rect 25044 32224 25096 32230
rect 25044 32166 25096 32172
rect 24860 31136 24912 31142
rect 24860 31078 24912 31084
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 24872 30666 24900 31078
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24952 30116 25004 30122
rect 24952 30058 25004 30064
rect 24964 29850 24992 30058
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 24676 29776 24728 29782
rect 24676 29718 24728 29724
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24596 29306 24624 29446
rect 24584 29300 24636 29306
rect 24584 29242 24636 29248
rect 24676 29232 24728 29238
rect 24398 29200 24454 29209
rect 24216 29164 24268 29170
rect 24676 29174 24728 29180
rect 24398 29135 24454 29144
rect 24216 29106 24268 29112
rect 24124 29028 24176 29034
rect 24124 28970 24176 28976
rect 24124 28552 24176 28558
rect 24124 28494 24176 28500
rect 23860 22066 24072 22094
rect 23860 13394 23888 22066
rect 23940 20868 23992 20874
rect 23940 20810 23992 20816
rect 23952 19514 23980 20810
rect 23940 19508 23992 19514
rect 23940 19450 23992 19456
rect 24136 17678 24164 28494
rect 24412 27538 24440 29135
rect 24688 29016 24716 29174
rect 24952 29164 25004 29170
rect 24952 29106 25004 29112
rect 24596 28988 24716 29016
rect 24596 28422 24624 28988
rect 24964 28762 24992 29106
rect 24952 28756 25004 28762
rect 24952 28698 25004 28704
rect 24584 28416 24636 28422
rect 24584 28358 24636 28364
rect 24400 27532 24452 27538
rect 24400 27474 24452 27480
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24688 26994 24716 27270
rect 24676 26988 24728 26994
rect 24676 26930 24728 26936
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24320 18630 24348 26522
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24596 25906 24624 26318
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24688 25498 24716 26930
rect 24768 26920 24820 26926
rect 24768 26862 24820 26868
rect 24780 25498 24808 26862
rect 24872 26518 24900 27270
rect 24860 26512 24912 26518
rect 24860 26454 24912 26460
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24676 25492 24728 25498
rect 24676 25434 24728 25440
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24688 23662 24716 24822
rect 24964 24818 24992 25842
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24952 24336 25004 24342
rect 24952 24278 25004 24284
rect 25056 24290 25084 32166
rect 25136 30592 25188 30598
rect 25136 30534 25188 30540
rect 25148 30326 25176 30534
rect 25136 30320 25188 30326
rect 25136 30262 25188 30268
rect 25136 28484 25188 28490
rect 25136 28426 25188 28432
rect 25148 27946 25176 28426
rect 25136 27940 25188 27946
rect 25136 27882 25188 27888
rect 25136 26852 25188 26858
rect 25136 26794 25188 26800
rect 25148 26450 25176 26794
rect 25136 26444 25188 26450
rect 25136 26386 25188 26392
rect 25148 25974 25176 26386
rect 25136 25968 25188 25974
rect 25136 25910 25188 25916
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25148 24410 25176 24754
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 24964 23866 24992 24278
rect 25056 24262 25176 24290
rect 24768 23860 24820 23866
rect 24768 23802 24820 23808
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 24780 23746 24808 23802
rect 24780 23730 24992 23746
rect 24780 23724 25004 23730
rect 24780 23718 24952 23724
rect 24952 23666 25004 23672
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 24688 23118 24716 23598
rect 24676 23112 24728 23118
rect 24676 23054 24728 23060
rect 25044 22636 25096 22642
rect 25044 22578 25096 22584
rect 25056 21622 25084 22578
rect 25044 21616 25096 21622
rect 25044 21558 25096 21564
rect 24676 21548 24728 21554
rect 24676 21490 24728 21496
rect 24688 21350 24716 21490
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24400 20800 24452 20806
rect 24400 20742 24452 20748
rect 24412 20262 24440 20742
rect 24400 20256 24452 20262
rect 24400 20198 24452 20204
rect 24412 19378 24440 20198
rect 24584 19780 24636 19786
rect 24584 19722 24636 19728
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24596 18902 24624 19722
rect 24584 18896 24636 18902
rect 24584 18838 24636 18844
rect 24308 18624 24360 18630
rect 24308 18566 24360 18572
rect 24216 18352 24268 18358
rect 24216 18294 24268 18300
rect 24124 17672 24176 17678
rect 24124 17614 24176 17620
rect 24228 17202 24256 18294
rect 24688 18290 24716 21286
rect 25056 20874 25084 21558
rect 25044 20868 25096 20874
rect 25044 20810 25096 20816
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24780 18358 24808 19382
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 24964 18290 24992 19246
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24964 17202 24992 18226
rect 24216 17196 24268 17202
rect 24216 17138 24268 17144
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24032 17128 24084 17134
rect 24032 17070 24084 17076
rect 24044 16114 24072 17070
rect 25044 16992 25096 16998
rect 25044 16934 25096 16940
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24492 16720 24544 16726
rect 24492 16662 24544 16668
rect 24032 16108 24084 16114
rect 24032 16050 24084 16056
rect 24030 15600 24086 15609
rect 24030 15535 24086 15544
rect 24044 14822 24072 15535
rect 24308 15496 24360 15502
rect 24308 15438 24360 15444
rect 24320 14822 24348 15438
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24032 14816 24084 14822
rect 24032 14758 24084 14764
rect 24216 14816 24268 14822
rect 24216 14758 24268 14764
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24228 14618 24256 14758
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23952 13841 23980 14010
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 23938 13832 23994 13841
rect 23938 13767 23994 13776
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23860 12986 23888 13330
rect 24044 12986 24072 13874
rect 23848 12980 23900 12986
rect 23848 12922 23900 12928
rect 24032 12980 24084 12986
rect 24032 12922 24084 12928
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23756 11144 23808 11150
rect 23756 11086 23808 11092
rect 23768 10810 23796 11086
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 24032 8900 24084 8906
rect 24032 8842 24084 8848
rect 23848 7472 23900 7478
rect 23848 7414 23900 7420
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23768 5914 23796 6734
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23860 5642 23888 7414
rect 24044 6458 24072 8842
rect 24136 8022 24164 13874
rect 24412 13190 24440 14962
rect 24504 14618 24532 16662
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24400 13184 24452 13190
rect 24400 13126 24452 13132
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24124 8016 24176 8022
rect 24124 7958 24176 7964
rect 24228 7546 24256 12922
rect 24596 12306 24624 16730
rect 25056 14958 25084 16934
rect 25044 14952 25096 14958
rect 25044 14894 25096 14900
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24872 12434 24900 14350
rect 25148 14074 25176 24262
rect 25240 24138 25268 25230
rect 25228 24132 25280 24138
rect 25228 24074 25280 24080
rect 25240 22778 25268 24074
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25332 23050 25360 23734
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25228 22772 25280 22778
rect 25228 22714 25280 22720
rect 25320 19712 25372 19718
rect 25320 19654 25372 19660
rect 25332 19446 25360 19654
rect 25320 19440 25372 19446
rect 25320 19382 25372 19388
rect 25424 16726 25452 32506
rect 25516 29753 25544 33254
rect 25780 33108 25832 33114
rect 25780 33050 25832 33056
rect 25688 31136 25740 31142
rect 25688 31078 25740 31084
rect 25700 30258 25728 31078
rect 25688 30252 25740 30258
rect 25688 30194 25740 30200
rect 25502 29744 25558 29753
rect 25502 29679 25558 29688
rect 25516 29306 25544 29679
rect 25596 29572 25648 29578
rect 25596 29514 25648 29520
rect 25504 29300 25556 29306
rect 25504 29242 25556 29248
rect 25608 29034 25636 29514
rect 25596 29028 25648 29034
rect 25596 28970 25648 28976
rect 25792 28762 25820 33050
rect 26240 30660 26292 30666
rect 26240 30602 26292 30608
rect 26252 30326 26280 30602
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 25872 30048 25924 30054
rect 25872 29990 25924 29996
rect 25884 28966 25912 29990
rect 26344 29850 26372 37810
rect 26424 35488 26476 35494
rect 26424 35430 26476 35436
rect 26436 35086 26464 35430
rect 26424 35080 26476 35086
rect 26424 35022 26476 35028
rect 26332 29844 26384 29850
rect 26332 29786 26384 29792
rect 26424 29504 26476 29510
rect 26424 29446 26476 29452
rect 26148 29164 26200 29170
rect 26148 29106 26200 29112
rect 26160 29073 26188 29106
rect 26146 29064 26202 29073
rect 26146 28999 26148 29008
rect 26200 28999 26202 29008
rect 26148 28970 26200 28976
rect 25872 28960 25924 28966
rect 25872 28902 25924 28908
rect 25780 28756 25832 28762
rect 25780 28698 25832 28704
rect 25608 27130 25820 27146
rect 25596 27124 25820 27130
rect 25648 27118 25820 27124
rect 25596 27066 25648 27072
rect 25792 27062 25820 27118
rect 25780 27056 25832 27062
rect 25780 26998 25832 27004
rect 25884 26790 25912 28902
rect 26436 28082 26464 29446
rect 26620 28994 26648 40870
rect 27252 40520 27304 40526
rect 27252 40462 27304 40468
rect 27160 40452 27212 40458
rect 27160 40394 27212 40400
rect 27172 39098 27200 40394
rect 27264 39438 27292 40462
rect 28172 40384 28224 40390
rect 28172 40326 28224 40332
rect 28184 40118 28212 40326
rect 28172 40112 28224 40118
rect 28172 40054 28224 40060
rect 29184 40112 29236 40118
rect 29184 40054 29236 40060
rect 27620 39840 27672 39846
rect 27620 39782 27672 39788
rect 27252 39432 27304 39438
rect 27304 39392 27476 39420
rect 27252 39374 27304 39380
rect 27160 39092 27212 39098
rect 27160 39034 27212 39040
rect 27344 38344 27396 38350
rect 27344 38286 27396 38292
rect 27356 37670 27384 38286
rect 27448 37806 27476 39392
rect 27528 39364 27580 39370
rect 27528 39306 27580 39312
rect 27540 38554 27568 39306
rect 27632 38962 27660 39782
rect 27896 39092 27948 39098
rect 27896 39034 27948 39040
rect 27620 38956 27672 38962
rect 27620 38898 27672 38904
rect 27712 38888 27764 38894
rect 27712 38830 27764 38836
rect 27528 38548 27580 38554
rect 27528 38490 27580 38496
rect 27436 37800 27488 37806
rect 27436 37742 27488 37748
rect 27344 37664 27396 37670
rect 27344 37606 27396 37612
rect 27068 36032 27120 36038
rect 27068 35974 27120 35980
rect 27080 35834 27108 35974
rect 27068 35828 27120 35834
rect 27068 35770 27120 35776
rect 27080 35222 27108 35770
rect 27068 35216 27120 35222
rect 27068 35158 27120 35164
rect 27080 34746 27108 35158
rect 27068 34740 27120 34746
rect 27068 34682 27120 34688
rect 27080 34066 27108 34682
rect 27068 34060 27120 34066
rect 27068 34002 27120 34008
rect 27356 33998 27384 37606
rect 27448 35698 27476 37742
rect 27528 36576 27580 36582
rect 27528 36518 27580 36524
rect 27540 36174 27568 36518
rect 27528 36168 27580 36174
rect 27528 36110 27580 36116
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27620 35692 27672 35698
rect 27620 35634 27672 35640
rect 27528 35488 27580 35494
rect 27528 35430 27580 35436
rect 27540 35154 27568 35430
rect 27632 35290 27660 35634
rect 27620 35284 27672 35290
rect 27620 35226 27672 35232
rect 27528 35148 27580 35154
rect 27528 35090 27580 35096
rect 27620 35148 27672 35154
rect 27620 35090 27672 35096
rect 27632 34626 27660 35090
rect 27724 35086 27752 38830
rect 27908 38486 27936 39034
rect 28080 38956 28132 38962
rect 28080 38898 28132 38904
rect 27896 38480 27948 38486
rect 27896 38422 27948 38428
rect 28092 38350 28120 38898
rect 28080 38344 28132 38350
rect 28080 38286 28132 38292
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 27804 35760 27856 35766
rect 27804 35702 27856 35708
rect 27712 35080 27764 35086
rect 27712 35022 27764 35028
rect 27724 34746 27752 35022
rect 27712 34740 27764 34746
rect 27712 34682 27764 34688
rect 27816 34626 27844 35702
rect 27632 34598 27844 34626
rect 26700 33992 26752 33998
rect 26698 33960 26700 33969
rect 27344 33992 27396 33998
rect 26752 33960 26754 33969
rect 27344 33934 27396 33940
rect 26698 33895 26754 33904
rect 27632 33862 27660 34598
rect 27712 33992 27764 33998
rect 27712 33934 27764 33940
rect 27252 33856 27304 33862
rect 27252 33798 27304 33804
rect 27620 33856 27672 33862
rect 27620 33798 27672 33804
rect 27264 33590 27292 33798
rect 27252 33584 27304 33590
rect 27252 33526 27304 33532
rect 27160 33448 27212 33454
rect 27160 33390 27212 33396
rect 27172 32366 27200 33390
rect 27724 33114 27752 33934
rect 27712 33108 27764 33114
rect 27712 33050 27764 33056
rect 27160 32360 27212 32366
rect 27160 32302 27212 32308
rect 27172 31890 27200 32302
rect 27160 31884 27212 31890
rect 27160 31826 27212 31832
rect 27172 31754 27200 31826
rect 27080 31726 27200 31754
rect 27080 30734 27108 31726
rect 27908 30938 27936 36246
rect 28184 32434 28212 40054
rect 28816 39296 28868 39302
rect 28816 39238 28868 39244
rect 29000 39296 29052 39302
rect 29000 39238 29052 39244
rect 28828 38282 28856 39238
rect 29012 38962 29040 39238
rect 29000 38956 29052 38962
rect 29000 38898 29052 38904
rect 28816 38276 28868 38282
rect 28816 38218 28868 38224
rect 28724 36304 28776 36310
rect 28724 36246 28776 36252
rect 28448 36236 28500 36242
rect 28448 36178 28500 36184
rect 28460 35766 28488 36178
rect 28736 36174 28764 36246
rect 28724 36168 28776 36174
rect 28724 36110 28776 36116
rect 28448 35760 28500 35766
rect 28448 35702 28500 35708
rect 28448 35488 28500 35494
rect 28448 35430 28500 35436
rect 28460 35086 28488 35430
rect 28448 35080 28500 35086
rect 28448 35022 28500 35028
rect 28460 32502 28488 35022
rect 28540 33312 28592 33318
rect 28540 33254 28592 33260
rect 28552 32910 28580 33254
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28552 32502 28580 32846
rect 28828 32570 28856 38218
rect 29012 36786 29040 38898
rect 29092 38752 29144 38758
rect 29092 38694 29144 38700
rect 29104 38418 29132 38694
rect 29092 38412 29144 38418
rect 29092 38354 29144 38360
rect 29104 37806 29132 38354
rect 29196 38350 29224 40054
rect 29184 38344 29236 38350
rect 29184 38286 29236 38292
rect 29196 38010 29224 38286
rect 29184 38004 29236 38010
rect 29184 37946 29236 37952
rect 29184 37868 29236 37874
rect 29184 37810 29236 37816
rect 29092 37800 29144 37806
rect 29092 37742 29144 37748
rect 29000 36780 29052 36786
rect 29000 36722 29052 36728
rect 29012 36378 29040 36722
rect 29000 36372 29052 36378
rect 29000 36314 29052 36320
rect 29196 36242 29224 37810
rect 29184 36236 29236 36242
rect 29184 36178 29236 36184
rect 28816 32564 28868 32570
rect 28816 32506 28868 32512
rect 28448 32496 28500 32502
rect 28448 32438 28500 32444
rect 28540 32496 28592 32502
rect 28540 32438 28592 32444
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 29012 32230 29040 32302
rect 29000 32224 29052 32230
rect 29000 32166 29052 32172
rect 29288 31754 29316 41386
rect 30668 41386 30880 41414
rect 30564 40044 30616 40050
rect 30564 39986 30616 39992
rect 30012 39840 30064 39846
rect 30012 39782 30064 39788
rect 29736 36372 29788 36378
rect 29736 36314 29788 36320
rect 29644 36032 29696 36038
rect 29564 35992 29644 36020
rect 29564 35018 29592 35992
rect 29644 35974 29696 35980
rect 29552 35012 29604 35018
rect 29552 34954 29604 34960
rect 29564 34610 29592 34954
rect 29644 34944 29696 34950
rect 29644 34886 29696 34892
rect 29552 34604 29604 34610
rect 29552 34546 29604 34552
rect 29564 33930 29592 34546
rect 29656 34542 29684 34886
rect 29644 34536 29696 34542
rect 29644 34478 29696 34484
rect 29552 33924 29604 33930
rect 29552 33866 29604 33872
rect 29564 32842 29592 33866
rect 29656 33522 29684 34478
rect 29644 33516 29696 33522
rect 29644 33458 29696 33464
rect 29656 33318 29684 33458
rect 29644 33312 29696 33318
rect 29644 33254 29696 33260
rect 29552 32836 29604 32842
rect 29552 32778 29604 32784
rect 28080 31748 28132 31754
rect 28080 31690 28132 31696
rect 29196 31726 29316 31754
rect 27896 30932 27948 30938
rect 27896 30874 27948 30880
rect 27908 30734 27936 30874
rect 27068 30728 27120 30734
rect 27068 30670 27120 30676
rect 27896 30728 27948 30734
rect 27896 30670 27948 30676
rect 27080 30258 27108 30670
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 27080 29714 27108 30194
rect 27068 29708 27120 29714
rect 27068 29650 27120 29656
rect 27526 29064 27582 29073
rect 27526 28999 27582 29008
rect 26620 28966 26740 28994
rect 26424 28076 26476 28082
rect 26424 28018 26476 28024
rect 26608 27940 26660 27946
rect 26608 27882 26660 27888
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 25608 26382 25636 26726
rect 25596 26376 25648 26382
rect 25596 26318 25648 26324
rect 26160 26314 26188 27338
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 25780 26240 25832 26246
rect 25780 26182 25832 26188
rect 25792 25906 25820 26182
rect 25780 25900 25832 25906
rect 25780 25842 25832 25848
rect 25872 25900 25924 25906
rect 25872 25842 25924 25848
rect 25884 24886 25912 25842
rect 26160 25294 26188 26250
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 25872 24880 25924 24886
rect 25872 24822 25924 24828
rect 25596 24744 25648 24750
rect 25596 24686 25648 24692
rect 25504 24200 25556 24206
rect 25504 24142 25556 24148
rect 25516 23186 25544 24142
rect 25608 24138 25636 24686
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25504 23180 25556 23186
rect 25504 23122 25556 23128
rect 25700 22438 25728 23666
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26160 23118 26188 23462
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 26424 21412 26476 21418
rect 26424 21354 26476 21360
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25792 20058 25820 20402
rect 25780 20052 25832 20058
rect 25780 19994 25832 20000
rect 26056 19848 26108 19854
rect 26056 19790 26108 19796
rect 26436 19836 26464 21354
rect 26516 19848 26568 19854
rect 26436 19808 26516 19836
rect 25594 19680 25650 19689
rect 25594 19615 25650 19624
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25516 18766 25544 19382
rect 25608 19378 25636 19615
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25688 19236 25740 19242
rect 25688 19178 25740 19184
rect 25700 18834 25728 19178
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25516 17882 25544 18702
rect 26068 18630 26096 19790
rect 26436 19514 26464 19808
rect 26516 19790 26568 19796
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26436 19174 26464 19450
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 26620 18766 26648 27882
rect 26712 27878 26740 28966
rect 26700 27872 26752 27878
rect 26700 27814 26752 27820
rect 27068 27872 27120 27878
rect 27068 27814 27120 27820
rect 26700 27464 26752 27470
rect 26752 27412 26832 27418
rect 26700 27406 26832 27412
rect 26712 27390 26832 27406
rect 26804 26382 26832 27390
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 26896 27130 26924 27338
rect 26884 27124 26936 27130
rect 26884 27066 26936 27072
rect 26792 26376 26844 26382
rect 26792 26318 26844 26324
rect 26804 25226 26832 26318
rect 27080 25974 27108 27814
rect 27160 27396 27212 27402
rect 27160 27338 27212 27344
rect 27068 25968 27120 25974
rect 27068 25910 27120 25916
rect 26792 25220 26844 25226
rect 26792 25162 26844 25168
rect 26804 24818 26832 25162
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26804 24206 26832 24754
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26884 24064 26936 24070
rect 26884 24006 26936 24012
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26332 18692 26384 18698
rect 26332 18634 26384 18640
rect 25780 18624 25832 18630
rect 25780 18566 25832 18572
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 25504 17876 25556 17882
rect 25504 17818 25556 17824
rect 25688 17604 25740 17610
rect 25688 17546 25740 17552
rect 25700 17338 25728 17546
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25792 17270 25820 18566
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25872 18216 25924 18222
rect 25872 18158 25924 18164
rect 25780 17264 25832 17270
rect 25780 17206 25832 17212
rect 25688 17196 25740 17202
rect 25688 17138 25740 17144
rect 25700 16726 25728 17138
rect 25412 16720 25464 16726
rect 25412 16662 25464 16668
rect 25688 16720 25740 16726
rect 25688 16662 25740 16668
rect 25884 15348 25912 18158
rect 25976 17241 26004 18226
rect 25962 17232 26018 17241
rect 25962 17167 26018 17176
rect 26240 17128 26292 17134
rect 26240 17070 26292 17076
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 25700 15320 25912 15348
rect 25504 14952 25556 14958
rect 25504 14894 25556 14900
rect 25516 14482 25544 14894
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25136 14068 25188 14074
rect 25136 14010 25188 14016
rect 25228 13252 25280 13258
rect 25228 13194 25280 13200
rect 24780 12406 24900 12434
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24780 9654 24808 12406
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11830 24992 12038
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24872 11218 24900 11630
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 24860 11212 24912 11218
rect 24860 11154 24912 11160
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24964 10538 24992 11086
rect 25056 10674 25084 11494
rect 25240 10674 25268 13194
rect 25596 12708 25648 12714
rect 25596 12650 25648 12656
rect 25320 12232 25372 12238
rect 25504 12232 25556 12238
rect 25320 12174 25372 12180
rect 25502 12200 25504 12209
rect 25556 12200 25558 12209
rect 25332 11898 25360 12174
rect 25502 12135 25558 12144
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25332 11150 25360 11834
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 24952 10532 25004 10538
rect 24952 10474 25004 10480
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24492 9104 24544 9110
rect 24492 9046 24544 9052
rect 24504 8838 24532 9046
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24504 8634 24532 8774
rect 24492 8628 24544 8634
rect 24492 8570 24544 8576
rect 24964 8566 24992 10474
rect 25056 9654 25084 10610
rect 25240 9738 25268 10610
rect 25332 10130 25360 11086
rect 25608 11082 25636 12650
rect 25596 11076 25648 11082
rect 25596 11018 25648 11024
rect 25608 10674 25636 11018
rect 25412 10668 25464 10674
rect 25412 10610 25464 10616
rect 25596 10668 25648 10674
rect 25596 10610 25648 10616
rect 25424 10266 25452 10610
rect 25412 10260 25464 10266
rect 25412 10202 25464 10208
rect 25608 10198 25636 10610
rect 25596 10192 25648 10198
rect 25596 10134 25648 10140
rect 25320 10124 25372 10130
rect 25320 10066 25372 10072
rect 25148 9710 25268 9738
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 24952 8560 25004 8566
rect 24952 8502 25004 8508
rect 25148 8498 25176 9710
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 25240 9178 25268 9522
rect 25424 9382 25452 9522
rect 25700 9450 25728 15320
rect 25780 12300 25832 12306
rect 25780 12242 25832 12248
rect 25792 10810 25820 12242
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 26068 9450 26096 16594
rect 26252 15706 26280 17070
rect 26344 16522 26372 18634
rect 26608 18352 26660 18358
rect 26608 18294 26660 18300
rect 26620 17882 26648 18294
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26240 15700 26292 15706
rect 26240 15642 26292 15648
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 26252 15162 26280 15438
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26344 14006 26372 15846
rect 26436 15502 26464 16050
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 26528 14482 26556 17614
rect 26620 16590 26648 17818
rect 26712 17202 26740 22646
rect 26896 22098 26924 24006
rect 26884 22092 26936 22098
rect 26884 22034 26936 22040
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 26974 19952 27030 19961
rect 26974 19887 27030 19896
rect 26884 19780 26936 19786
rect 26884 19722 26936 19728
rect 26896 18902 26924 19722
rect 26988 19514 27016 19887
rect 27080 19854 27108 20198
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 27172 19530 27200 27338
rect 27252 24064 27304 24070
rect 27252 24006 27304 24012
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 27080 19502 27200 19530
rect 26884 18896 26936 18902
rect 27080 18850 27108 19502
rect 27264 19446 27292 24006
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 27448 20874 27476 21966
rect 27436 20868 27488 20874
rect 27436 20810 27488 20816
rect 27448 20330 27476 20810
rect 27540 20466 27568 28999
rect 27908 28994 27936 30670
rect 27816 28966 27936 28994
rect 27620 27328 27672 27334
rect 27620 27270 27672 27276
rect 27632 26450 27660 27270
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 27724 26042 27752 26930
rect 27712 26036 27764 26042
rect 27712 25978 27764 25984
rect 27816 25430 27844 28966
rect 27988 27328 28040 27334
rect 27988 27270 28040 27276
rect 27804 25424 27856 25430
rect 27804 25366 27856 25372
rect 28000 25158 28028 27270
rect 27988 25152 28040 25158
rect 27988 25094 28040 25100
rect 27620 22976 27672 22982
rect 27620 22918 27672 22924
rect 27632 22710 27660 22918
rect 27620 22704 27672 22710
rect 27620 22646 27672 22652
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 27252 19440 27304 19446
rect 27252 19382 27304 19388
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27172 18902 27200 19314
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 26884 18838 26936 18844
rect 26988 18822 27108 18850
rect 27160 18896 27212 18902
rect 27160 18838 27212 18844
rect 26988 17954 27016 18822
rect 27068 18692 27120 18698
rect 27068 18634 27120 18640
rect 27080 18086 27108 18634
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 26896 17926 27016 17954
rect 26700 17196 26752 17202
rect 26700 17138 26752 17144
rect 26608 16584 26660 16590
rect 26608 16526 26660 16532
rect 26700 16516 26752 16522
rect 26700 16458 26752 16464
rect 26712 15978 26740 16458
rect 26896 16182 26924 17926
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 26988 17338 27016 17546
rect 26976 17332 27028 17338
rect 26976 17274 27028 17280
rect 27080 17218 27108 18022
rect 26988 17190 27108 17218
rect 27160 17196 27212 17202
rect 26884 16176 26936 16182
rect 26884 16118 26936 16124
rect 26700 15972 26752 15978
rect 26700 15914 26752 15920
rect 26608 15428 26660 15434
rect 26608 15370 26660 15376
rect 26620 15094 26648 15370
rect 26608 15088 26660 15094
rect 26608 15030 26660 15036
rect 26620 14618 26648 15030
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26516 14476 26568 14482
rect 26516 14418 26568 14424
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26252 11354 26280 13330
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26252 10810 26280 11018
rect 26436 10810 26464 13874
rect 26528 13394 26556 14418
rect 26516 13388 26568 13394
rect 26516 13330 26568 13336
rect 26988 12434 27016 17190
rect 27160 17138 27212 17144
rect 27172 16522 27200 17138
rect 27264 16658 27292 19246
rect 27356 18970 27384 19314
rect 27344 18964 27396 18970
rect 27344 18906 27396 18912
rect 27448 17678 27476 20266
rect 27632 19854 27660 22646
rect 28092 22094 28120 31690
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 28736 30734 28764 31078
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 28356 30592 28408 30598
rect 28356 30534 28408 30540
rect 28368 30258 28396 30534
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28724 27872 28776 27878
rect 28724 27814 28776 27820
rect 28736 27402 28764 27814
rect 29012 27606 29040 30670
rect 29000 27600 29052 27606
rect 29052 27548 29132 27554
rect 29000 27542 29132 27548
rect 29012 27526 29132 27542
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 28724 27396 28776 27402
rect 28724 27338 28776 27344
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28172 26784 28224 26790
rect 28172 26726 28224 26732
rect 28184 26314 28212 26726
rect 28644 26586 28672 27270
rect 29012 26586 29040 27406
rect 29104 27062 29132 27526
rect 29092 27056 29144 27062
rect 29092 26998 29144 27004
rect 28632 26580 28684 26586
rect 28632 26522 28684 26528
rect 29000 26580 29052 26586
rect 29000 26522 29052 26528
rect 28724 26444 28776 26450
rect 28724 26386 28776 26392
rect 28172 26308 28224 26314
rect 28172 26250 28224 26256
rect 28632 25968 28684 25974
rect 28632 25910 28684 25916
rect 28540 24676 28592 24682
rect 28540 24618 28592 24624
rect 28552 24206 28580 24618
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28644 24138 28672 25910
rect 28632 24132 28684 24138
rect 28632 24074 28684 24080
rect 28264 23656 28316 23662
rect 28264 23598 28316 23604
rect 28092 22066 28212 22094
rect 27896 21956 27948 21962
rect 27896 21898 27948 21904
rect 27908 21622 27936 21898
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 27712 21548 27764 21554
rect 27712 21490 27764 21496
rect 27724 21146 27752 21490
rect 27712 21140 27764 21146
rect 27764 21100 27844 21128
rect 27712 21082 27764 21088
rect 27712 20800 27764 20806
rect 27712 20742 27764 20748
rect 27724 20058 27752 20742
rect 27816 20602 27844 21100
rect 28184 20806 28212 22066
rect 28276 21554 28304 23598
rect 28448 23044 28500 23050
rect 28448 22986 28500 22992
rect 28460 22710 28488 22986
rect 28448 22704 28500 22710
rect 28448 22646 28500 22652
rect 28356 22432 28408 22438
rect 28356 22374 28408 22380
rect 28368 21604 28396 22374
rect 28460 21894 28488 22646
rect 28644 22642 28672 24074
rect 28632 22636 28684 22642
rect 28632 22578 28684 22584
rect 28448 21888 28500 21894
rect 28448 21830 28500 21836
rect 28448 21616 28500 21622
rect 28368 21576 28448 21604
rect 28448 21558 28500 21564
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28172 20800 28224 20806
rect 28172 20742 28224 20748
rect 27804 20596 27856 20602
rect 27804 20538 27856 20544
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27528 18624 27580 18630
rect 27528 18566 27580 18572
rect 27540 18426 27568 18566
rect 27528 18420 27580 18426
rect 27528 18362 27580 18368
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27356 16658 27384 17274
rect 27436 17196 27488 17202
rect 27436 17138 27488 17144
rect 27448 16794 27476 17138
rect 27436 16788 27488 16794
rect 27436 16730 27488 16736
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27160 16516 27212 16522
rect 27160 16458 27212 16464
rect 27068 14340 27120 14346
rect 27068 14282 27120 14288
rect 27080 13530 27108 14282
rect 27068 13524 27120 13530
rect 27068 13466 27120 13472
rect 27172 12442 27200 16458
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27264 15094 27292 15370
rect 27252 15088 27304 15094
rect 27252 15030 27304 15036
rect 27448 14346 27476 15982
rect 27528 15360 27580 15366
rect 27528 15302 27580 15308
rect 27252 14340 27304 14346
rect 27252 14282 27304 14288
rect 27436 14340 27488 14346
rect 27436 14282 27488 14288
rect 27264 14074 27292 14282
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27436 13796 27488 13802
rect 27436 13738 27488 13744
rect 27448 13326 27476 13738
rect 27540 13326 27568 15302
rect 27724 14618 27752 19994
rect 27908 19174 27936 20402
rect 28276 19990 28304 21490
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28552 20466 28580 20742
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28264 19984 28316 19990
rect 28264 19926 28316 19932
rect 28264 19440 28316 19446
rect 28264 19382 28316 19388
rect 27896 19168 27948 19174
rect 27896 19110 27948 19116
rect 27804 14816 27856 14822
rect 27804 14758 27856 14764
rect 27712 14612 27764 14618
rect 27712 14554 27764 14560
rect 27724 13530 27752 14554
rect 27816 13938 27844 14758
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27252 13320 27304 13326
rect 27252 13262 27304 13268
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 27264 12646 27292 13262
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 27160 12436 27212 12442
rect 26988 12406 27108 12434
rect 26240 10804 26292 10810
rect 26240 10746 26292 10752
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26240 9988 26292 9994
rect 26240 9930 26292 9936
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 26056 9444 26108 9450
rect 26056 9386 26108 9392
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25424 8838 25452 9318
rect 25964 8900 26016 8906
rect 25964 8842 26016 8848
rect 25412 8832 25464 8838
rect 25412 8774 25464 8780
rect 25504 8560 25556 8566
rect 25504 8502 25556 8508
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 25136 8492 25188 8498
rect 25136 8434 25188 8440
rect 24872 8090 24900 8434
rect 24860 8084 24912 8090
rect 24860 8026 24912 8032
rect 24308 7812 24360 7818
rect 24308 7754 24360 7760
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24320 7410 24348 7754
rect 24400 7472 24452 7478
rect 24400 7414 24452 7420
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23860 4826 23888 5578
rect 24320 5574 24348 7346
rect 24412 6390 24440 7414
rect 25148 7410 25176 8434
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 24596 6798 24624 7142
rect 25148 6866 25176 7346
rect 25516 7342 25544 8502
rect 25688 8424 25740 8430
rect 25688 8366 25740 8372
rect 25596 8288 25648 8294
rect 25596 8230 25648 8236
rect 25608 7410 25636 8230
rect 25700 7954 25728 8366
rect 25976 8362 26004 8842
rect 26252 8498 26280 9930
rect 26240 8492 26292 8498
rect 26240 8434 26292 8440
rect 25964 8356 26016 8362
rect 25964 8298 26016 8304
rect 25688 7948 25740 7954
rect 25688 7890 25740 7896
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25504 7336 25556 7342
rect 25504 7278 25556 7284
rect 25136 6860 25188 6866
rect 25136 6802 25188 6808
rect 24584 6792 24636 6798
rect 24584 6734 24636 6740
rect 24768 6792 24820 6798
rect 24768 6734 24820 6740
rect 24780 6458 24808 6734
rect 25516 6730 25544 7278
rect 25504 6724 25556 6730
rect 25504 6666 25556 6672
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24768 6452 24820 6458
rect 24768 6394 24820 6400
rect 24400 6384 24452 6390
rect 24400 6326 24452 6332
rect 24308 5568 24360 5574
rect 24308 5510 24360 5516
rect 24412 4826 24440 6326
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 25056 4554 25084 6598
rect 25700 6458 25728 7890
rect 25780 7744 25832 7750
rect 25780 7686 25832 7692
rect 25792 6866 25820 7686
rect 25976 7410 26004 8298
rect 26252 7886 26280 8434
rect 26436 8430 26464 10746
rect 26976 10464 27028 10470
rect 26976 10406 27028 10412
rect 26988 9994 27016 10406
rect 26976 9988 27028 9994
rect 26976 9930 27028 9936
rect 27080 9874 27108 12406
rect 27160 12378 27212 12384
rect 26988 9846 27108 9874
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26056 7812 26108 7818
rect 26056 7754 26108 7760
rect 26068 7546 26096 7754
rect 26056 7540 26108 7546
rect 26056 7482 26108 7488
rect 25964 7404 26016 7410
rect 25964 7346 26016 7352
rect 25976 7206 26004 7346
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 25780 6860 25832 6866
rect 25780 6802 25832 6808
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25688 6452 25740 6458
rect 25688 6394 25740 6400
rect 25148 4622 25176 6394
rect 26988 6361 27016 9846
rect 27264 6866 27292 12582
rect 27712 11076 27764 11082
rect 27712 11018 27764 11024
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 27356 10606 27384 10950
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27620 10668 27672 10674
rect 27620 10610 27672 10616
rect 27344 10600 27396 10606
rect 27344 10542 27396 10548
rect 27356 10062 27384 10542
rect 27448 10062 27476 10610
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27436 10056 27488 10062
rect 27436 9998 27488 10004
rect 27436 8900 27488 8906
rect 27436 8842 27488 8848
rect 27448 8566 27476 8842
rect 27436 8560 27488 8566
rect 27436 8502 27488 8508
rect 27448 8090 27476 8502
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27632 7698 27660 10610
rect 27724 9178 27752 11018
rect 27804 10668 27856 10674
rect 27804 10610 27856 10616
rect 27712 9172 27764 9178
rect 27712 9114 27764 9120
rect 27816 9110 27844 10610
rect 27804 9104 27856 9110
rect 27804 9046 27856 9052
rect 27632 7670 27844 7698
rect 27712 7540 27764 7546
rect 27712 7482 27764 7488
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 27632 7002 27660 7346
rect 27620 6996 27672 7002
rect 27620 6938 27672 6944
rect 27252 6860 27304 6866
rect 27252 6802 27304 6808
rect 27436 6792 27488 6798
rect 27436 6734 27488 6740
rect 27068 6656 27120 6662
rect 27068 6598 27120 6604
rect 27080 6390 27108 6598
rect 27448 6390 27476 6734
rect 27528 6724 27580 6730
rect 27528 6666 27580 6672
rect 27540 6458 27568 6666
rect 27528 6452 27580 6458
rect 27528 6394 27580 6400
rect 27068 6384 27120 6390
rect 26974 6352 27030 6361
rect 27068 6326 27120 6332
rect 27436 6384 27488 6390
rect 27436 6326 27488 6332
rect 26974 6287 26976 6296
rect 27028 6287 27030 6296
rect 26976 6258 27028 6264
rect 27448 5930 27476 6326
rect 27356 5902 27476 5930
rect 27356 5778 27384 5902
rect 27344 5772 27396 5778
rect 27344 5714 27396 5720
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25424 5370 25452 5646
rect 25412 5364 25464 5370
rect 25412 5306 25464 5312
rect 26424 5296 26476 5302
rect 26422 5264 26424 5273
rect 26476 5264 26478 5273
rect 26422 5199 26478 5208
rect 27356 5098 27384 5714
rect 27724 5710 27752 7482
rect 27816 5846 27844 7670
rect 27804 5840 27856 5846
rect 27804 5782 27856 5788
rect 27712 5704 27764 5710
rect 27712 5646 27764 5652
rect 27436 5568 27488 5574
rect 27436 5510 27488 5516
rect 27448 5234 27476 5510
rect 27908 5302 27936 19110
rect 28080 17060 28132 17066
rect 28080 17002 28132 17008
rect 27988 14884 28040 14890
rect 27988 14826 28040 14832
rect 28000 14482 28028 14826
rect 27988 14476 28040 14482
rect 27988 14418 28040 14424
rect 28092 13938 28120 17002
rect 28276 16182 28304 19382
rect 28264 16176 28316 16182
rect 28264 16118 28316 16124
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28184 15094 28212 16050
rect 28276 15706 28304 16118
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 28172 15088 28224 15094
rect 28172 15030 28224 15036
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 14550 28396 14894
rect 28356 14544 28408 14550
rect 28356 14486 28408 14492
rect 28080 13932 28132 13938
rect 28080 13874 28132 13880
rect 28092 13326 28120 13874
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 28264 12164 28316 12170
rect 28264 12106 28316 12112
rect 28276 11762 28304 12106
rect 28264 11756 28316 11762
rect 28264 11698 28316 11704
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28460 10742 28488 10950
rect 28448 10736 28500 10742
rect 28448 10678 28500 10684
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 28092 9586 28120 10610
rect 28552 10577 28580 20402
rect 28644 19922 28672 22578
rect 28736 21962 28764 26386
rect 28908 25900 28960 25906
rect 28908 25842 28960 25848
rect 28920 24614 28948 25842
rect 29012 25294 29040 26522
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 29000 25152 29052 25158
rect 29000 25094 29052 25100
rect 28908 24608 28960 24614
rect 28908 24550 28960 24556
rect 28920 24410 28948 24550
rect 28908 24404 28960 24410
rect 28908 24346 28960 24352
rect 28816 23724 28868 23730
rect 28816 23666 28868 23672
rect 28828 23526 28856 23666
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28724 21956 28776 21962
rect 28724 21898 28776 21904
rect 28828 20602 28856 23462
rect 28816 20596 28868 20602
rect 28816 20538 28868 20544
rect 29012 20466 29040 25094
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29104 23866 29132 24754
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 29196 23746 29224 31726
rect 29460 31408 29512 31414
rect 29460 31350 29512 31356
rect 29472 30394 29500 31350
rect 29460 30388 29512 30394
rect 29460 30330 29512 30336
rect 29276 30048 29328 30054
rect 29276 29990 29328 29996
rect 29104 23718 29224 23746
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28632 19916 28684 19922
rect 28632 19858 28684 19864
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28632 19780 28684 19786
rect 28632 19722 28684 19728
rect 28644 19514 28672 19722
rect 28920 19689 28948 19790
rect 28906 19680 28962 19689
rect 28906 19615 28962 19624
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 28828 15978 28856 17614
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 28816 15972 28868 15978
rect 28816 15914 28868 15920
rect 28828 15502 28856 15914
rect 28816 15496 28868 15502
rect 28816 15438 28868 15444
rect 28632 15088 28684 15094
rect 28632 15030 28684 15036
rect 28644 14006 28672 15030
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28828 14006 28856 14214
rect 28632 14000 28684 14006
rect 28632 13942 28684 13948
rect 28816 14000 28868 14006
rect 28816 13942 28868 13948
rect 28828 13530 28856 13942
rect 28816 13524 28868 13530
rect 28816 13466 28868 13472
rect 28538 10568 28594 10577
rect 28538 10503 28594 10512
rect 28552 9722 28580 10503
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28080 9580 28132 9586
rect 28080 9522 28132 9528
rect 28092 8974 28120 9522
rect 28724 9444 28776 9450
rect 28724 9386 28776 9392
rect 28736 9042 28764 9386
rect 28724 9036 28776 9042
rect 28724 8978 28776 8984
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28080 8832 28132 8838
rect 28080 8774 28132 8780
rect 28092 8566 28120 8774
rect 28080 8560 28132 8566
rect 28080 8502 28132 8508
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28368 7410 28396 8434
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 28000 6322 28028 7142
rect 27988 6316 28040 6322
rect 27988 6258 28040 6264
rect 28172 6316 28224 6322
rect 28172 6258 28224 6264
rect 28184 5642 28212 6258
rect 28172 5636 28224 5642
rect 28172 5578 28224 5584
rect 27896 5296 27948 5302
rect 27896 5238 27948 5244
rect 28184 5234 28212 5578
rect 28552 5574 28580 8910
rect 28736 8498 28764 8978
rect 28920 8634 28948 16730
rect 29012 16250 29040 17138
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 29012 15638 29040 16186
rect 29000 15632 29052 15638
rect 29000 15574 29052 15580
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 29012 8566 29040 9590
rect 29000 8560 29052 8566
rect 29000 8502 29052 8508
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 29012 8090 29040 8502
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 27344 5092 27396 5098
rect 27344 5034 27396 5040
rect 27252 5024 27304 5030
rect 27252 4966 27304 4972
rect 25136 4616 25188 4622
rect 25136 4558 25188 4564
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 25044 4548 25096 4554
rect 25044 4490 25096 4496
rect 25792 4146 25820 4558
rect 27264 4214 27292 4966
rect 27252 4208 27304 4214
rect 27252 4150 27304 4156
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 28552 4010 28580 5510
rect 29104 5370 29132 23718
rect 29288 23610 29316 29990
rect 29368 28076 29420 28082
rect 29368 28018 29420 28024
rect 29196 23582 29316 23610
rect 29196 16998 29224 23582
rect 29380 23474 29408 28018
rect 29656 27334 29684 33254
rect 29748 32570 29776 36314
rect 30024 33998 30052 39782
rect 30576 39370 30604 39986
rect 30564 39364 30616 39370
rect 30564 39306 30616 39312
rect 30380 39296 30432 39302
rect 30380 39238 30432 39244
rect 30392 38962 30420 39238
rect 30380 38956 30432 38962
rect 30380 38898 30432 38904
rect 30392 38196 30420 38898
rect 30472 38752 30524 38758
rect 30472 38694 30524 38700
rect 30484 38350 30512 38694
rect 30472 38344 30524 38350
rect 30472 38286 30524 38292
rect 30576 38282 30604 39306
rect 30564 38276 30616 38282
rect 30564 38218 30616 38224
rect 30392 38168 30512 38196
rect 30380 37664 30432 37670
rect 30380 37606 30432 37612
rect 30392 36174 30420 37606
rect 30380 36168 30432 36174
rect 30380 36110 30432 36116
rect 30288 35692 30340 35698
rect 30288 35634 30340 35640
rect 30196 34944 30248 34950
rect 30196 34886 30248 34892
rect 30208 34678 30236 34886
rect 30300 34746 30328 35634
rect 30288 34740 30340 34746
rect 30288 34682 30340 34688
rect 30196 34672 30248 34678
rect 30196 34614 30248 34620
rect 30012 33992 30064 33998
rect 30012 33934 30064 33940
rect 30288 33856 30340 33862
rect 30288 33798 30340 33804
rect 29828 33652 29880 33658
rect 29828 33594 29880 33600
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 29748 31822 29776 32506
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 29840 29850 29868 33594
rect 30300 32842 30328 33798
rect 29920 32836 29972 32842
rect 29920 32778 29972 32784
rect 30288 32836 30340 32842
rect 30288 32778 30340 32784
rect 29932 32026 29960 32778
rect 30104 32224 30156 32230
rect 30104 32166 30156 32172
rect 29920 32020 29972 32026
rect 29920 31962 29972 31968
rect 29920 30320 29972 30326
rect 29920 30262 29972 30268
rect 29828 29844 29880 29850
rect 29828 29786 29880 29792
rect 29840 29646 29868 29786
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29644 27328 29696 27334
rect 29644 27270 29696 27276
rect 29736 26308 29788 26314
rect 29736 26250 29788 26256
rect 29552 25696 29604 25702
rect 29552 25638 29604 25644
rect 29564 23730 29592 25638
rect 29644 24744 29696 24750
rect 29644 24686 29696 24692
rect 29656 24410 29684 24686
rect 29644 24404 29696 24410
rect 29644 24346 29696 24352
rect 29552 23724 29604 23730
rect 29552 23666 29604 23672
rect 29460 23588 29512 23594
rect 29460 23530 29512 23536
rect 29288 23446 29408 23474
rect 29288 20942 29316 23446
rect 29368 22976 29420 22982
rect 29472 22964 29500 23530
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 29420 22936 29500 22964
rect 29368 22918 29420 22924
rect 29276 20936 29328 20942
rect 29276 20878 29328 20884
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29184 16448 29236 16454
rect 29184 16390 29236 16396
rect 29196 16096 29224 16390
rect 29276 16108 29328 16114
rect 29196 16068 29276 16096
rect 29196 14550 29224 16068
rect 29276 16050 29328 16056
rect 29184 14544 29236 14550
rect 29184 14486 29236 14492
rect 29196 12714 29224 14486
rect 29184 12708 29236 12714
rect 29184 12650 29236 12656
rect 29380 12374 29408 22918
rect 29564 21418 29592 23258
rect 29748 22642 29776 26250
rect 29828 25152 29880 25158
rect 29828 25094 29880 25100
rect 29840 24682 29868 25094
rect 29828 24676 29880 24682
rect 29828 24618 29880 24624
rect 29840 23662 29868 24618
rect 29932 24410 29960 30262
rect 30116 30258 30144 32166
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 30300 31414 30328 31826
rect 30288 31408 30340 31414
rect 30288 31350 30340 31356
rect 30104 30252 30156 30258
rect 30104 30194 30156 30200
rect 30012 29504 30064 29510
rect 30012 29446 30064 29452
rect 30024 29238 30052 29446
rect 30012 29232 30064 29238
rect 30012 29174 30064 29180
rect 30116 29170 30144 30194
rect 30104 29164 30156 29170
rect 30104 29106 30156 29112
rect 30116 28490 30144 29106
rect 30104 28484 30156 28490
rect 30104 28426 30156 28432
rect 30116 28082 30144 28426
rect 30104 28076 30156 28082
rect 30104 28018 30156 28024
rect 30300 26586 30328 31350
rect 30392 30326 30420 36110
rect 30484 35698 30512 38168
rect 30668 37369 30696 41386
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 30840 40180 30892 40186
rect 30840 40122 30892 40128
rect 30852 39098 30880 40122
rect 31024 40044 31076 40050
rect 31024 39986 31076 39992
rect 31036 39846 31064 39986
rect 31116 39908 31168 39914
rect 31116 39850 31168 39856
rect 31024 39840 31076 39846
rect 31024 39782 31076 39788
rect 31024 39364 31076 39370
rect 31024 39306 31076 39312
rect 30840 39092 30892 39098
rect 30840 39034 30892 39040
rect 30852 38826 30880 39034
rect 31036 38962 31064 39306
rect 31024 38956 31076 38962
rect 31024 38898 31076 38904
rect 30840 38820 30892 38826
rect 30840 38762 30892 38768
rect 30654 37360 30710 37369
rect 30654 37295 30710 37304
rect 30656 35760 30708 35766
rect 30656 35702 30708 35708
rect 30472 35692 30524 35698
rect 30472 35634 30524 35640
rect 30484 35562 30512 35634
rect 30472 35556 30524 35562
rect 30472 35498 30524 35504
rect 30668 33998 30696 35702
rect 30748 35488 30800 35494
rect 30748 35430 30800 35436
rect 30760 35086 30788 35430
rect 30748 35080 30800 35086
rect 30748 35022 30800 35028
rect 30656 33992 30708 33998
rect 30656 33934 30708 33940
rect 30564 33448 30616 33454
rect 30564 33390 30616 33396
rect 30576 32502 30604 33390
rect 30564 32496 30616 32502
rect 30564 32438 30616 32444
rect 30564 32292 30616 32298
rect 30564 32234 30616 32240
rect 30472 32224 30524 32230
rect 30472 32166 30524 32172
rect 30484 30802 30512 32166
rect 30576 30870 30604 32234
rect 30564 30864 30616 30870
rect 30564 30806 30616 30812
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 30380 30320 30432 30326
rect 30380 30262 30432 30268
rect 30576 30190 30604 30806
rect 30668 30802 30696 33934
rect 30748 32496 30800 32502
rect 30748 32438 30800 32444
rect 30760 31906 30788 32438
rect 30852 32230 30880 38762
rect 31128 38010 31156 39850
rect 31300 39840 31352 39846
rect 31300 39782 31352 39788
rect 31312 39438 31340 39782
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 32680 39636 32732 39642
rect 32680 39578 32732 39584
rect 31300 39432 31352 39438
rect 31300 39374 31352 39380
rect 31300 39296 31352 39302
rect 31300 39238 31352 39244
rect 31116 38004 31168 38010
rect 31116 37946 31168 37952
rect 31312 37874 31340 39238
rect 31576 38956 31628 38962
rect 31576 38898 31628 38904
rect 31760 38956 31812 38962
rect 31760 38898 31812 38904
rect 31588 37874 31616 38898
rect 31772 38214 31800 38898
rect 32692 38350 32720 39578
rect 32772 38956 32824 38962
rect 32772 38898 32824 38904
rect 32680 38344 32732 38350
rect 32680 38286 32732 38292
rect 31760 38208 31812 38214
rect 31760 38150 31812 38156
rect 31300 37868 31352 37874
rect 31300 37810 31352 37816
rect 31576 37868 31628 37874
rect 31576 37810 31628 37816
rect 30932 35624 30984 35630
rect 30932 35566 30984 35572
rect 30944 34610 30972 35566
rect 31116 34944 31168 34950
rect 31116 34886 31168 34892
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30944 33998 30972 34546
rect 30932 33992 30984 33998
rect 30932 33934 30984 33940
rect 30944 33318 30972 33934
rect 30932 33312 30984 33318
rect 30932 33254 30984 33260
rect 31024 33108 31076 33114
rect 31024 33050 31076 33056
rect 30840 32224 30892 32230
rect 30840 32166 30892 32172
rect 30760 31878 30880 31906
rect 30748 31816 30800 31822
rect 30748 31758 30800 31764
rect 30656 30796 30708 30802
rect 30656 30738 30708 30744
rect 30564 30184 30616 30190
rect 30564 30126 30616 30132
rect 30576 29238 30604 30126
rect 30656 30048 30708 30054
rect 30656 29990 30708 29996
rect 30564 29232 30616 29238
rect 30564 29174 30616 29180
rect 30576 28626 30604 29174
rect 30668 29102 30696 29990
rect 30760 29306 30788 31758
rect 30852 29782 30880 31878
rect 31036 31822 31064 33050
rect 30932 31816 30984 31822
rect 30932 31758 30984 31764
rect 31024 31816 31076 31822
rect 31024 31758 31076 31764
rect 30944 31346 30972 31758
rect 31128 31414 31156 34886
rect 31312 31822 31340 37810
rect 31484 37460 31536 37466
rect 31484 37402 31536 37408
rect 31496 35494 31524 37402
rect 31588 37330 31616 37810
rect 31576 37324 31628 37330
rect 31576 37266 31628 37272
rect 31484 35488 31536 35494
rect 31484 35430 31536 35436
rect 31496 34542 31524 35430
rect 31484 34536 31536 34542
rect 31484 34478 31536 34484
rect 31576 33924 31628 33930
rect 31576 33866 31628 33872
rect 31588 33114 31616 33866
rect 31576 33108 31628 33114
rect 31576 33050 31628 33056
rect 31668 31952 31720 31958
rect 31668 31894 31720 31900
rect 31300 31816 31352 31822
rect 31300 31758 31352 31764
rect 31208 31748 31260 31754
rect 31208 31690 31260 31696
rect 31220 31414 31248 31690
rect 31116 31408 31168 31414
rect 31116 31350 31168 31356
rect 31208 31408 31260 31414
rect 31208 31350 31260 31356
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 30840 29776 30892 29782
rect 30840 29718 30892 29724
rect 30852 29306 30880 29718
rect 30748 29300 30800 29306
rect 30748 29242 30800 29248
rect 30840 29300 30892 29306
rect 30840 29242 30892 29248
rect 30760 29102 30788 29242
rect 30840 29164 30892 29170
rect 30840 29106 30892 29112
rect 30656 29096 30708 29102
rect 30656 29038 30708 29044
rect 30748 29096 30800 29102
rect 30748 29038 30800 29044
rect 30852 28966 30880 29106
rect 30840 28960 30892 28966
rect 30840 28902 30892 28908
rect 30564 28620 30616 28626
rect 30564 28562 30616 28568
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 30760 28082 30788 28494
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 30472 28008 30524 28014
rect 30472 27950 30524 27956
rect 30484 27606 30512 27950
rect 30472 27600 30524 27606
rect 30472 27542 30524 27548
rect 30288 26580 30340 26586
rect 30288 26522 30340 26528
rect 30012 25900 30064 25906
rect 30012 25842 30064 25848
rect 30024 25430 30052 25842
rect 30472 25696 30524 25702
rect 30472 25638 30524 25644
rect 30012 25424 30064 25430
rect 30012 25366 30064 25372
rect 30484 25294 30512 25638
rect 30472 25288 30524 25294
rect 30472 25230 30524 25236
rect 30564 25288 30616 25294
rect 30564 25230 30616 25236
rect 30576 25140 30604 25230
rect 30484 25112 30604 25140
rect 30484 24886 30512 25112
rect 30472 24880 30524 24886
rect 30472 24822 30524 24828
rect 30380 24608 30432 24614
rect 30380 24550 30432 24556
rect 29920 24404 29972 24410
rect 29920 24346 29972 24352
rect 30392 24206 30420 24550
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 29828 23656 29880 23662
rect 29828 23598 29880 23604
rect 30484 23526 30512 24822
rect 30564 24812 30616 24818
rect 30564 24754 30616 24760
rect 30576 24614 30604 24754
rect 30564 24608 30616 24614
rect 30564 24550 30616 24556
rect 30840 23860 30892 23866
rect 30840 23802 30892 23808
rect 30472 23520 30524 23526
rect 30472 23462 30524 23468
rect 30852 22930 30880 23802
rect 30760 22902 30880 22930
rect 29920 22704 29972 22710
rect 29920 22646 29972 22652
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29552 21412 29604 21418
rect 29552 21354 29604 21360
rect 29828 21344 29880 21350
rect 29828 21286 29880 21292
rect 29840 20602 29868 21286
rect 29552 20596 29604 20602
rect 29552 20538 29604 20544
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29460 20460 29512 20466
rect 29460 20402 29512 20408
rect 29472 19446 29500 20402
rect 29564 19700 29592 20538
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29656 19854 29684 20402
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29564 19672 29684 19700
rect 29460 19440 29512 19446
rect 29460 19382 29512 19388
rect 29656 18358 29684 19672
rect 29932 19310 29960 22646
rect 30104 21480 30156 21486
rect 30104 21422 30156 21428
rect 30012 19848 30064 19854
rect 30012 19790 30064 19796
rect 29920 19304 29972 19310
rect 29840 19264 29920 19292
rect 29840 19174 29868 19264
rect 29920 19246 29972 19252
rect 30024 19242 30052 19790
rect 30012 19236 30064 19242
rect 30012 19178 30064 19184
rect 29828 19168 29880 19174
rect 29828 19110 29880 19116
rect 29840 18766 29868 19110
rect 30024 18766 30052 19178
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 30012 18760 30064 18766
rect 30012 18702 30064 18708
rect 29920 18692 29972 18698
rect 29920 18634 29972 18640
rect 29644 18352 29696 18358
rect 29644 18294 29696 18300
rect 29460 16040 29512 16046
rect 29460 15982 29512 15988
rect 29472 14890 29500 15982
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29564 15502 29592 15846
rect 29552 15496 29604 15502
rect 29552 15438 29604 15444
rect 29552 15020 29604 15026
rect 29552 14962 29604 14968
rect 29460 14884 29512 14890
rect 29460 14826 29512 14832
rect 29472 13938 29500 14826
rect 29564 14822 29592 14962
rect 29552 14816 29604 14822
rect 29552 14758 29604 14764
rect 29460 13932 29512 13938
rect 29460 13874 29512 13880
rect 29368 12368 29420 12374
rect 29368 12310 29420 12316
rect 29184 9716 29236 9722
rect 29184 9658 29236 9664
rect 29196 6458 29224 9658
rect 29564 8362 29592 14758
rect 29656 11898 29684 18294
rect 29932 17270 29960 18634
rect 30012 18624 30064 18630
rect 30012 18566 30064 18572
rect 29920 17264 29972 17270
rect 29920 17206 29972 17212
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 29840 16130 29868 16526
rect 29932 16250 29960 17206
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 29840 16114 29960 16130
rect 29840 16108 29972 16114
rect 29840 16102 29920 16108
rect 29920 16050 29972 16056
rect 29932 14958 29960 16050
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 29840 14074 29868 14350
rect 29828 14068 29880 14074
rect 29828 14010 29880 14016
rect 29932 13870 29960 14894
rect 29920 13864 29972 13870
rect 29920 13806 29972 13812
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 29920 11280 29972 11286
rect 29920 11222 29972 11228
rect 29552 8356 29604 8362
rect 29552 8298 29604 8304
rect 29828 7200 29880 7206
rect 29828 7142 29880 7148
rect 29184 6452 29236 6458
rect 29184 6394 29236 6400
rect 29840 6322 29868 7142
rect 29828 6316 29880 6322
rect 29828 6258 29880 6264
rect 29932 5914 29960 11222
rect 30024 11082 30052 18566
rect 30012 11076 30064 11082
rect 30012 11018 30064 11024
rect 30116 9178 30144 21422
rect 30196 21004 30248 21010
rect 30196 20946 30248 20952
rect 30208 11286 30236 20946
rect 30760 20534 30788 22902
rect 30932 22432 30984 22438
rect 30932 22374 30984 22380
rect 30838 21992 30894 22001
rect 30838 21927 30840 21936
rect 30892 21927 30894 21936
rect 30840 21898 30892 21904
rect 30840 20868 30892 20874
rect 30944 20856 30972 22374
rect 31036 22094 31064 31078
rect 31220 30326 31248 31350
rect 31392 30728 31444 30734
rect 31392 30670 31444 30676
rect 31208 30320 31260 30326
rect 31208 30262 31260 30268
rect 31404 30054 31432 30670
rect 31392 30048 31444 30054
rect 31392 29990 31444 29996
rect 31484 29844 31536 29850
rect 31484 29786 31536 29792
rect 31496 29753 31524 29786
rect 31482 29744 31538 29753
rect 31482 29679 31538 29688
rect 31208 29640 31260 29646
rect 31208 29582 31260 29588
rect 31220 29510 31248 29582
rect 31208 29504 31260 29510
rect 31208 29446 31260 29452
rect 31220 27062 31248 29446
rect 31392 28960 31444 28966
rect 31392 28902 31444 28908
rect 31404 28558 31432 28902
rect 31392 28552 31444 28558
rect 31392 28494 31444 28500
rect 31404 27130 31432 28494
rect 31392 27124 31444 27130
rect 31392 27066 31444 27072
rect 31208 27056 31260 27062
rect 31208 26998 31260 27004
rect 31300 25696 31352 25702
rect 31300 25638 31352 25644
rect 31312 25498 31340 25638
rect 31300 25492 31352 25498
rect 31300 25434 31352 25440
rect 31312 25294 31340 25434
rect 31300 25288 31352 25294
rect 31300 25230 31352 25236
rect 31116 24404 31168 24410
rect 31116 24346 31168 24352
rect 31128 22234 31156 24346
rect 31208 22704 31260 22710
rect 31208 22646 31260 22652
rect 31116 22228 31168 22234
rect 31116 22170 31168 22176
rect 31036 22066 31156 22094
rect 30892 20828 30972 20856
rect 30840 20810 30892 20816
rect 30748 20528 30800 20534
rect 30748 20470 30800 20476
rect 30564 20392 30616 20398
rect 30564 20334 30616 20340
rect 30472 20256 30524 20262
rect 30472 20198 30524 20204
rect 30484 20058 30512 20198
rect 30472 20052 30524 20058
rect 30472 19994 30524 20000
rect 30380 18896 30432 18902
rect 30380 18838 30432 18844
rect 30392 16454 30420 18838
rect 30472 16992 30524 16998
rect 30472 16934 30524 16940
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30392 15162 30420 16050
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30484 15026 30512 16934
rect 30576 16794 30604 20334
rect 30656 18896 30708 18902
rect 30654 18864 30656 18873
rect 30708 18864 30710 18873
rect 30654 18799 30710 18808
rect 30564 16788 30616 16794
rect 30564 16730 30616 16736
rect 30564 16516 30616 16522
rect 30564 16458 30616 16464
rect 30576 16182 30604 16458
rect 30564 16176 30616 16182
rect 30564 16118 30616 16124
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30380 14612 30432 14618
rect 30380 14554 30432 14560
rect 30392 14346 30420 14554
rect 30380 14340 30432 14346
rect 30380 14282 30432 14288
rect 30392 12434 30420 14282
rect 30656 14000 30708 14006
rect 30656 13942 30708 13948
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30576 13258 30604 13806
rect 30564 13252 30616 13258
rect 30564 13194 30616 13200
rect 30668 12434 30696 13942
rect 30392 12406 30512 12434
rect 30668 12406 30788 12434
rect 30288 11552 30340 11558
rect 30288 11494 30340 11500
rect 30196 11280 30248 11286
rect 30196 11222 30248 11228
rect 30300 11150 30328 11494
rect 30196 11144 30248 11150
rect 30196 11086 30248 11092
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30104 9172 30156 9178
rect 30104 9114 30156 9120
rect 30208 8634 30236 11086
rect 30484 10606 30512 12406
rect 30564 11756 30616 11762
rect 30564 11698 30616 11704
rect 30576 10810 30604 11698
rect 30564 10804 30616 10810
rect 30564 10746 30616 10752
rect 30472 10600 30524 10606
rect 30472 10542 30524 10548
rect 30380 9920 30432 9926
rect 30380 9862 30432 9868
rect 30392 9586 30420 9862
rect 30380 9580 30432 9586
rect 30380 9522 30432 9528
rect 30392 9382 30420 9522
rect 30380 9376 30432 9382
rect 30380 9318 30432 9324
rect 30484 8634 30512 10542
rect 30012 8628 30064 8634
rect 30012 8570 30064 8576
rect 30196 8628 30248 8634
rect 30196 8570 30248 8576
rect 30472 8628 30524 8634
rect 30472 8570 30524 8576
rect 30024 6866 30052 8570
rect 30012 6860 30064 6866
rect 30012 6802 30064 6808
rect 30380 6724 30432 6730
rect 30380 6666 30432 6672
rect 30392 6458 30420 6666
rect 30656 6656 30708 6662
rect 30656 6598 30708 6604
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 30116 6322 30144 6394
rect 30104 6316 30156 6322
rect 30104 6258 30156 6264
rect 30104 6180 30156 6186
rect 30104 6122 30156 6128
rect 30012 6112 30064 6118
rect 30012 6054 30064 6060
rect 29920 5908 29972 5914
rect 29920 5850 29972 5856
rect 29932 5574 29960 5850
rect 30024 5778 30052 6054
rect 30012 5772 30064 5778
rect 30012 5714 30064 5720
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29920 5568 29972 5574
rect 29920 5510 29972 5516
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 28540 4004 28592 4010
rect 28540 3946 28592 3952
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 23584 2378 23612 2518
rect 23572 2372 23624 2378
rect 23572 2314 23624 2320
rect 23676 800 23704 3470
rect 23952 800 23980 3470
rect 24228 800 24256 3878
rect 25516 3670 25544 3878
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24504 800 24532 2926
rect 24780 800 24808 3470
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25320 2848 25372 2854
rect 25320 2790 25372 2796
rect 25056 800 25084 2790
rect 25332 800 25360 2790
rect 25608 800 25636 3470
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 25884 800 25912 2382
rect 26160 800 26188 2790
rect 26424 2576 26476 2582
rect 26424 2518 26476 2524
rect 26436 800 26464 2518
rect 26712 800 26740 3470
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 26896 898 26924 2790
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 27356 2446 27384 2586
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 26896 870 27016 898
rect 26988 800 27016 870
rect 27264 800 27292 2382
rect 27540 800 27568 3470
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 27816 800 27844 2790
rect 28092 800 28120 2790
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28368 800 28396 2518
rect 28644 800 28672 3470
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 28920 800 28948 2382
rect 29196 800 29224 2790
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 29472 800 29500 2382
rect 29564 1902 29592 5510
rect 29736 5364 29788 5370
rect 29736 5306 29788 5312
rect 29748 4282 29776 5306
rect 30024 5166 30052 5714
rect 30116 5710 30144 6122
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 30196 5840 30248 5846
rect 30196 5782 30248 5788
rect 30208 5710 30236 5782
rect 30104 5704 30156 5710
rect 30104 5646 30156 5652
rect 30196 5704 30248 5710
rect 30196 5646 30248 5652
rect 30116 5234 30144 5646
rect 30392 5234 30420 6054
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30576 5642 30604 5850
rect 30668 5710 30696 6598
rect 30656 5704 30708 5710
rect 30656 5646 30708 5652
rect 30564 5636 30616 5642
rect 30564 5578 30616 5584
rect 30760 5370 30788 12406
rect 30852 12374 30880 20810
rect 30930 19816 30986 19825
rect 30930 19751 30986 19760
rect 30944 19514 30972 19751
rect 30932 19508 30984 19514
rect 30932 19450 30984 19456
rect 31128 18766 31156 22066
rect 31220 21962 31248 22646
rect 31208 21956 31260 21962
rect 31208 21898 31260 21904
rect 31208 19372 31260 19378
rect 31208 19314 31260 19320
rect 31116 18760 31168 18766
rect 31116 18702 31168 18708
rect 31024 13252 31076 13258
rect 31024 13194 31076 13200
rect 30840 12368 30892 12374
rect 30840 12310 30892 12316
rect 31036 12186 31064 13194
rect 30852 12170 31064 12186
rect 30852 12164 31076 12170
rect 30852 12158 31024 12164
rect 30852 11830 30880 12158
rect 31024 12106 31076 12112
rect 31036 12075 31064 12106
rect 30840 11824 30892 11830
rect 30840 11766 30892 11772
rect 30852 9926 30880 11766
rect 31024 11008 31076 11014
rect 31024 10950 31076 10956
rect 31036 10742 31064 10950
rect 31024 10736 31076 10742
rect 31024 10678 31076 10684
rect 30932 10056 30984 10062
rect 30932 9998 30984 10004
rect 30840 9920 30892 9926
rect 30840 9862 30892 9868
rect 30944 9654 30972 9998
rect 31036 9722 31064 10678
rect 31220 10538 31248 19314
rect 31312 17066 31340 25230
rect 31484 24608 31536 24614
rect 31484 24550 31536 24556
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31404 22166 31432 22578
rect 31496 22438 31524 24550
rect 31576 23792 31628 23798
rect 31576 23734 31628 23740
rect 31484 22432 31536 22438
rect 31484 22374 31536 22380
rect 31484 22228 31536 22234
rect 31484 22170 31536 22176
rect 31392 22160 31444 22166
rect 31392 22102 31444 22108
rect 31404 19854 31432 22102
rect 31392 19848 31444 19854
rect 31392 19790 31444 19796
rect 31300 17060 31352 17066
rect 31300 17002 31352 17008
rect 31312 13938 31340 17002
rect 31496 14074 31524 22170
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31300 13932 31352 13938
rect 31300 13874 31352 13880
rect 31312 13530 31340 13874
rect 31300 13524 31352 13530
rect 31300 13466 31352 13472
rect 31484 12368 31536 12374
rect 31484 12310 31536 12316
rect 31496 12238 31524 12310
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 31484 12232 31536 12238
rect 31484 12174 31536 12180
rect 31312 11898 31340 12174
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 31300 10736 31352 10742
rect 31300 10678 31352 10684
rect 31208 10532 31260 10538
rect 31208 10474 31260 10480
rect 31208 10056 31260 10062
rect 31128 10016 31208 10044
rect 31024 9716 31076 9722
rect 31024 9658 31076 9664
rect 30932 9648 30984 9654
rect 30932 9590 30984 9596
rect 31024 9580 31076 9586
rect 31024 9522 31076 9528
rect 31036 7478 31064 9522
rect 31128 9518 31156 10016
rect 31208 9998 31260 10004
rect 31208 9580 31260 9586
rect 31208 9522 31260 9528
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 31220 9042 31248 9522
rect 31312 9382 31340 10678
rect 31484 9920 31536 9926
rect 31484 9862 31536 9868
rect 31300 9376 31352 9382
rect 31300 9318 31352 9324
rect 31208 9036 31260 9042
rect 31208 8978 31260 8984
rect 31312 8974 31340 9318
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 31116 8492 31168 8498
rect 31116 8434 31168 8440
rect 31024 7472 31076 7478
rect 31024 7414 31076 7420
rect 30932 7200 30984 7206
rect 30932 7142 30984 7148
rect 30944 7002 30972 7142
rect 31036 7002 31064 7414
rect 30932 6996 30984 7002
rect 30932 6938 30984 6944
rect 31024 6996 31076 7002
rect 31024 6938 31076 6944
rect 31128 6662 31156 8434
rect 31496 7886 31524 9862
rect 31588 9450 31616 23734
rect 31680 19446 31708 31894
rect 31772 31346 31800 38150
rect 32784 38010 32812 38898
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 33048 38276 33100 38282
rect 33048 38218 33100 38224
rect 33140 38276 33192 38282
rect 33140 38218 33192 38224
rect 33060 38010 33088 38218
rect 32772 38004 32824 38010
rect 32772 37946 32824 37952
rect 33048 38004 33100 38010
rect 33048 37946 33100 37952
rect 32588 37868 32640 37874
rect 32588 37810 32640 37816
rect 32600 37466 32628 37810
rect 32588 37460 32640 37466
rect 32588 37402 32640 37408
rect 32784 35086 32812 37946
rect 33048 37868 33100 37874
rect 33048 37810 33100 37816
rect 33060 37670 33088 37810
rect 33048 37664 33100 37670
rect 33048 37606 33100 37612
rect 32128 35080 32180 35086
rect 32128 35022 32180 35028
rect 32772 35080 32824 35086
rect 32772 35022 32824 35028
rect 32140 34610 32168 35022
rect 32128 34604 32180 34610
rect 32128 34546 32180 34552
rect 32140 32842 32168 34546
rect 32128 32836 32180 32842
rect 32128 32778 32180 32784
rect 31760 31340 31812 31346
rect 31760 31282 31812 31288
rect 31852 30660 31904 30666
rect 31852 30602 31904 30608
rect 31864 28422 31892 30602
rect 32140 30598 32168 32778
rect 32404 32768 32456 32774
rect 32404 32710 32456 32716
rect 32416 31822 32444 32710
rect 32404 31816 32456 31822
rect 32404 31758 32456 31764
rect 32784 31482 32812 35022
rect 33060 34678 33088 37606
rect 33152 36582 33180 38218
rect 33508 38208 33560 38214
rect 33508 38150 33560 38156
rect 33324 37324 33376 37330
rect 33324 37266 33376 37272
rect 33140 36576 33192 36582
rect 33140 36518 33192 36524
rect 33152 35154 33180 36518
rect 33336 36242 33364 37266
rect 33416 37256 33468 37262
rect 33416 37198 33468 37204
rect 33324 36236 33376 36242
rect 33324 36178 33376 36184
rect 33336 35630 33364 36178
rect 33428 36106 33456 37198
rect 33520 37126 33548 38150
rect 33784 37800 33836 37806
rect 33784 37742 33836 37748
rect 33796 37262 33824 37742
rect 34336 37664 34388 37670
rect 34336 37606 34388 37612
rect 34244 37324 34296 37330
rect 34244 37266 34296 37272
rect 33692 37256 33744 37262
rect 33692 37198 33744 37204
rect 33784 37256 33836 37262
rect 33784 37198 33836 37204
rect 33508 37120 33560 37126
rect 33508 37062 33560 37068
rect 33416 36100 33468 36106
rect 33416 36042 33468 36048
rect 33428 35698 33456 36042
rect 33416 35692 33468 35698
rect 33416 35634 33468 35640
rect 33324 35624 33376 35630
rect 33324 35566 33376 35572
rect 33140 35148 33192 35154
rect 33140 35090 33192 35096
rect 33048 34672 33100 34678
rect 33048 34614 33100 34620
rect 32956 33380 33008 33386
rect 32956 33322 33008 33328
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32876 32026 32904 32370
rect 32864 32020 32916 32026
rect 32864 31962 32916 31968
rect 32968 31890 32996 33322
rect 33060 32502 33088 34614
rect 33152 32910 33180 35090
rect 33336 34542 33364 35566
rect 33428 34610 33456 35634
rect 33416 34604 33468 34610
rect 33416 34546 33468 34552
rect 33324 34536 33376 34542
rect 33324 34478 33376 34484
rect 33336 33998 33364 34478
rect 33324 33992 33376 33998
rect 33324 33934 33376 33940
rect 33232 33924 33284 33930
rect 33232 33866 33284 33872
rect 33244 33454 33272 33866
rect 33232 33448 33284 33454
rect 33232 33390 33284 33396
rect 33140 32904 33192 32910
rect 33140 32846 33192 32852
rect 33232 32836 33284 32842
rect 33232 32778 33284 32784
rect 33048 32496 33100 32502
rect 33048 32438 33100 32444
rect 33244 32230 33272 32778
rect 33232 32224 33284 32230
rect 33232 32166 33284 32172
rect 33336 31958 33364 33934
rect 33428 33522 33456 34546
rect 33416 33516 33468 33522
rect 33416 33458 33468 33464
rect 33324 31952 33376 31958
rect 33324 31894 33376 31900
rect 32956 31884 33008 31890
rect 32956 31826 33008 31832
rect 32864 31816 32916 31822
rect 32864 31758 32916 31764
rect 32772 31476 32824 31482
rect 32772 31418 32824 31424
rect 32876 31142 32904 31758
rect 33140 31272 33192 31278
rect 33140 31214 33192 31220
rect 33232 31272 33284 31278
rect 33232 31214 33284 31220
rect 32864 31136 32916 31142
rect 32864 31078 32916 31084
rect 32588 30660 32640 30666
rect 32588 30602 32640 30608
rect 32128 30592 32180 30598
rect 32128 30534 32180 30540
rect 32312 30592 32364 30598
rect 32312 30534 32364 30540
rect 31944 29640 31996 29646
rect 31944 29582 31996 29588
rect 31852 28416 31904 28422
rect 31852 28358 31904 28364
rect 31864 26858 31892 28358
rect 31956 26926 31984 29582
rect 32324 29578 32352 30534
rect 32600 30326 32628 30602
rect 32588 30320 32640 30326
rect 32588 30262 32640 30268
rect 32876 30122 32904 31078
rect 33152 30734 33180 31214
rect 33244 30734 33272 31214
rect 33520 30734 33548 37062
rect 33704 36378 33732 37198
rect 33692 36372 33744 36378
rect 33692 36314 33744 36320
rect 34256 36038 34284 37266
rect 34348 37262 34376 37606
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34336 37256 34388 37262
rect 34336 37198 34388 37204
rect 34244 36032 34296 36038
rect 34244 35974 34296 35980
rect 34060 34944 34112 34950
rect 34060 34886 34112 34892
rect 34072 34406 34100 34886
rect 34256 34474 34284 35974
rect 34244 34468 34296 34474
rect 34244 34410 34296 34416
rect 34060 34400 34112 34406
rect 34060 34342 34112 34348
rect 33692 33992 33744 33998
rect 33692 33934 33744 33940
rect 33704 33658 33732 33934
rect 33968 33856 34020 33862
rect 33968 33798 34020 33804
rect 33692 33652 33744 33658
rect 33692 33594 33744 33600
rect 33980 33522 34008 33798
rect 33968 33516 34020 33522
rect 33968 33458 34020 33464
rect 33784 32224 33836 32230
rect 33784 32166 33836 32172
rect 33140 30728 33192 30734
rect 33140 30670 33192 30676
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 32956 30592 33008 30598
rect 32956 30534 33008 30540
rect 32864 30116 32916 30122
rect 32864 30058 32916 30064
rect 32312 29572 32364 29578
rect 32312 29514 32364 29520
rect 32772 27464 32824 27470
rect 32772 27406 32824 27412
rect 32312 27328 32364 27334
rect 32312 27270 32364 27276
rect 31944 26920 31996 26926
rect 31944 26862 31996 26868
rect 31852 26852 31904 26858
rect 31852 26794 31904 26800
rect 31956 26450 31984 26862
rect 31944 26444 31996 26450
rect 31944 26386 31996 26392
rect 31956 25294 31984 26386
rect 31944 25288 31996 25294
rect 31944 25230 31996 25236
rect 31956 24274 31984 25230
rect 31944 24268 31996 24274
rect 31944 24210 31996 24216
rect 32324 24070 32352 27270
rect 32404 27124 32456 27130
rect 32404 27066 32456 27072
rect 32416 26994 32444 27066
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 32588 26988 32640 26994
rect 32588 26930 32640 26936
rect 32600 24818 32628 26930
rect 32784 26042 32812 27406
rect 32876 26858 32904 30058
rect 32864 26852 32916 26858
rect 32864 26794 32916 26800
rect 32772 26036 32824 26042
rect 32772 25978 32824 25984
rect 32784 24886 32812 25978
rect 32772 24880 32824 24886
rect 32772 24822 32824 24828
rect 32588 24812 32640 24818
rect 32588 24754 32640 24760
rect 32312 24064 32364 24070
rect 32312 24006 32364 24012
rect 32968 23798 32996 30534
rect 33152 30258 33180 30670
rect 33416 30660 33468 30666
rect 33416 30602 33468 30608
rect 33140 30252 33192 30258
rect 33140 30194 33192 30200
rect 33324 30048 33376 30054
rect 33324 29990 33376 29996
rect 33232 29504 33284 29510
rect 33232 29446 33284 29452
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33152 27402 33180 27950
rect 33244 27470 33272 29446
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33140 27396 33192 27402
rect 33140 27338 33192 27344
rect 33336 23798 33364 29990
rect 33428 29170 33456 30602
rect 33692 30320 33744 30326
rect 33692 30262 33744 30268
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33416 29164 33468 29170
rect 33416 29106 33468 29112
rect 33520 28626 33548 30194
rect 33704 30122 33732 30262
rect 33692 30116 33744 30122
rect 33692 30058 33744 30064
rect 33600 29096 33652 29102
rect 33600 29038 33652 29044
rect 33508 28620 33560 28626
rect 33508 28562 33560 28568
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33428 28082 33456 28494
rect 33612 28490 33640 29038
rect 33600 28484 33652 28490
rect 33600 28426 33652 28432
rect 33416 28076 33468 28082
rect 33416 28018 33468 28024
rect 33428 27470 33456 28018
rect 33612 28014 33640 28426
rect 33600 28008 33652 28014
rect 33600 27950 33652 27956
rect 33796 27470 33824 32166
rect 33980 30818 34008 33458
rect 34072 31686 34100 34342
rect 34256 33998 34284 34410
rect 34244 33992 34296 33998
rect 34244 33934 34296 33940
rect 34060 31680 34112 31686
rect 34060 31622 34112 31628
rect 34072 30938 34100 31622
rect 34060 30932 34112 30938
rect 34060 30874 34112 30880
rect 33980 30790 34100 30818
rect 33876 30660 33928 30666
rect 33876 30602 33928 30608
rect 33888 30258 33916 30602
rect 34072 30258 34100 30790
rect 33876 30252 33928 30258
rect 33876 30194 33928 30200
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 33876 30048 33928 30054
rect 33876 29990 33928 29996
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 33784 27464 33836 27470
rect 33784 27406 33836 27412
rect 33508 27328 33560 27334
rect 33508 27270 33560 27276
rect 33520 24698 33548 27270
rect 33600 26784 33652 26790
rect 33600 26726 33652 26732
rect 33612 25974 33640 26726
rect 33600 25968 33652 25974
rect 33600 25910 33652 25916
rect 33520 24670 33640 24698
rect 32956 23792 33008 23798
rect 32956 23734 33008 23740
rect 33324 23792 33376 23798
rect 33324 23734 33376 23740
rect 32496 23520 32548 23526
rect 32496 23462 32548 23468
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32772 23520 32824 23526
rect 32772 23462 32824 23468
rect 33508 23520 33560 23526
rect 33508 23462 33560 23468
rect 32312 22976 32364 22982
rect 32312 22918 32364 22924
rect 32324 22710 32352 22918
rect 32312 22704 32364 22710
rect 32312 22646 32364 22652
rect 32508 22574 32536 23462
rect 32588 22636 32640 22642
rect 32588 22578 32640 22584
rect 32496 22568 32548 22574
rect 31758 22536 31814 22545
rect 32496 22510 32548 22516
rect 31758 22471 31760 22480
rect 31812 22471 31814 22480
rect 31760 22442 31812 22448
rect 31852 22024 31904 22030
rect 31852 21966 31904 21972
rect 31668 19440 31720 19446
rect 31668 19382 31720 19388
rect 31864 19334 31892 21966
rect 32600 20466 32628 22578
rect 32692 21894 32720 23462
rect 32784 22778 32812 23462
rect 33416 23044 33468 23050
rect 33416 22986 33468 22992
rect 32864 22976 32916 22982
rect 32864 22918 32916 22924
rect 32772 22772 32824 22778
rect 32772 22714 32824 22720
rect 32772 22024 32824 22030
rect 32770 21992 32772 22001
rect 32824 21992 32826 22001
rect 32770 21927 32826 21936
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 32876 21622 32904 22918
rect 33428 22778 33456 22986
rect 33416 22772 33468 22778
rect 33416 22714 33468 22720
rect 32956 22500 33008 22506
rect 32956 22442 33008 22448
rect 33048 22500 33100 22506
rect 33048 22442 33100 22448
rect 32864 21616 32916 21622
rect 32864 21558 32916 21564
rect 32968 21486 32996 22442
rect 32956 21480 33008 21486
rect 32956 21422 33008 21428
rect 32956 21344 33008 21350
rect 32956 21286 33008 21292
rect 32968 21146 32996 21286
rect 32956 21140 33008 21146
rect 32956 21082 33008 21088
rect 32968 20466 32996 21082
rect 33060 20516 33088 22442
rect 33140 22160 33192 22166
rect 33140 22102 33192 22108
rect 33152 22030 33180 22102
rect 33140 22024 33192 22030
rect 33140 21966 33192 21972
rect 33520 21690 33548 23462
rect 33508 21684 33560 21690
rect 33508 21626 33560 21632
rect 33324 21548 33376 21554
rect 33324 21490 33376 21496
rect 33140 20528 33192 20534
rect 33060 20488 33140 20516
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32772 20460 32824 20466
rect 32956 20460 33008 20466
rect 32824 20420 32904 20448
rect 32772 20402 32824 20408
rect 32600 19334 32628 20402
rect 32772 20324 32824 20330
rect 32772 20266 32824 20272
rect 32784 19854 32812 20266
rect 32876 20058 32904 20420
rect 32956 20402 33008 20408
rect 32864 20052 32916 20058
rect 32864 19994 32916 20000
rect 32772 19848 32824 19854
rect 32772 19790 32824 19796
rect 32680 19780 32732 19786
rect 32680 19722 32732 19728
rect 31864 19306 32076 19334
rect 32048 18902 32076 19306
rect 32416 19306 32628 19334
rect 32036 18896 32088 18902
rect 32036 18838 32088 18844
rect 31852 18420 31904 18426
rect 31852 18362 31904 18368
rect 32128 18420 32180 18426
rect 32128 18362 32180 18368
rect 31760 16040 31812 16046
rect 31760 15982 31812 15988
rect 31772 15502 31800 15982
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31772 14278 31800 15438
rect 31760 14272 31812 14278
rect 31760 14214 31812 14220
rect 31772 13394 31800 14214
rect 31760 13388 31812 13394
rect 31760 13330 31812 13336
rect 31668 12844 31720 12850
rect 31668 12786 31720 12792
rect 31680 11830 31708 12786
rect 31760 12300 31812 12306
rect 31760 12242 31812 12248
rect 31668 11824 31720 11830
rect 31668 11766 31720 11772
rect 31680 10742 31708 11766
rect 31772 11762 31800 12242
rect 31760 11756 31812 11762
rect 31760 11698 31812 11704
rect 31668 10736 31720 10742
rect 31668 10678 31720 10684
rect 31772 10130 31800 11698
rect 31760 10124 31812 10130
rect 31760 10066 31812 10072
rect 31668 9988 31720 9994
rect 31668 9930 31720 9936
rect 31680 9654 31708 9930
rect 31668 9648 31720 9654
rect 31668 9590 31720 9596
rect 31772 9586 31800 10066
rect 31864 10062 31892 18362
rect 32140 18154 32168 18362
rect 32416 18290 32444 19306
rect 32692 19242 32720 19722
rect 32968 19718 32996 20402
rect 32956 19712 33008 19718
rect 32956 19654 33008 19660
rect 32680 19236 32732 19242
rect 32680 19178 32732 19184
rect 32692 18766 32720 19178
rect 32864 18896 32916 18902
rect 32864 18838 32916 18844
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32600 18290 32628 18566
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32588 18284 32640 18290
rect 32588 18226 32640 18232
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32128 18148 32180 18154
rect 32128 18090 32180 18096
rect 32416 17338 32444 18226
rect 32784 18154 32812 18226
rect 32772 18148 32824 18154
rect 32772 18090 32824 18096
rect 32876 17678 32904 18838
rect 32864 17672 32916 17678
rect 32864 17614 32916 17620
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32128 17128 32180 17134
rect 32128 17070 32180 17076
rect 32140 16658 32168 17070
rect 32128 16652 32180 16658
rect 32128 16594 32180 16600
rect 32496 13320 32548 13326
rect 32496 13262 32548 13268
rect 32680 13320 32732 13326
rect 32680 13262 32732 13268
rect 32508 12306 32536 13262
rect 32692 12986 32720 13262
rect 32680 12980 32732 12986
rect 32680 12922 32732 12928
rect 32496 12300 32548 12306
rect 32496 12242 32548 12248
rect 32404 12096 32456 12102
rect 32404 12038 32456 12044
rect 32416 11762 32444 12038
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 31852 10056 31904 10062
rect 31852 9998 31904 10004
rect 32036 10056 32088 10062
rect 32036 9998 32088 10004
rect 31760 9580 31812 9586
rect 31760 9522 31812 9528
rect 31576 9444 31628 9450
rect 31576 9386 31628 9392
rect 31576 8900 31628 8906
rect 31576 8842 31628 8848
rect 31484 7880 31536 7886
rect 31484 7822 31536 7828
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 31116 6656 31168 6662
rect 31116 6598 31168 6604
rect 31220 6322 31248 7346
rect 31588 7274 31616 8842
rect 31576 7268 31628 7274
rect 31576 7210 31628 7216
rect 32048 6322 32076 9998
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 32232 9042 32260 9862
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 32324 9178 32352 9522
rect 32312 9172 32364 9178
rect 32312 9114 32364 9120
rect 32220 9036 32272 9042
rect 32220 8978 32272 8984
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 31208 6316 31260 6322
rect 31208 6258 31260 6264
rect 32036 6316 32088 6322
rect 32036 6258 32088 6264
rect 31220 5642 31248 6258
rect 31668 5704 31720 5710
rect 31668 5646 31720 5652
rect 31208 5636 31260 5642
rect 31208 5578 31260 5584
rect 31116 5568 31168 5574
rect 31116 5510 31168 5516
rect 30748 5364 30800 5370
rect 30748 5306 30800 5312
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 30380 5228 30432 5234
rect 30380 5170 30432 5176
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 29736 4276 29788 4282
rect 29736 4218 29788 4224
rect 30852 3534 30880 4966
rect 31128 4622 31156 5510
rect 31680 5370 31708 5646
rect 31668 5364 31720 5370
rect 31668 5306 31720 5312
rect 30932 4616 30984 4622
rect 30932 4558 30984 4564
rect 31116 4616 31168 4622
rect 31116 4558 31168 4564
rect 30944 4146 30972 4558
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30944 3602 30972 4082
rect 32048 3738 32076 6258
rect 32140 5642 32168 8910
rect 32232 8906 32260 8978
rect 32416 8974 32444 11698
rect 32508 11218 32536 12242
rect 32496 11212 32548 11218
rect 32496 11154 32548 11160
rect 32588 10056 32640 10062
rect 32588 9998 32640 10004
rect 32600 9518 32628 9998
rect 32968 9654 32996 19654
rect 33060 18222 33088 20488
rect 33140 20470 33192 20476
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 33152 19854 33180 20198
rect 33336 19854 33364 21490
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 33324 19848 33376 19854
rect 33324 19790 33376 19796
rect 33232 19372 33284 19378
rect 33232 19314 33284 19320
rect 33244 18426 33272 19314
rect 33336 18698 33364 19790
rect 33324 18692 33376 18698
rect 33324 18634 33376 18640
rect 33508 18692 33560 18698
rect 33508 18634 33560 18640
rect 33232 18420 33284 18426
rect 33232 18362 33284 18368
rect 33048 18216 33100 18222
rect 33048 18158 33100 18164
rect 33060 17202 33088 18158
rect 33336 17610 33364 18634
rect 33520 18426 33548 18634
rect 33508 18420 33560 18426
rect 33508 18362 33560 18368
rect 33612 18086 33640 24670
rect 33888 22710 33916 29990
rect 34244 29096 34296 29102
rect 34244 29038 34296 29044
rect 33968 27872 34020 27878
rect 33968 27814 34020 27820
rect 33980 23866 34008 27814
rect 34256 27130 34284 29038
rect 34348 28762 34376 37198
rect 34520 37120 34572 37126
rect 34520 37062 34572 37068
rect 34428 36780 34480 36786
rect 34428 36722 34480 36728
rect 34440 36174 34468 36722
rect 34428 36168 34480 36174
rect 34428 36110 34480 36116
rect 34440 33998 34468 36110
rect 34532 36106 34560 37062
rect 35348 36780 35400 36786
rect 35348 36722 35400 36728
rect 34796 36576 34848 36582
rect 34796 36518 34848 36524
rect 34808 36242 34836 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35360 36378 35388 36722
rect 35440 36576 35492 36582
rect 35440 36518 35492 36524
rect 35348 36372 35400 36378
rect 35348 36314 35400 36320
rect 35452 36258 35480 36518
rect 34796 36236 34848 36242
rect 34796 36178 34848 36184
rect 35360 36230 35480 36258
rect 34888 36168 34940 36174
rect 34888 36110 34940 36116
rect 34520 36100 34572 36106
rect 34520 36042 34572 36048
rect 34428 33992 34480 33998
rect 34428 33934 34480 33940
rect 34336 28756 34388 28762
rect 34336 28698 34388 28704
rect 34532 28082 34560 36042
rect 34900 35834 34928 36110
rect 34888 35828 34940 35834
rect 34888 35770 34940 35776
rect 35360 35698 35388 36230
rect 35348 35692 35400 35698
rect 35348 35634 35400 35640
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34796 34740 34848 34746
rect 34796 34682 34848 34688
rect 34808 33658 34836 34682
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34796 33652 34848 33658
rect 34796 33594 34848 33600
rect 34808 30190 34836 33594
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35164 31748 35216 31754
rect 35164 31690 35216 31696
rect 35176 31414 35204 31690
rect 35164 31408 35216 31414
rect 35164 31350 35216 31356
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34796 30184 34848 30190
rect 34796 30126 34848 30132
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34624 29306 34652 29582
rect 34612 29300 34664 29306
rect 34612 29242 34664 29248
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 34624 27402 34652 29242
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28558 35388 35634
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 35452 31142 35480 31758
rect 35820 31754 35848 56306
rect 39868 55690 39896 57394
rect 40776 57384 40828 57390
rect 40776 57326 40828 57332
rect 40788 57050 40816 57326
rect 40776 57044 40828 57050
rect 40776 56986 40828 56992
rect 42536 56982 42564 57394
rect 42524 56976 42576 56982
rect 42524 56918 42576 56924
rect 42892 56364 42944 56370
rect 42892 56306 42944 56312
rect 43536 56364 43588 56370
rect 43536 56306 43588 56312
rect 43996 56364 44048 56370
rect 43996 56306 44048 56312
rect 39856 55684 39908 55690
rect 39856 55626 39908 55632
rect 42904 55622 42932 56306
rect 43548 55622 43576 56306
rect 44008 55622 44036 56306
rect 44100 56234 44128 57394
rect 44192 56506 44220 57394
rect 45468 56704 45520 56710
rect 45468 56646 45520 56652
rect 44180 56500 44232 56506
rect 44180 56442 44232 56448
rect 45480 56370 45508 56646
rect 46216 56506 46244 57462
rect 47584 57452 47636 57458
rect 47584 57394 47636 57400
rect 47676 57452 47728 57458
rect 47676 57394 47728 57400
rect 53472 57452 53524 57458
rect 53472 57394 53524 57400
rect 55312 57452 55364 57458
rect 55312 57394 55364 57400
rect 56048 57452 56100 57458
rect 56048 57394 56100 57400
rect 47596 56506 47624 57394
rect 46204 56500 46256 56506
rect 46204 56442 46256 56448
rect 47584 56500 47636 56506
rect 47584 56442 47636 56448
rect 44732 56364 44784 56370
rect 44732 56306 44784 56312
rect 45468 56364 45520 56370
rect 45468 56306 45520 56312
rect 46112 56364 46164 56370
rect 46112 56306 46164 56312
rect 46756 56364 46808 56370
rect 46756 56306 46808 56312
rect 44088 56228 44140 56234
rect 44088 56170 44140 56176
rect 44744 55622 44772 56306
rect 42892 55616 42944 55622
rect 42892 55558 42944 55564
rect 43536 55616 43588 55622
rect 43536 55558 43588 55564
rect 43996 55616 44048 55622
rect 43996 55558 44048 55564
rect 44732 55616 44784 55622
rect 44732 55558 44784 55564
rect 36728 37256 36780 37262
rect 36728 37198 36780 37204
rect 36740 36718 36768 37198
rect 36728 36712 36780 36718
rect 36728 36654 36780 36660
rect 36636 36168 36688 36174
rect 36636 36110 36688 36116
rect 35900 34536 35952 34542
rect 35900 34478 35952 34484
rect 35912 33590 35940 34478
rect 36268 34196 36320 34202
rect 36268 34138 36320 34144
rect 36176 33992 36228 33998
rect 36176 33934 36228 33940
rect 35900 33584 35952 33590
rect 35900 33526 35952 33532
rect 36188 33454 36216 33934
rect 36176 33448 36228 33454
rect 36176 33390 36228 33396
rect 35992 33312 36044 33318
rect 35992 33254 36044 33260
rect 35900 32224 35952 32230
rect 35900 32166 35952 32172
rect 35912 31958 35940 32166
rect 35900 31952 35952 31958
rect 35900 31894 35952 31900
rect 36004 31822 36032 33254
rect 36188 32434 36216 33390
rect 36176 32428 36228 32434
rect 36176 32370 36228 32376
rect 36084 31884 36136 31890
rect 36084 31826 36136 31832
rect 35992 31816 36044 31822
rect 35992 31758 36044 31764
rect 35728 31726 35848 31754
rect 35532 31408 35584 31414
rect 35532 31350 35584 31356
rect 35440 31136 35492 31142
rect 35440 31078 35492 31084
rect 35452 30122 35480 31078
rect 35544 30258 35572 31350
rect 35532 30252 35584 30258
rect 35532 30194 35584 30200
rect 35440 30116 35492 30122
rect 35440 30058 35492 30064
rect 35544 29510 35572 30194
rect 35624 29640 35676 29646
rect 35624 29582 35676 29588
rect 35532 29504 35584 29510
rect 35532 29446 35584 29452
rect 35544 29238 35572 29446
rect 35532 29232 35584 29238
rect 35532 29174 35584 29180
rect 35440 29164 35492 29170
rect 35440 29106 35492 29112
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 35452 28422 35480 29106
rect 35544 28558 35572 29174
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 34796 28416 34848 28422
rect 34796 28358 34848 28364
rect 35440 28416 35492 28422
rect 35440 28358 35492 28364
rect 34704 27532 34756 27538
rect 34704 27474 34756 27480
rect 34612 27396 34664 27402
rect 34612 27338 34664 27344
rect 34428 27328 34480 27334
rect 34428 27270 34480 27276
rect 34244 27124 34296 27130
rect 34244 27066 34296 27072
rect 34256 26994 34284 27066
rect 34440 26994 34468 27270
rect 34244 26988 34296 26994
rect 34244 26930 34296 26936
rect 34428 26988 34480 26994
rect 34428 26930 34480 26936
rect 34152 25832 34204 25838
rect 34152 25774 34204 25780
rect 34164 25294 34192 25774
rect 34152 25288 34204 25294
rect 34152 25230 34204 25236
rect 33968 23860 34020 23866
rect 33968 23802 34020 23808
rect 34164 23186 34192 25230
rect 34624 24750 34652 27338
rect 34716 26586 34744 27474
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34612 24744 34664 24750
rect 34612 24686 34664 24692
rect 34244 23656 34296 23662
rect 34244 23598 34296 23604
rect 34152 23180 34204 23186
rect 34152 23122 34204 23128
rect 34152 22976 34204 22982
rect 34152 22918 34204 22924
rect 33876 22704 33928 22710
rect 33876 22646 33928 22652
rect 34164 22642 34192 22918
rect 34152 22636 34204 22642
rect 34152 22578 34204 22584
rect 33784 22568 33836 22574
rect 33784 22510 33836 22516
rect 33692 22092 33744 22098
rect 33692 22034 33744 22040
rect 33600 18080 33652 18086
rect 33600 18022 33652 18028
rect 33416 17740 33468 17746
rect 33416 17682 33468 17688
rect 33324 17604 33376 17610
rect 33324 17546 33376 17552
rect 33428 17202 33456 17682
rect 33704 17678 33732 22034
rect 33692 17672 33744 17678
rect 33692 17614 33744 17620
rect 33600 17536 33652 17542
rect 33600 17478 33652 17484
rect 33612 17202 33640 17478
rect 33048 17196 33100 17202
rect 33048 17138 33100 17144
rect 33416 17196 33468 17202
rect 33416 17138 33468 17144
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33324 17060 33376 17066
rect 33324 17002 33376 17008
rect 33336 16794 33364 17002
rect 33324 16788 33376 16794
rect 33324 16730 33376 16736
rect 33324 15496 33376 15502
rect 33324 15438 33376 15444
rect 33336 15366 33364 15438
rect 33324 15360 33376 15366
rect 33324 15302 33376 15308
rect 33428 15026 33456 17138
rect 33704 16250 33732 17614
rect 33692 16244 33744 16250
rect 33692 16186 33744 16192
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 33600 15360 33652 15366
rect 33600 15302 33652 15308
rect 33416 15020 33468 15026
rect 33416 14962 33468 14968
rect 33140 13932 33192 13938
rect 33140 13874 33192 13880
rect 33152 13530 33180 13874
rect 33324 13728 33376 13734
rect 33324 13670 33376 13676
rect 33140 13524 33192 13530
rect 33140 13466 33192 13472
rect 33336 12918 33364 13670
rect 33612 13190 33640 15302
rect 33704 14958 33732 15438
rect 33692 14952 33744 14958
rect 33692 14894 33744 14900
rect 33600 13184 33652 13190
rect 33600 13126 33652 13132
rect 33140 12912 33192 12918
rect 33140 12854 33192 12860
rect 33324 12912 33376 12918
rect 33324 12854 33376 12860
rect 33152 9994 33180 12854
rect 33612 12850 33640 13126
rect 33600 12844 33652 12850
rect 33600 12786 33652 12792
rect 33416 12776 33468 12782
rect 33416 12718 33468 12724
rect 33428 11762 33456 12718
rect 33232 11756 33284 11762
rect 33232 11698 33284 11704
rect 33416 11756 33468 11762
rect 33416 11698 33468 11704
rect 33244 11218 33272 11698
rect 33232 11212 33284 11218
rect 33232 11154 33284 11160
rect 33796 10266 33824 22510
rect 33876 22432 33928 22438
rect 33876 22374 33928 22380
rect 33888 22234 33916 22374
rect 33876 22228 33928 22234
rect 33876 22170 33928 22176
rect 34152 20256 34204 20262
rect 34152 20198 34204 20204
rect 34164 19378 34192 20198
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 34164 18834 34192 19314
rect 34152 18828 34204 18834
rect 34152 18770 34204 18776
rect 34152 18284 34204 18290
rect 34152 18226 34204 18232
rect 34164 17746 34192 18226
rect 34152 17740 34204 17746
rect 34152 17682 34204 17688
rect 34060 16992 34112 16998
rect 34060 16934 34112 16940
rect 34072 16182 34100 16934
rect 34060 16176 34112 16182
rect 34060 16118 34112 16124
rect 33968 11620 34020 11626
rect 33968 11562 34020 11568
rect 33980 10810 34008 11562
rect 33968 10804 34020 10810
rect 33968 10746 34020 10752
rect 33784 10260 33836 10266
rect 33784 10202 33836 10208
rect 33140 9988 33192 9994
rect 33140 9930 33192 9936
rect 32956 9648 33008 9654
rect 32956 9590 33008 9596
rect 32588 9512 32640 9518
rect 32588 9454 32640 9460
rect 32600 8974 32628 9454
rect 33140 9376 33192 9382
rect 33140 9318 33192 9324
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32220 8900 32272 8906
rect 32220 8842 32272 8848
rect 33152 7478 33180 9318
rect 34256 9178 34284 23598
rect 34334 22536 34390 22545
rect 34334 22471 34336 22480
rect 34388 22471 34390 22480
rect 34336 22442 34388 22448
rect 34808 21622 34836 28358
rect 35452 28150 35480 28358
rect 35440 28144 35492 28150
rect 35440 28086 35492 28092
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35636 27062 35664 29582
rect 35624 27056 35676 27062
rect 35624 26998 35676 27004
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35624 23724 35676 23730
rect 35624 23666 35676 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35636 22778 35664 23666
rect 35624 22772 35676 22778
rect 35624 22714 35676 22720
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34796 21616 34848 21622
rect 34796 21558 34848 21564
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 34348 17882 34376 18158
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34336 17876 34388 17882
rect 34336 17818 34388 17824
rect 35728 17218 35756 31726
rect 36004 31414 36032 31758
rect 35992 31408 36044 31414
rect 35992 31350 36044 31356
rect 36004 30870 36032 31350
rect 36096 31346 36124 31826
rect 36176 31816 36228 31822
rect 36176 31758 36228 31764
rect 36188 31482 36216 31758
rect 36176 31476 36228 31482
rect 36176 31418 36228 31424
rect 36280 31346 36308 34138
rect 36360 31680 36412 31686
rect 36360 31622 36412 31628
rect 36372 31414 36400 31622
rect 36360 31408 36412 31414
rect 36360 31350 36412 31356
rect 36084 31340 36136 31346
rect 36084 31282 36136 31288
rect 36268 31340 36320 31346
rect 36268 31282 36320 31288
rect 35992 30864 36044 30870
rect 35992 30806 36044 30812
rect 36372 30802 36400 31350
rect 36360 30796 36412 30802
rect 36360 30738 36412 30744
rect 35992 30728 36044 30734
rect 35992 30670 36044 30676
rect 36004 30394 36032 30670
rect 35992 30388 36044 30394
rect 35992 30330 36044 30336
rect 36372 29714 36400 30738
rect 36648 30054 36676 36110
rect 36740 33998 36768 36654
rect 36728 33992 36780 33998
rect 36728 33934 36780 33940
rect 37280 33924 37332 33930
rect 37280 33866 37332 33872
rect 37292 33318 37320 33866
rect 37280 33312 37332 33318
rect 37280 33254 37332 33260
rect 36636 30048 36688 30054
rect 36636 29990 36688 29996
rect 36648 29850 36676 29990
rect 36636 29844 36688 29850
rect 36636 29786 36688 29792
rect 36360 29708 36412 29714
rect 36360 29650 36412 29656
rect 36084 29640 36136 29646
rect 36084 29582 36136 29588
rect 36096 29170 36124 29582
rect 36268 29300 36320 29306
rect 36268 29242 36320 29248
rect 36084 29164 36136 29170
rect 36084 29106 36136 29112
rect 36280 28558 36308 29242
rect 36372 29050 36400 29650
rect 37004 29640 37056 29646
rect 37004 29582 37056 29588
rect 36544 29164 36596 29170
rect 36544 29106 36596 29112
rect 36372 29034 36492 29050
rect 36372 29028 36504 29034
rect 36372 29022 36452 29028
rect 36452 28970 36504 28976
rect 36556 28966 36584 29106
rect 36360 28960 36412 28966
rect 36360 28902 36412 28908
rect 36544 28960 36596 28966
rect 36544 28902 36596 28908
rect 36372 28762 36400 28902
rect 37016 28762 37044 29582
rect 36360 28756 36412 28762
rect 36360 28698 36412 28704
rect 37004 28756 37056 28762
rect 37004 28698 37056 28704
rect 36268 28552 36320 28558
rect 36268 28494 36320 28500
rect 35808 26784 35860 26790
rect 35808 26726 35860 26732
rect 37096 26784 37148 26790
rect 37096 26726 37148 26732
rect 35820 26382 35848 26726
rect 35808 26376 35860 26382
rect 35808 26318 35860 26324
rect 36176 25152 36228 25158
rect 36176 25094 36228 25100
rect 36188 24750 36216 25094
rect 36176 24744 36228 24750
rect 36176 24686 36228 24692
rect 36084 23792 36136 23798
rect 36084 23734 36136 23740
rect 35808 23724 35860 23730
rect 35808 23666 35860 23672
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 35820 23186 35848 23666
rect 35900 23520 35952 23526
rect 35900 23462 35952 23468
rect 35808 23180 35860 23186
rect 35808 23122 35860 23128
rect 35820 22642 35848 23122
rect 35912 22710 35940 23462
rect 36004 23050 36032 23666
rect 36096 23254 36124 23734
rect 36188 23730 36216 24686
rect 36176 23724 36228 23730
rect 36176 23666 36228 23672
rect 36084 23248 36136 23254
rect 36084 23190 36136 23196
rect 35992 23044 36044 23050
rect 35992 22986 36044 22992
rect 35900 22704 35952 22710
rect 35900 22646 35952 22652
rect 36004 22642 36032 22986
rect 36096 22710 36124 23190
rect 36084 22704 36136 22710
rect 36084 22646 36136 22652
rect 37108 22642 37136 26726
rect 37188 26376 37240 26382
rect 37188 26318 37240 26324
rect 37200 25770 37228 26318
rect 37292 26042 37320 33254
rect 37464 32428 37516 32434
rect 37464 32370 37516 32376
rect 37556 32428 37608 32434
rect 37556 32370 37608 32376
rect 37476 31346 37504 32370
rect 37568 32026 37596 32370
rect 38660 32224 38712 32230
rect 38660 32166 38712 32172
rect 37556 32020 37608 32026
rect 37556 31962 37608 31968
rect 38672 31346 38700 32166
rect 37464 31340 37516 31346
rect 37464 31282 37516 31288
rect 37924 31340 37976 31346
rect 37924 31282 37976 31288
rect 38660 31340 38712 31346
rect 38660 31282 38712 31288
rect 37936 30802 37964 31282
rect 37924 30796 37976 30802
rect 37924 30738 37976 30744
rect 37372 30592 37424 30598
rect 37372 30534 37424 30540
rect 37384 30326 37412 30534
rect 37372 30320 37424 30326
rect 37372 30262 37424 30268
rect 37464 29504 37516 29510
rect 37464 29446 37516 29452
rect 37476 29238 37504 29446
rect 37464 29232 37516 29238
rect 37464 29174 37516 29180
rect 39488 29096 39540 29102
rect 39488 29038 39540 29044
rect 38384 29028 38436 29034
rect 38384 28970 38436 28976
rect 38396 28558 38424 28970
rect 39500 28558 39528 29038
rect 38384 28552 38436 28558
rect 38384 28494 38436 28500
rect 39488 28552 39540 28558
rect 39488 28494 39540 28500
rect 39948 28552 40000 28558
rect 39948 28494 40000 28500
rect 39856 28076 39908 28082
rect 39856 28018 39908 28024
rect 39028 27872 39080 27878
rect 39080 27820 39160 27826
rect 39028 27814 39160 27820
rect 39040 27798 39160 27814
rect 37372 26376 37424 26382
rect 37372 26318 37424 26324
rect 37280 26036 37332 26042
rect 37280 25978 37332 25984
rect 37188 25764 37240 25770
rect 37188 25706 37240 25712
rect 37200 25294 37228 25706
rect 37188 25288 37240 25294
rect 37188 25230 37240 25236
rect 37200 23118 37228 25230
rect 37384 24818 37412 26318
rect 39132 26314 39160 27798
rect 39120 26308 39172 26314
rect 39120 26250 39172 26256
rect 37832 25696 37884 25702
rect 37832 25638 37884 25644
rect 37844 25294 37872 25638
rect 37832 25288 37884 25294
rect 38016 25288 38068 25294
rect 37884 25248 37964 25276
rect 37832 25230 37884 25236
rect 37372 24812 37424 24818
rect 37372 24754 37424 24760
rect 37188 23112 37240 23118
rect 37188 23054 37240 23060
rect 37384 22642 37412 24754
rect 37936 23662 37964 25248
rect 38016 25230 38068 25236
rect 38028 24954 38056 25230
rect 38016 24948 38068 24954
rect 38016 24890 38068 24896
rect 38752 24608 38804 24614
rect 38752 24550 38804 24556
rect 38764 24206 38792 24550
rect 38752 24200 38804 24206
rect 38752 24142 38804 24148
rect 37924 23656 37976 23662
rect 37924 23598 37976 23604
rect 37936 23118 37964 23598
rect 38384 23588 38436 23594
rect 38384 23530 38436 23536
rect 38396 23118 38424 23530
rect 37924 23112 37976 23118
rect 37924 23054 37976 23060
rect 38200 23112 38252 23118
rect 38200 23054 38252 23060
rect 38384 23112 38436 23118
rect 38384 23054 38436 23060
rect 35808 22636 35860 22642
rect 35808 22578 35860 22584
rect 35992 22636 36044 22642
rect 35992 22578 36044 22584
rect 37096 22636 37148 22642
rect 37096 22578 37148 22584
rect 37372 22636 37424 22642
rect 37372 22578 37424 22584
rect 35820 19378 35848 22578
rect 36268 22568 36320 22574
rect 36268 22510 36320 22516
rect 36280 19922 36308 22510
rect 37832 22228 37884 22234
rect 37832 22170 37884 22176
rect 37280 21412 37332 21418
rect 37280 21354 37332 21360
rect 37292 20602 37320 21354
rect 37464 20800 37516 20806
rect 37464 20742 37516 20748
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 37372 20528 37424 20534
rect 37372 20470 37424 20476
rect 37280 20460 37332 20466
rect 37280 20402 37332 20408
rect 36268 19916 36320 19922
rect 36268 19858 36320 19864
rect 36084 19712 36136 19718
rect 36084 19654 36136 19660
rect 36096 19446 36124 19654
rect 36280 19446 36308 19858
rect 36084 19440 36136 19446
rect 36084 19382 36136 19388
rect 36268 19440 36320 19446
rect 36268 19382 36320 19388
rect 35808 19372 35860 19378
rect 35808 19314 35860 19320
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 36004 18766 36032 19314
rect 36280 18766 36308 19382
rect 37292 19310 37320 20402
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37292 18766 37320 19246
rect 37384 18970 37412 20470
rect 37476 19854 37504 20742
rect 37648 20528 37700 20534
rect 37648 20470 37700 20476
rect 37556 20460 37608 20466
rect 37556 20402 37608 20408
rect 37464 19848 37516 19854
rect 37464 19790 37516 19796
rect 37372 18964 37424 18970
rect 37372 18906 37424 18912
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 36912 18760 36964 18766
rect 36912 18702 36964 18708
rect 37280 18760 37332 18766
rect 37280 18702 37332 18708
rect 36268 17604 36320 17610
rect 36268 17546 36320 17552
rect 36176 17536 36228 17542
rect 36176 17478 36228 17484
rect 35624 17196 35676 17202
rect 35728 17190 35848 17218
rect 35624 17138 35676 17144
rect 34520 17128 34572 17134
rect 34520 17070 34572 17076
rect 34532 16046 34560 17070
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35636 16794 35664 17138
rect 35624 16788 35676 16794
rect 35624 16730 35676 16736
rect 35624 16584 35676 16590
rect 35624 16526 35676 16532
rect 34520 16040 34572 16046
rect 34520 15982 34572 15988
rect 35532 16040 35584 16046
rect 35532 15982 35584 15988
rect 34532 14278 34560 15982
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35440 15428 35492 15434
rect 35440 15370 35492 15376
rect 35452 15026 35480 15370
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35440 14884 35492 14890
rect 35440 14826 35492 14832
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35164 14408 35216 14414
rect 35164 14350 35216 14356
rect 35348 14408 35400 14414
rect 35348 14350 35400 14356
rect 34520 14272 34572 14278
rect 34520 14214 34572 14220
rect 34532 13920 34560 14214
rect 35176 13938 35204 14350
rect 34612 13932 34664 13938
rect 34532 13892 34612 13920
rect 34532 12238 34560 13892
rect 34612 13874 34664 13880
rect 35164 13932 35216 13938
rect 35164 13874 35216 13880
rect 35360 13802 35388 14350
rect 35452 13938 35480 14826
rect 35544 14482 35572 15982
rect 35532 14476 35584 14482
rect 35532 14418 35584 14424
rect 35440 13932 35492 13938
rect 35440 13874 35492 13880
rect 35348 13796 35400 13802
rect 35348 13738 35400 13744
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35360 13394 35388 13738
rect 35348 13388 35400 13394
rect 35348 13330 35400 13336
rect 34704 13252 34756 13258
rect 34704 13194 34756 13200
rect 34520 12232 34572 12238
rect 34520 12174 34572 12180
rect 34532 11218 34560 12174
rect 34612 12096 34664 12102
rect 34612 12038 34664 12044
rect 34520 11212 34572 11218
rect 34520 11154 34572 11160
rect 34244 9172 34296 9178
rect 34244 9114 34296 9120
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 33140 7472 33192 7478
rect 33140 7414 33192 7420
rect 33888 7410 33916 7822
rect 33876 7404 33928 7410
rect 33876 7346 33928 7352
rect 33888 5914 33916 7346
rect 34624 6746 34652 12038
rect 34716 11898 34744 13194
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34704 11892 34756 11898
rect 34704 11834 34756 11840
rect 35360 11762 35388 13330
rect 35452 12434 35480 13874
rect 35636 12442 35664 16526
rect 35716 13320 35768 13326
rect 35716 13262 35768 13268
rect 35728 12850 35756 13262
rect 35716 12844 35768 12850
rect 35716 12786 35768 12792
rect 35624 12436 35676 12442
rect 35452 12406 35572 12434
rect 35544 11762 35572 12406
rect 35624 12378 35676 12384
rect 35728 11778 35756 12786
rect 35820 12102 35848 17190
rect 36188 16590 36216 17478
rect 36280 17338 36308 17546
rect 36268 17332 36320 17338
rect 36268 17274 36320 17280
rect 36360 16992 36412 16998
rect 36360 16934 36412 16940
rect 36372 16590 36400 16934
rect 36176 16584 36228 16590
rect 36176 16526 36228 16532
rect 36360 16584 36412 16590
rect 36360 16526 36412 16532
rect 36176 15700 36228 15706
rect 36176 15642 36228 15648
rect 35992 14816 36044 14822
rect 35992 14758 36044 14764
rect 36004 14074 36032 14758
rect 36188 14414 36216 15642
rect 36728 15020 36780 15026
rect 36728 14962 36780 14968
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 35900 13864 35952 13870
rect 35900 13806 35952 13812
rect 35912 13530 35940 13806
rect 35900 13524 35952 13530
rect 35900 13466 35952 13472
rect 35912 12986 35940 13466
rect 36004 13326 36032 14010
rect 36740 13326 36768 14962
rect 35992 13320 36044 13326
rect 35992 13262 36044 13268
rect 36728 13320 36780 13326
rect 36728 13262 36780 13268
rect 36360 13184 36412 13190
rect 36360 13126 36412 13132
rect 35900 12980 35952 12986
rect 35900 12922 35952 12928
rect 36372 12850 36400 13126
rect 36740 12986 36768 13262
rect 36728 12980 36780 12986
rect 36728 12922 36780 12928
rect 36360 12844 36412 12850
rect 36360 12786 36412 12792
rect 36544 12844 36596 12850
rect 36544 12786 36596 12792
rect 36556 12442 36584 12786
rect 36728 12640 36780 12646
rect 36728 12582 36780 12588
rect 36544 12436 36596 12442
rect 36544 12378 36596 12384
rect 36740 12170 36768 12582
rect 36728 12164 36780 12170
rect 36728 12106 36780 12112
rect 35808 12096 35860 12102
rect 35808 12038 35860 12044
rect 36268 11824 36320 11830
rect 35348 11756 35400 11762
rect 35348 11698 35400 11704
rect 35532 11756 35584 11762
rect 35532 11698 35584 11704
rect 35624 11756 35676 11762
rect 35728 11750 35848 11778
rect 36268 11766 36320 11772
rect 35624 11698 35676 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35164 11076 35216 11082
rect 35164 11018 35216 11024
rect 35176 10810 35204 11018
rect 35164 10804 35216 10810
rect 35164 10746 35216 10752
rect 34796 10668 34848 10674
rect 34796 10610 34848 10616
rect 34704 9512 34756 9518
rect 34704 9454 34756 9460
rect 34716 8362 34744 9454
rect 34808 8974 34836 10610
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35440 9920 35492 9926
rect 35440 9862 35492 9868
rect 35348 9648 35400 9654
rect 35348 9590 35400 9596
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 35360 9178 35388 9590
rect 35348 9172 35400 9178
rect 35348 9114 35400 9120
rect 35452 9110 35480 9862
rect 35440 9104 35492 9110
rect 35440 9046 35492 9052
rect 34796 8968 34848 8974
rect 34796 8910 34848 8916
rect 34808 8566 34836 8910
rect 35348 8832 35400 8838
rect 35544 8786 35572 11698
rect 35636 10062 35664 11698
rect 35716 11620 35768 11626
rect 35716 11562 35768 11568
rect 35624 10056 35676 10062
rect 35624 9998 35676 10004
rect 35636 9382 35664 9998
rect 35624 9376 35676 9382
rect 35624 9318 35676 9324
rect 35624 8968 35676 8974
rect 35624 8910 35676 8916
rect 35348 8774 35400 8780
rect 34796 8560 34848 8566
rect 34796 8502 34848 8508
rect 34704 8356 34756 8362
rect 34704 8298 34756 8304
rect 34532 6718 34652 6746
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 32128 5636 32180 5642
rect 32128 5578 32180 5584
rect 32140 4758 32168 5578
rect 32128 4752 32180 4758
rect 32128 4694 32180 4700
rect 33888 4146 33916 5850
rect 33876 4140 33928 4146
rect 33876 4082 33928 4088
rect 32036 3732 32088 3738
rect 32036 3674 32088 3680
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30840 3528 30892 3534
rect 30840 3470 30892 3476
rect 34532 3058 34560 6718
rect 34612 6656 34664 6662
rect 34612 6598 34664 6604
rect 34624 4162 34652 6598
rect 34716 6322 34744 8298
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35256 7404 35308 7410
rect 35360 7392 35388 8774
rect 35452 8758 35572 8786
rect 35452 7818 35480 8758
rect 35636 8650 35664 8910
rect 35544 8622 35664 8650
rect 35544 8430 35572 8622
rect 35532 8424 35584 8430
rect 35532 8366 35584 8372
rect 35440 7812 35492 7818
rect 35440 7754 35492 7760
rect 35452 7478 35480 7754
rect 35440 7472 35492 7478
rect 35440 7414 35492 7420
rect 35544 7410 35572 8366
rect 35624 7880 35676 7886
rect 35624 7822 35676 7828
rect 35308 7364 35388 7392
rect 35256 7346 35308 7352
rect 34796 7200 34848 7206
rect 34796 7142 34848 7148
rect 34808 6390 34836 7142
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6848 35388 7364
rect 35532 7404 35584 7410
rect 35532 7346 35584 7352
rect 35440 6860 35492 6866
rect 35360 6820 35440 6848
rect 35440 6802 35492 6808
rect 35544 6798 35572 7346
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35348 6656 35400 6662
rect 35348 6598 35400 6604
rect 34796 6384 34848 6390
rect 34796 6326 34848 6332
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 35360 5914 35388 6598
rect 35348 5908 35400 5914
rect 35348 5850 35400 5856
rect 35636 5710 35664 7822
rect 35728 7750 35756 11562
rect 35820 8974 35848 11750
rect 36280 11354 36308 11766
rect 36268 11348 36320 11354
rect 36268 11290 36320 11296
rect 36280 10742 36308 11290
rect 36268 10736 36320 10742
rect 36268 10678 36320 10684
rect 36924 8974 36952 18702
rect 37188 18216 37240 18222
rect 37188 18158 37240 18164
rect 37200 17610 37228 18158
rect 37188 17604 37240 17610
rect 37188 17546 37240 17552
rect 37004 16584 37056 16590
rect 37004 16526 37056 16532
rect 37016 16114 37044 16526
rect 37004 16108 37056 16114
rect 37004 16050 37056 16056
rect 37200 15434 37228 17546
rect 37292 16114 37320 18702
rect 37372 17332 37424 17338
rect 37372 17274 37424 17280
rect 37384 16590 37412 17274
rect 37372 16584 37424 16590
rect 37372 16526 37424 16532
rect 37372 16448 37424 16454
rect 37372 16390 37424 16396
rect 37280 16108 37332 16114
rect 37280 16050 37332 16056
rect 37278 16008 37334 16017
rect 37278 15943 37280 15952
rect 37332 15943 37334 15952
rect 37280 15914 37332 15920
rect 37188 15428 37240 15434
rect 37188 15370 37240 15376
rect 37200 14006 37228 15370
rect 37188 14000 37240 14006
rect 37188 13942 37240 13948
rect 37200 13852 37228 13942
rect 37280 13864 37332 13870
rect 37200 13824 37280 13852
rect 37280 13806 37332 13812
rect 37280 13252 37332 13258
rect 37280 13194 37332 13200
rect 37292 10062 37320 13194
rect 37384 12918 37412 16390
rect 37476 15706 37504 19790
rect 37568 19514 37596 20402
rect 37660 19786 37688 20470
rect 37844 20466 37872 22170
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37648 19780 37700 19786
rect 37648 19722 37700 19728
rect 37556 19508 37608 19514
rect 37556 19450 37608 19456
rect 37660 18698 37688 19722
rect 37648 18692 37700 18698
rect 37648 18634 37700 18640
rect 37660 16522 37688 18634
rect 37936 18426 37964 23054
rect 38212 22778 38240 23054
rect 38200 22772 38252 22778
rect 38200 22714 38252 22720
rect 38108 22636 38160 22642
rect 38108 22578 38160 22584
rect 38292 22636 38344 22642
rect 38292 22578 38344 22584
rect 38016 19440 38068 19446
rect 38016 19382 38068 19388
rect 37924 18420 37976 18426
rect 37924 18362 37976 18368
rect 37832 17604 37884 17610
rect 37832 17546 37884 17552
rect 37844 16658 37872 17546
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 37648 16516 37700 16522
rect 37648 16458 37700 16464
rect 37660 16114 37688 16458
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 37464 15700 37516 15706
rect 37464 15642 37516 15648
rect 37660 15570 37688 16050
rect 37844 15638 37872 16594
rect 37832 15632 37884 15638
rect 37832 15574 37884 15580
rect 37648 15564 37700 15570
rect 37648 15506 37700 15512
rect 37844 15094 37872 15574
rect 37832 15088 37884 15094
rect 37832 15030 37884 15036
rect 37648 14884 37700 14890
rect 37648 14826 37700 14832
rect 37660 14006 37688 14826
rect 37740 14612 37792 14618
rect 37740 14554 37792 14560
rect 37648 14000 37700 14006
rect 37648 13942 37700 13948
rect 37556 13864 37608 13870
rect 37556 13806 37608 13812
rect 37568 13258 37596 13806
rect 37556 13252 37608 13258
rect 37556 13194 37608 13200
rect 37372 12912 37424 12918
rect 37424 12860 37504 12866
rect 37372 12854 37504 12860
rect 37384 12838 37504 12854
rect 37476 12442 37504 12838
rect 37464 12436 37516 12442
rect 37464 12378 37516 12384
rect 37280 10056 37332 10062
rect 37280 9998 37332 10004
rect 35808 8968 35860 8974
rect 35808 8910 35860 8916
rect 36912 8968 36964 8974
rect 36912 8910 36964 8916
rect 36084 8288 36136 8294
rect 36084 8230 36136 8236
rect 36096 8090 36124 8230
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 35716 7744 35768 7750
rect 35716 7686 35768 7692
rect 35728 7410 35756 7686
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 36096 6882 36124 8026
rect 36924 8022 36952 8910
rect 37292 8906 37320 9998
rect 37556 9376 37608 9382
rect 37556 9318 37608 9324
rect 37568 8974 37596 9318
rect 37660 9042 37688 13942
rect 37752 13734 37780 14554
rect 37740 13728 37792 13734
rect 37740 13670 37792 13676
rect 37752 12918 37780 13670
rect 38028 13326 38056 19382
rect 38120 18698 38148 22578
rect 38304 22234 38332 22578
rect 38292 22228 38344 22234
rect 38292 22170 38344 22176
rect 38108 18692 38160 18698
rect 38108 18634 38160 18640
rect 38120 18290 38148 18634
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 38200 16992 38252 16998
rect 38200 16934 38252 16940
rect 38212 15502 38240 16934
rect 38200 15496 38252 15502
rect 38200 15438 38252 15444
rect 38016 13320 38068 13326
rect 38016 13262 38068 13268
rect 38028 12986 38056 13262
rect 38016 12980 38068 12986
rect 38016 12922 38068 12928
rect 37740 12912 37792 12918
rect 37740 12854 37792 12860
rect 37752 11762 37780 12854
rect 38396 12434 38424 23054
rect 38764 22982 38792 24142
rect 39132 23322 39160 26250
rect 39868 25498 39896 28018
rect 39960 28014 39988 28494
rect 39948 28008 40000 28014
rect 39948 27950 40000 27956
rect 39960 26926 39988 27950
rect 40500 26988 40552 26994
rect 40500 26930 40552 26936
rect 39948 26920 40000 26926
rect 39948 26862 40000 26868
rect 39960 25770 39988 26862
rect 40040 26784 40092 26790
rect 40040 26726 40092 26732
rect 40052 26314 40080 26726
rect 40316 26376 40368 26382
rect 40316 26318 40368 26324
rect 40040 26308 40092 26314
rect 40040 26250 40092 26256
rect 39948 25764 40000 25770
rect 39948 25706 40000 25712
rect 39856 25492 39908 25498
rect 39856 25434 39908 25440
rect 39764 25220 39816 25226
rect 39764 25162 39816 25168
rect 39120 23316 39172 23322
rect 39120 23258 39172 23264
rect 38752 22976 38804 22982
rect 38752 22918 38804 22924
rect 38936 22432 38988 22438
rect 38936 22374 38988 22380
rect 38844 22024 38896 22030
rect 38764 21972 38844 21978
rect 38764 21966 38896 21972
rect 38476 21956 38528 21962
rect 38476 21898 38528 21904
rect 38764 21950 38884 21966
rect 38488 21690 38516 21898
rect 38476 21684 38528 21690
rect 38476 21626 38528 21632
rect 38660 21548 38712 21554
rect 38660 21490 38712 21496
rect 38672 20058 38700 21490
rect 38764 20398 38792 21950
rect 38948 21554 38976 22374
rect 39776 21554 39804 25162
rect 39960 24834 39988 25706
rect 40132 25424 40184 25430
rect 40132 25366 40184 25372
rect 40144 25294 40172 25366
rect 40328 25294 40356 26318
rect 40512 25498 40540 26930
rect 41144 26240 41196 26246
rect 41144 26182 41196 26188
rect 40500 25492 40552 25498
rect 40500 25434 40552 25440
rect 40868 25356 40920 25362
rect 40868 25298 40920 25304
rect 40132 25288 40184 25294
rect 40132 25230 40184 25236
rect 40316 25288 40368 25294
rect 40316 25230 40368 25236
rect 40144 24970 40172 25230
rect 40144 24942 40356 24970
rect 39960 24818 40080 24834
rect 39960 24812 40092 24818
rect 39960 24806 40040 24812
rect 39960 23746 39988 24806
rect 40040 24754 40092 24760
rect 40224 24812 40276 24818
rect 40224 24754 40276 24760
rect 40132 24132 40184 24138
rect 40132 24074 40184 24080
rect 39960 23730 40080 23746
rect 39960 23724 40092 23730
rect 39960 23718 40040 23724
rect 40040 23666 40092 23672
rect 40144 22710 40172 24074
rect 40236 23322 40264 24754
rect 40224 23316 40276 23322
rect 40224 23258 40276 23264
rect 40328 23100 40356 24942
rect 40408 24132 40460 24138
rect 40408 24074 40460 24080
rect 40420 23526 40448 24074
rect 40408 23520 40460 23526
rect 40408 23462 40460 23468
rect 40408 23112 40460 23118
rect 40328 23072 40408 23100
rect 40328 22778 40356 23072
rect 40408 23054 40460 23060
rect 40316 22772 40368 22778
rect 40316 22714 40368 22720
rect 40132 22704 40184 22710
rect 40132 22646 40184 22652
rect 40592 22704 40644 22710
rect 40592 22646 40644 22652
rect 38936 21548 38988 21554
rect 38936 21490 38988 21496
rect 39764 21548 39816 21554
rect 39764 21490 39816 21496
rect 38752 20392 38804 20398
rect 38752 20334 38804 20340
rect 38660 20052 38712 20058
rect 38660 19994 38712 20000
rect 38764 19718 38792 20334
rect 38752 19712 38804 19718
rect 38752 19654 38804 19660
rect 38764 19310 38792 19654
rect 38752 19304 38804 19310
rect 38752 19246 38804 19252
rect 38764 18222 38792 19246
rect 39396 18624 39448 18630
rect 39396 18566 39448 18572
rect 38752 18216 38804 18222
rect 38752 18158 38804 18164
rect 38660 18148 38712 18154
rect 38660 18090 38712 18096
rect 38672 17746 38700 18090
rect 38660 17740 38712 17746
rect 38660 17682 38712 17688
rect 38568 16244 38620 16250
rect 38568 16186 38620 16192
rect 38580 15502 38608 16186
rect 38764 16114 38792 18158
rect 38936 17672 38988 17678
rect 38936 17614 38988 17620
rect 38948 16590 38976 17614
rect 38936 16584 38988 16590
rect 38936 16526 38988 16532
rect 38660 16108 38712 16114
rect 38660 16050 38712 16056
rect 38752 16108 38804 16114
rect 38752 16050 38804 16056
rect 38568 15496 38620 15502
rect 38568 15438 38620 15444
rect 38672 15434 38700 16050
rect 38660 15428 38712 15434
rect 38660 15370 38712 15376
rect 38672 15162 38700 15370
rect 38844 15360 38896 15366
rect 38844 15302 38896 15308
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38856 15094 38884 15302
rect 38844 15088 38896 15094
rect 38844 15030 38896 15036
rect 38660 14952 38712 14958
rect 38660 14894 38712 14900
rect 38672 14278 38700 14894
rect 38948 14618 38976 16526
rect 38936 14612 38988 14618
rect 38936 14554 38988 14560
rect 38936 14476 38988 14482
rect 38936 14418 38988 14424
rect 38660 14272 38712 14278
rect 38660 14214 38712 14220
rect 38672 12850 38700 14214
rect 38948 13938 38976 14418
rect 38752 13932 38804 13938
rect 38752 13874 38804 13880
rect 38936 13932 38988 13938
rect 38936 13874 38988 13880
rect 38764 13530 38792 13874
rect 38752 13524 38804 13530
rect 38752 13466 38804 13472
rect 38660 12844 38712 12850
rect 38660 12786 38712 12792
rect 38120 12406 38424 12434
rect 37740 11756 37792 11762
rect 37740 11698 37792 11704
rect 38120 11558 38148 12406
rect 38384 12232 38436 12238
rect 38384 12174 38436 12180
rect 38292 11688 38344 11694
rect 38292 11630 38344 11636
rect 38108 11552 38160 11558
rect 38108 11494 38160 11500
rect 38120 11354 38148 11494
rect 38108 11348 38160 11354
rect 38108 11290 38160 11296
rect 38304 11082 38332 11630
rect 38292 11076 38344 11082
rect 38292 11018 38344 11024
rect 38304 10674 38332 11018
rect 38292 10668 38344 10674
rect 38292 10610 38344 10616
rect 38304 9994 38332 10610
rect 38396 10606 38424 12174
rect 38948 11150 38976 13874
rect 39212 13728 39264 13734
rect 39212 13670 39264 13676
rect 39224 12918 39252 13670
rect 39212 12912 39264 12918
rect 39212 12854 39264 12860
rect 39120 11620 39172 11626
rect 39120 11562 39172 11568
rect 39132 11286 39160 11562
rect 39304 11348 39356 11354
rect 39304 11290 39356 11296
rect 39120 11280 39172 11286
rect 39120 11222 39172 11228
rect 38936 11144 38988 11150
rect 38936 11086 38988 11092
rect 38660 11008 38712 11014
rect 38660 10950 38712 10956
rect 38672 10742 38700 10950
rect 38660 10736 38712 10742
rect 38660 10678 38712 10684
rect 38384 10600 38436 10606
rect 38384 10542 38436 10548
rect 38292 9988 38344 9994
rect 38292 9930 38344 9936
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 37648 9036 37700 9042
rect 37648 8978 37700 8984
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 37280 8900 37332 8906
rect 37332 8860 37412 8888
rect 37280 8842 37332 8848
rect 37096 8832 37148 8838
rect 37096 8774 37148 8780
rect 37108 8566 37136 8774
rect 37096 8560 37148 8566
rect 37096 8502 37148 8508
rect 37278 8528 37334 8537
rect 37278 8463 37280 8472
rect 37332 8463 37334 8472
rect 37280 8434 37332 8440
rect 37292 8090 37320 8434
rect 37280 8084 37332 8090
rect 37280 8026 37332 8032
rect 36912 8016 36964 8022
rect 36912 7958 36964 7964
rect 36268 7404 36320 7410
rect 36268 7346 36320 7352
rect 37096 7404 37148 7410
rect 37096 7346 37148 7352
rect 36176 7268 36228 7274
rect 36176 7210 36228 7216
rect 35912 6854 36124 6882
rect 35912 6730 35940 6854
rect 36188 6798 36216 7210
rect 35992 6792 36044 6798
rect 35992 6734 36044 6740
rect 36176 6792 36228 6798
rect 36176 6734 36228 6740
rect 35900 6724 35952 6730
rect 35900 6666 35952 6672
rect 36004 5914 36032 6734
rect 36084 6656 36136 6662
rect 36084 6598 36136 6604
rect 36096 6322 36124 6598
rect 36188 6390 36216 6734
rect 36176 6384 36228 6390
rect 36176 6326 36228 6332
rect 36084 6316 36136 6322
rect 36084 6258 36136 6264
rect 35992 5908 36044 5914
rect 35992 5850 36044 5856
rect 36280 5710 36308 7346
rect 36912 7336 36964 7342
rect 36912 7278 36964 7284
rect 36924 7002 36952 7278
rect 36912 6996 36964 7002
rect 36912 6938 36964 6944
rect 37004 6928 37056 6934
rect 37004 6870 37056 6876
rect 37016 6798 37044 6870
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 37108 6730 37136 7346
rect 37384 6730 37412 8860
rect 37568 8634 37596 8910
rect 37556 8628 37608 8634
rect 37556 8570 37608 8576
rect 37660 8480 37688 8978
rect 37936 8838 37964 9454
rect 37924 8832 37976 8838
rect 37924 8774 37976 8780
rect 37740 8492 37792 8498
rect 37660 8452 37740 8480
rect 37740 8434 37792 8440
rect 37936 8362 37964 8774
rect 37924 8356 37976 8362
rect 37924 8298 37976 8304
rect 37936 7954 37964 8298
rect 38200 8288 38252 8294
rect 38200 8230 38252 8236
rect 37924 7948 37976 7954
rect 37924 7890 37976 7896
rect 37096 6724 37148 6730
rect 37096 6666 37148 6672
rect 37372 6724 37424 6730
rect 37372 6666 37424 6672
rect 37108 6458 37136 6666
rect 37096 6452 37148 6458
rect 37096 6394 37148 6400
rect 35624 5704 35676 5710
rect 35624 5646 35676 5652
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34624 4146 34744 4162
rect 34624 4140 34756 4146
rect 34624 4134 34704 4140
rect 34704 4082 34756 4088
rect 35636 4010 35664 5646
rect 36280 5370 36308 5646
rect 37384 5574 37412 6666
rect 37936 6322 37964 7890
rect 38212 7886 38240 8230
rect 38200 7880 38252 7886
rect 38200 7822 38252 7828
rect 38304 7410 38332 9930
rect 38396 9518 38424 10542
rect 39132 10470 39160 11222
rect 39316 11150 39344 11290
rect 39304 11144 39356 11150
rect 39304 11086 39356 11092
rect 39120 10464 39172 10470
rect 39120 10406 39172 10412
rect 38752 9920 38804 9926
rect 38752 9862 38804 9868
rect 38660 9580 38712 9586
rect 38660 9522 38712 9528
rect 38384 9512 38436 9518
rect 38384 9454 38436 9460
rect 38672 8634 38700 9522
rect 38660 8628 38712 8634
rect 38660 8570 38712 8576
rect 38764 8566 38792 9862
rect 38752 8560 38804 8566
rect 38752 8502 38804 8508
rect 38842 8528 38898 8537
rect 38842 8463 38844 8472
rect 38896 8463 38898 8472
rect 38844 8434 38896 8440
rect 39132 8430 39160 10406
rect 39316 8498 39344 11086
rect 39408 10062 39436 18566
rect 39776 14074 39804 21490
rect 40040 21480 40092 21486
rect 40040 21422 40092 21428
rect 40052 17814 40080 21422
rect 40224 20936 40276 20942
rect 40224 20878 40276 20884
rect 40236 20262 40264 20878
rect 40500 20868 40552 20874
rect 40500 20810 40552 20816
rect 40512 20754 40540 20810
rect 40604 20754 40632 22646
rect 40880 21486 40908 25298
rect 41156 25294 41184 26182
rect 41144 25288 41196 25294
rect 41144 25230 41196 25236
rect 41236 25152 41288 25158
rect 41236 25094 41288 25100
rect 41248 24614 41276 25094
rect 41236 24608 41288 24614
rect 41236 24550 41288 24556
rect 40960 24064 41012 24070
rect 41012 24024 41092 24052
rect 40960 24006 41012 24012
rect 41064 23730 41092 24024
rect 41248 23866 41276 24550
rect 41420 24064 41472 24070
rect 41420 24006 41472 24012
rect 41236 23860 41288 23866
rect 41236 23802 41288 23808
rect 41052 23724 41104 23730
rect 41052 23666 41104 23672
rect 40960 23588 41012 23594
rect 40960 23530 41012 23536
rect 41052 23588 41104 23594
rect 41052 23530 41104 23536
rect 40972 23050 41000 23530
rect 41064 23118 41092 23530
rect 41052 23112 41104 23118
rect 41052 23054 41104 23060
rect 40960 23044 41012 23050
rect 40960 22986 41012 22992
rect 40868 21480 40920 21486
rect 40868 21422 40920 21428
rect 40684 20868 40736 20874
rect 40684 20810 40736 20816
rect 40512 20726 40632 20754
rect 40500 20324 40552 20330
rect 40500 20266 40552 20272
rect 40224 20256 40276 20262
rect 40224 20198 40276 20204
rect 40236 18834 40264 20198
rect 40512 19922 40540 20266
rect 40500 19916 40552 19922
rect 40500 19858 40552 19864
rect 40408 19780 40460 19786
rect 40408 19722 40460 19728
rect 40316 19712 40368 19718
rect 40316 19654 40368 19660
rect 40328 19446 40356 19654
rect 40316 19440 40368 19446
rect 40316 19382 40368 19388
rect 40224 18828 40276 18834
rect 40224 18770 40276 18776
rect 40132 18760 40184 18766
rect 40132 18702 40184 18708
rect 40144 18426 40172 18702
rect 40132 18420 40184 18426
rect 40132 18362 40184 18368
rect 40132 18284 40184 18290
rect 40132 18226 40184 18232
rect 40040 17808 40092 17814
rect 40040 17750 40092 17756
rect 39948 17196 40000 17202
rect 39948 17138 40000 17144
rect 39856 16108 39908 16114
rect 39856 16050 39908 16056
rect 39868 15706 39896 16050
rect 39856 15700 39908 15706
rect 39856 15642 39908 15648
rect 39960 15434 39988 17138
rect 40144 16998 40172 18226
rect 40132 16992 40184 16998
rect 40132 16934 40184 16940
rect 40040 16516 40092 16522
rect 40040 16458 40092 16464
rect 40052 16182 40080 16458
rect 40040 16176 40092 16182
rect 40040 16118 40092 16124
rect 39948 15428 40000 15434
rect 39948 15370 40000 15376
rect 39764 14068 39816 14074
rect 39764 14010 39816 14016
rect 39776 13870 39804 14010
rect 39764 13864 39816 13870
rect 39764 13806 39816 13812
rect 39960 13190 39988 15370
rect 40144 14618 40172 16934
rect 40224 16448 40276 16454
rect 40224 16390 40276 16396
rect 40236 15366 40264 16390
rect 40224 15360 40276 15366
rect 40224 15302 40276 15308
rect 40132 14612 40184 14618
rect 40132 14554 40184 14560
rect 39488 13184 39540 13190
rect 39488 13126 39540 13132
rect 39948 13184 40000 13190
rect 39948 13126 40000 13132
rect 39500 11830 39528 13126
rect 39488 11824 39540 11830
rect 39488 11766 39540 11772
rect 40420 11150 40448 19722
rect 40512 17338 40540 19858
rect 40604 19378 40632 20726
rect 40696 20448 40724 20810
rect 40972 20602 41000 22986
rect 40960 20596 41012 20602
rect 40960 20538 41012 20544
rect 40957 20460 41009 20466
rect 40696 20420 40957 20448
rect 40592 19372 40644 19378
rect 40592 19314 40644 19320
rect 40604 17882 40632 19314
rect 40696 18222 40724 20420
rect 40957 20402 41009 20408
rect 41064 20330 41092 23054
rect 41248 22506 41276 23802
rect 41432 23186 41460 24006
rect 41420 23180 41472 23186
rect 41420 23122 41472 23128
rect 41236 22500 41288 22506
rect 41236 22442 41288 22448
rect 41144 20800 41196 20806
rect 41196 20760 41276 20788
rect 41144 20742 41196 20748
rect 41248 20398 41276 20760
rect 41236 20392 41288 20398
rect 41236 20334 41288 20340
rect 41052 20324 41104 20330
rect 41052 20266 41104 20272
rect 40776 19848 40828 19854
rect 40776 19790 40828 19796
rect 40960 19848 41012 19854
rect 41064 19836 41092 20266
rect 41012 19808 41092 19836
rect 40960 19790 41012 19796
rect 40788 19514 40816 19790
rect 40776 19508 40828 19514
rect 40776 19450 40828 19456
rect 40776 18624 40828 18630
rect 40776 18566 40828 18572
rect 40788 18290 40816 18566
rect 40776 18284 40828 18290
rect 40776 18226 40828 18232
rect 40684 18216 40736 18222
rect 40684 18158 40736 18164
rect 40592 17876 40644 17882
rect 40592 17818 40644 17824
rect 40696 17746 40724 18158
rect 40684 17740 40736 17746
rect 40684 17682 40736 17688
rect 40500 17332 40552 17338
rect 40500 17274 40552 17280
rect 40972 16046 41000 19790
rect 41052 18352 41104 18358
rect 41052 18294 41104 18300
rect 41064 17814 41092 18294
rect 41052 17808 41104 17814
rect 41052 17750 41104 17756
rect 40684 16040 40736 16046
rect 40684 15982 40736 15988
rect 40960 16040 41012 16046
rect 40960 15982 41012 15988
rect 40696 14414 40724 15982
rect 40972 15502 41000 15982
rect 40960 15496 41012 15502
rect 40960 15438 41012 15444
rect 40684 14408 40736 14414
rect 40684 14350 40736 14356
rect 40696 14006 40724 14350
rect 40684 14000 40736 14006
rect 40684 13942 40736 13948
rect 40408 11144 40460 11150
rect 40408 11086 40460 11092
rect 40420 10810 40448 11086
rect 40408 10804 40460 10810
rect 40408 10746 40460 10752
rect 39396 10056 39448 10062
rect 39396 9998 39448 10004
rect 39408 9722 39436 9998
rect 39396 9716 39448 9722
rect 39396 9658 39448 9664
rect 39304 8492 39356 8498
rect 39304 8434 39356 8440
rect 38660 8424 38712 8430
rect 38660 8366 38712 8372
rect 39120 8424 39172 8430
rect 39120 8366 39172 8372
rect 38292 7404 38344 7410
rect 38292 7346 38344 7352
rect 37924 6316 37976 6322
rect 37924 6258 37976 6264
rect 37372 5568 37424 5574
rect 37372 5510 37424 5516
rect 36268 5364 36320 5370
rect 36268 5306 36320 5312
rect 37936 5302 37964 6258
rect 38304 5710 38332 7346
rect 38672 6866 38700 8366
rect 38844 7812 38896 7818
rect 38844 7754 38896 7760
rect 38856 7478 38884 7754
rect 38844 7472 38896 7478
rect 38844 7414 38896 7420
rect 38384 6860 38436 6866
rect 38384 6802 38436 6808
rect 38660 6860 38712 6866
rect 38660 6802 38712 6808
rect 38292 5704 38344 5710
rect 38292 5646 38344 5652
rect 37924 5296 37976 5302
rect 37924 5238 37976 5244
rect 38396 5234 38424 6802
rect 38568 6656 38620 6662
rect 38568 6598 38620 6604
rect 38580 6322 38608 6598
rect 38672 6390 38700 6802
rect 38856 6458 38884 7414
rect 38936 7200 38988 7206
rect 38936 7142 38988 7148
rect 38948 6798 38976 7142
rect 39316 6798 39344 8434
rect 38936 6792 38988 6798
rect 38936 6734 38988 6740
rect 39304 6792 39356 6798
rect 39304 6734 39356 6740
rect 39316 6662 39344 6734
rect 39304 6656 39356 6662
rect 39304 6598 39356 6604
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 38660 6384 38712 6390
rect 38660 6326 38712 6332
rect 38568 6316 38620 6322
rect 38568 6258 38620 6264
rect 38384 5228 38436 5234
rect 38384 5170 38436 5176
rect 35624 4004 35676 4010
rect 35624 3946 35676 3952
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 34520 3052 34572 3058
rect 34520 2994 34572 3000
rect 32772 2984 32824 2990
rect 32772 2926 32824 2932
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 29552 1896 29604 1902
rect 29552 1838 29604 1844
rect 29748 800 29776 2790
rect 30024 800 30052 2790
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30300 800 30328 2382
rect 30576 800 30604 2790
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 30852 800 30880 2382
rect 31128 800 31156 2382
rect 31404 800 31432 2382
rect 31680 800 31708 2790
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 31956 800 31984 2450
rect 32232 800 32260 2790
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32508 800 32536 2382
rect 32784 800 32812 2926
rect 33876 2916 33928 2922
rect 33876 2858 33928 2864
rect 33324 2848 33376 2854
rect 33324 2790 33376 2796
rect 33048 2508 33100 2514
rect 33048 2450 33100 2456
rect 33060 800 33088 2450
rect 33336 800 33364 2790
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33612 800 33640 2382
rect 33888 800 33916 2858
rect 34428 2848 34480 2854
rect 34428 2790 34480 2796
rect 34152 1420 34204 1426
rect 34152 1362 34204 1368
rect 34164 800 34192 1362
rect 34440 800 34468 2790
rect 34716 800 34744 3470
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 1850 35388 3470
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 34992 1822 35388 1850
rect 34992 800 35020 1822
rect 35452 1442 35480 2790
rect 35268 1414 35480 1442
rect 35544 2650 35664 2666
rect 35544 2644 35676 2650
rect 35544 2638 35624 2644
rect 35268 800 35296 1414
rect 35544 800 35572 2638
rect 35624 2586 35676 2592
rect 35624 2508 35676 2514
rect 35624 2450 35676 2456
rect 35636 2106 35664 2450
rect 35716 2440 35768 2446
rect 35716 2382 35768 2388
rect 35624 2100 35676 2106
rect 35624 2042 35676 2048
rect 35728 1426 35756 2382
rect 35716 1420 35768 1426
rect 35716 1362 35768 1368
rect 35820 800 35848 3470
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36096 800 36124 2382
rect 36372 800 36400 2790
rect 36544 2372 36596 2378
rect 36544 2314 36596 2320
rect 36556 2106 36584 2314
rect 36544 2100 36596 2106
rect 36544 2042 36596 2048
rect 36648 800 36676 3470
rect 37188 2916 37240 2922
rect 37188 2858 37240 2864
rect 36728 2576 36780 2582
rect 36728 2518 36780 2524
rect 36740 2378 36768 2518
rect 36912 2508 36964 2514
rect 36912 2450 36964 2456
rect 36728 2372 36780 2378
rect 36728 2314 36780 2320
rect 36924 800 36952 2450
rect 37200 800 37228 2858
rect 37476 800 37504 3470
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 37740 2848 37792 2854
rect 37740 2790 37792 2796
rect 37752 800 37780 2790
rect 38016 2576 38068 2582
rect 38016 2518 38068 2524
rect 38028 800 38056 2518
rect 38304 800 38332 2926
rect 38580 800 38608 3470
rect 39120 2916 39172 2922
rect 39120 2858 39172 2864
rect 38844 2508 38896 2514
rect 38844 2450 38896 2456
rect 38856 800 38884 2450
rect 39132 800 39160 2858
rect 39672 2848 39724 2854
rect 39672 2790 39724 2796
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39408 800 39436 2382
rect 39684 800 39712 2790
rect 39960 800 39988 3470
rect 40224 2916 40276 2922
rect 40224 2858 40276 2864
rect 40236 800 40264 2858
rect 40512 800 40540 3470
rect 40776 2508 40828 2514
rect 40776 2450 40828 2456
rect 40788 800 40816 2450
rect 41064 800 41092 3470
rect 42156 2984 42208 2990
rect 42156 2926 42208 2932
rect 41604 2848 41656 2854
rect 41604 2790 41656 2796
rect 41328 2440 41380 2446
rect 41328 2382 41380 2388
rect 41340 800 41368 2382
rect 41616 800 41644 2790
rect 41880 2576 41932 2582
rect 41880 2518 41932 2524
rect 41892 800 41920 2518
rect 42168 800 42196 2926
rect 42444 800 42472 3470
rect 42720 800 42748 3470
rect 42904 2650 42932 55558
rect 43168 51400 43220 51406
rect 43168 51342 43220 51348
rect 42984 2916 43036 2922
rect 42984 2858 43036 2864
rect 42892 2644 42944 2650
rect 42892 2586 42944 2592
rect 42996 800 43024 2858
rect 43180 2378 43208 51342
rect 43548 6914 43576 55558
rect 44008 55418 44036 55558
rect 43996 55412 44048 55418
rect 43996 55354 44048 55360
rect 43456 6886 43576 6914
rect 43260 2508 43312 2514
rect 43260 2450 43312 2456
rect 43168 2372 43220 2378
rect 43168 2314 43220 2320
rect 43272 800 43300 2450
rect 43456 2038 43484 6886
rect 44364 3528 44416 3534
rect 44364 3470 44416 3476
rect 44088 2916 44140 2922
rect 44088 2858 44140 2864
rect 43536 2848 43588 2854
rect 43536 2790 43588 2796
rect 43444 2032 43496 2038
rect 43444 1974 43496 1980
rect 43548 800 43576 2790
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 44100 800 44128 2858
rect 44376 800 44404 3470
rect 44640 2372 44692 2378
rect 44640 2314 44692 2320
rect 44652 800 44680 2314
rect 44744 2106 44772 55558
rect 45480 42265 45508 56306
rect 46124 55622 46152 56306
rect 46768 55622 46796 56306
rect 47688 56166 47716 57394
rect 48320 57384 48372 57390
rect 48320 57326 48372 57332
rect 48332 56234 48360 57326
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 53484 56438 53512 57394
rect 53472 56432 53524 56438
rect 53472 56374 53524 56380
rect 55324 56302 55352 57394
rect 56060 57254 56088 57394
rect 56048 57248 56100 57254
rect 56048 57190 56100 57196
rect 55312 56296 55364 56302
rect 55312 56238 55364 56244
rect 48320 56228 48372 56234
rect 48320 56170 48372 56176
rect 47676 56160 47728 56166
rect 47676 56102 47728 56108
rect 46112 55616 46164 55622
rect 46112 55558 46164 55564
rect 46756 55616 46808 55622
rect 46756 55558 46808 55564
rect 45466 42256 45522 42265
rect 45466 42191 45522 42200
rect 46124 42129 46152 55558
rect 46110 42120 46166 42129
rect 46110 42055 46166 42064
rect 46768 4826 46796 55558
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 56060 51270 56088 57190
rect 57532 57050 57560 57831
rect 58084 57594 58112 59200
rect 58438 59191 58494 59200
rect 58072 57588 58124 57594
rect 58072 57530 58124 57536
rect 57796 57452 57848 57458
rect 57796 57394 57848 57400
rect 57520 57044 57572 57050
rect 57520 56986 57572 56992
rect 56048 51264 56100 51270
rect 56048 51206 56100 51212
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 56324 45484 56376 45490
rect 56324 45426 56376 45432
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 53748 5160 53800 5166
rect 53748 5102 53800 5108
rect 53656 5024 53708 5030
rect 53656 4966 53708 4972
rect 46756 4820 46808 4826
rect 46756 4762 46808 4768
rect 52184 4752 52236 4758
rect 52184 4694 52236 4700
rect 52092 4616 52144 4622
rect 52092 4558 52144 4564
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 51816 4072 51868 4078
rect 51816 4014 51868 4020
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 51356 3936 51408 3942
rect 51356 3878 51408 3884
rect 46296 3664 46348 3670
rect 46296 3606 46348 3612
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44732 2100 44784 2106
rect 44732 2042 44784 2048
rect 44928 800 44956 2790
rect 45204 800 45232 3470
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 45480 800 45508 2790
rect 45744 2576 45796 2582
rect 45744 2518 45796 2524
rect 45756 800 45784 2518
rect 46032 800 46060 3470
rect 46308 800 46336 3606
rect 50804 3596 50856 3602
rect 50804 3538 50856 3544
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 47400 2916 47452 2922
rect 47400 2858 47452 2864
rect 46848 2848 46900 2854
rect 46848 2790 46900 2796
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 46584 800 46612 2450
rect 46860 800 46888 2790
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 47136 800 47164 2382
rect 47412 800 47440 2858
rect 47688 800 47716 3470
rect 47952 2848 48004 2854
rect 47952 2790 48004 2796
rect 47964 800 47992 2790
rect 48240 800 48268 3470
rect 48780 2916 48832 2922
rect 48780 2858 48832 2864
rect 49884 2916 49936 2922
rect 49884 2858 49936 2864
rect 48504 2508 48556 2514
rect 48504 2450 48556 2456
rect 48516 800 48544 2450
rect 48792 800 48820 2858
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 49068 800 49096 2382
rect 49344 800 49372 2790
rect 49608 2576 49660 2582
rect 49608 2518 49660 2524
rect 49620 800 49648 2518
rect 49896 800 49924 2858
rect 50172 800 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1850 50660 3470
rect 50712 2848 50764 2854
rect 50712 2790 50764 2796
rect 50448 1822 50660 1850
rect 50448 800 50476 1822
rect 50724 1442 50752 2790
rect 50632 1414 50752 1442
rect 50632 800 50660 1414
rect 50816 1306 50844 3538
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50896 2440 50948 2446
rect 50896 2382 50948 2388
rect 50724 1278 50844 1306
rect 50724 800 50752 1278
rect 50908 1170 50936 2382
rect 50816 1142 50936 1170
rect 50816 800 50844 1142
rect 51000 1034 51028 2858
rect 50908 1006 51028 1034
rect 50908 800 50936 1006
rect 50988 944 51040 950
rect 50988 886 51040 892
rect 51000 800 51028 886
rect 51092 800 51120 3878
rect 51172 3528 51224 3534
rect 51172 3470 51224 3476
rect 51184 800 51212 3470
rect 51264 2508 51316 2514
rect 51264 2450 51316 2456
rect 51276 800 51304 2450
rect 51368 800 51396 3878
rect 51448 3664 51500 3670
rect 51448 3606 51500 3612
rect 51460 800 51488 3606
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 51540 2848 51592 2854
rect 51540 2790 51592 2796
rect 51552 800 51580 2790
rect 51644 800 51672 3538
rect 51724 3052 51776 3058
rect 51724 2994 51776 3000
rect 51736 800 51764 2994
rect 51828 800 51856 4014
rect 51908 3120 51960 3126
rect 51908 3062 51960 3068
rect 51920 800 51948 3062
rect 52000 2644 52052 2650
rect 52000 2586 52052 2592
rect 52012 800 52040 2586
rect 52104 800 52132 4558
rect 52196 800 52224 4694
rect 53196 4684 53248 4690
rect 53196 4626 53248 4632
rect 52644 4616 52696 4622
rect 52644 4558 52696 4564
rect 52460 3936 52512 3942
rect 52460 3878 52512 3884
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 52288 800 52316 3470
rect 52368 2372 52420 2378
rect 52368 2314 52420 2320
rect 52380 800 52408 2314
rect 52472 800 52500 3878
rect 52552 2508 52604 2514
rect 52552 2450 52604 2456
rect 52564 1154 52592 2450
rect 52552 1148 52604 1154
rect 52552 1090 52604 1096
rect 52552 1012 52604 1018
rect 52552 954 52604 960
rect 52564 800 52592 954
rect 52656 800 52684 4558
rect 53012 4140 53064 4146
rect 53012 4082 53064 4088
rect 52828 4004 52880 4010
rect 52828 3946 52880 3952
rect 52736 3732 52788 3738
rect 52736 3674 52788 3680
rect 52748 2106 52776 3674
rect 52736 2100 52788 2106
rect 52736 2042 52788 2048
rect 52840 1986 52868 3946
rect 52920 2100 52972 2106
rect 52920 2042 52972 2048
rect 52748 1958 52868 1986
rect 52748 800 52776 1958
rect 52828 1488 52880 1494
rect 52828 1430 52880 1436
rect 52840 800 52868 1430
rect 52932 800 52960 2042
rect 53024 1494 53052 4082
rect 53104 2984 53156 2990
rect 53104 2926 53156 2932
rect 53012 1488 53064 1494
rect 53012 1430 53064 1436
rect 53012 1352 53064 1358
rect 53012 1294 53064 1300
rect 53024 800 53052 1294
rect 53116 800 53144 2926
rect 53208 800 53236 4626
rect 53288 3460 53340 3466
rect 53288 3402 53340 3408
rect 53300 800 53328 3402
rect 53378 2952 53434 2961
rect 53378 2887 53434 2896
rect 53392 800 53420 2887
rect 53470 2816 53526 2825
rect 53470 2751 53526 2760
rect 53484 800 53512 2751
rect 53564 2508 53616 2514
rect 53564 2450 53616 2456
rect 53576 800 53604 2450
rect 53668 800 53696 4966
rect 53760 800 53788 5102
rect 54116 5092 54168 5098
rect 54116 5034 54168 5040
rect 53932 4752 53984 4758
rect 53932 4694 53984 4700
rect 53840 3596 53892 3602
rect 53840 3538 53892 3544
rect 53852 800 53880 3538
rect 53944 800 53972 4694
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 54036 800 54064 4014
rect 54128 800 54156 5034
rect 54300 4684 54352 4690
rect 54300 4626 54352 4632
rect 54208 2916 54260 2922
rect 54208 2858 54260 2864
rect 54220 800 54248 2858
rect 54312 800 54340 4626
rect 55312 3936 55364 3942
rect 55312 3878 55364 3884
rect 54760 3052 54812 3058
rect 54760 2994 54812 3000
rect 54392 2576 54444 2582
rect 54392 2518 54444 2524
rect 54404 2106 54432 2518
rect 54392 2100 54444 2106
rect 54392 2042 54444 2048
rect 54772 1018 54800 2994
rect 55324 2825 55352 3878
rect 55310 2816 55366 2825
rect 55310 2751 55366 2760
rect 56336 2310 56364 45426
rect 57808 45354 57836 57394
rect 57888 56840 57940 56846
rect 57888 56782 57940 56788
rect 57900 56545 57928 56782
rect 57886 56536 57942 56545
rect 57886 56471 57942 56480
rect 58452 56370 58480 59191
rect 58440 56364 58492 56370
rect 58440 56306 58492 56312
rect 58162 55176 58218 55185
rect 58162 55111 58164 55120
rect 58216 55111 58218 55120
rect 58164 55082 58216 55088
rect 57888 53984 57940 53990
rect 57888 53926 57940 53932
rect 57900 53825 57928 53926
rect 57886 53816 57942 53825
rect 57886 53751 57942 53760
rect 57888 52488 57940 52494
rect 57886 52456 57888 52465
rect 57940 52456 57942 52465
rect 57886 52391 57942 52400
rect 58164 51400 58216 51406
rect 58164 51342 58216 51348
rect 58176 51105 58204 51342
rect 58162 51096 58218 51105
rect 58162 51031 58218 51040
rect 58164 49768 58216 49774
rect 58162 49736 58164 49745
rect 58216 49736 58218 49745
rect 58162 49671 58218 49680
rect 58164 48544 58216 48550
rect 58164 48486 58216 48492
rect 58176 48385 58204 48486
rect 58162 48376 58218 48385
rect 58162 48311 58218 48320
rect 58164 47048 58216 47054
rect 58162 47016 58164 47025
rect 58216 47016 58218 47025
rect 58162 46951 58218 46960
rect 58164 45960 58216 45966
rect 58164 45902 58216 45908
rect 58176 45665 58204 45902
rect 58162 45656 58218 45665
rect 58162 45591 58218 45600
rect 57796 45348 57848 45354
rect 57796 45290 57848 45296
rect 58162 44296 58218 44305
rect 58162 44231 58164 44240
rect 58216 44231 58218 44240
rect 58164 44202 58216 44208
rect 58164 43104 58216 43110
rect 58164 43046 58216 43052
rect 58176 42945 58204 43046
rect 58162 42936 58218 42945
rect 58162 42871 58218 42880
rect 58164 41608 58216 41614
rect 58162 41576 58164 41585
rect 58216 41576 58218 41585
rect 58162 41511 58218 41520
rect 58164 40520 58216 40526
rect 58164 40462 58216 40468
rect 58176 40225 58204 40462
rect 58162 40216 58218 40225
rect 58162 40151 58218 40160
rect 58162 38856 58218 38865
rect 58162 38791 58164 38800
rect 58216 38791 58218 38800
rect 58164 38762 58216 38768
rect 58164 37664 58216 37670
rect 58164 37606 58216 37612
rect 58176 37505 58204 37606
rect 58162 37496 58218 37505
rect 58162 37431 58218 37440
rect 58164 36168 58216 36174
rect 58162 36136 58164 36145
rect 58216 36136 58218 36145
rect 58162 36071 58218 36080
rect 58164 35080 58216 35086
rect 58164 35022 58216 35028
rect 58176 34785 58204 35022
rect 58162 34776 58218 34785
rect 58162 34711 58218 34720
rect 58162 33416 58218 33425
rect 58162 33351 58164 33360
rect 58216 33351 58218 33360
rect 58164 33322 58216 33328
rect 58164 32224 58216 32230
rect 58164 32166 58216 32172
rect 58176 32065 58204 32166
rect 58162 32056 58218 32065
rect 58162 31991 58218 32000
rect 58164 30728 58216 30734
rect 58162 30696 58164 30705
rect 58216 30696 58218 30705
rect 58162 30631 58218 30640
rect 58164 29640 58216 29646
rect 58164 29582 58216 29588
rect 58176 29345 58204 29582
rect 58162 29336 58218 29345
rect 58162 29271 58218 29280
rect 58162 27976 58218 27985
rect 58162 27911 58164 27920
rect 58216 27911 58218 27920
rect 58164 27882 58216 27888
rect 58164 26784 58216 26790
rect 58164 26726 58216 26732
rect 58176 26625 58204 26726
rect 58162 26616 58218 26625
rect 58162 26551 58218 26560
rect 58164 25288 58216 25294
rect 58162 25256 58164 25265
rect 58216 25256 58218 25265
rect 58162 25191 58218 25200
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 58176 23905 58204 24142
rect 58162 23896 58218 23905
rect 58162 23831 58218 23840
rect 58162 22536 58218 22545
rect 58162 22471 58164 22480
rect 58216 22471 58218 22480
rect 58164 22442 58216 22448
rect 58164 21344 58216 21350
rect 58164 21286 58216 21292
rect 58176 21185 58204 21286
rect 58162 21176 58218 21185
rect 58162 21111 58218 21120
rect 58164 19848 58216 19854
rect 58162 19816 58164 19825
rect 58216 19816 58218 19825
rect 58162 19751 58218 19760
rect 58164 18760 58216 18766
rect 58164 18702 58216 18708
rect 58176 18465 58204 18702
rect 58162 18456 58218 18465
rect 58162 18391 58218 18400
rect 58162 17096 58218 17105
rect 58162 17031 58164 17040
rect 58216 17031 58218 17040
rect 58164 17002 58216 17008
rect 58164 15904 58216 15910
rect 58164 15846 58216 15852
rect 58176 15745 58204 15846
rect 58162 15736 58218 15745
rect 58162 15671 58218 15680
rect 58164 14408 58216 14414
rect 58162 14376 58164 14385
rect 58216 14376 58218 14385
rect 58162 14311 58218 14320
rect 58164 13320 58216 13326
rect 58164 13262 58216 13268
rect 58176 13025 58204 13262
rect 58162 13016 58218 13025
rect 58162 12951 58218 12960
rect 58162 11656 58218 11665
rect 58162 11591 58164 11600
rect 58216 11591 58218 11600
rect 58164 11562 58216 11568
rect 58164 10464 58216 10470
rect 58164 10406 58216 10412
rect 58176 10305 58204 10406
rect 58162 10296 58218 10305
rect 58162 10231 58218 10240
rect 58164 8968 58216 8974
rect 58162 8936 58164 8945
rect 58216 8936 58218 8945
rect 58162 8871 58218 8880
rect 58164 7880 58216 7886
rect 58164 7822 58216 7828
rect 58176 7585 58204 7822
rect 58162 7576 58218 7585
rect 58162 7511 58218 7520
rect 58162 6216 58218 6225
rect 58162 6151 58164 6160
rect 58216 6151 58218 6160
rect 58164 6122 58216 6128
rect 58164 5024 58216 5030
rect 58164 4966 58216 4972
rect 58176 4865 58204 4966
rect 58162 4856 58218 4865
rect 58162 4791 58218 4800
rect 58440 3936 58492 3942
rect 58440 3878 58492 3884
rect 57520 3528 57572 3534
rect 58164 3528 58216 3534
rect 57520 3470 57572 3476
rect 58162 3496 58164 3505
rect 58216 3496 58218 3505
rect 56600 2984 56652 2990
rect 56598 2952 56600 2961
rect 56652 2952 56654 2961
rect 56598 2887 56654 2896
rect 56324 2304 56376 2310
rect 56324 2246 56376 2252
rect 57532 2145 57560 3470
rect 58162 3431 58218 3440
rect 57518 2136 57574 2145
rect 57518 2071 57574 2080
rect 54760 1012 54812 1018
rect 54760 954 54812 960
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 58452 785 58480 3878
rect 58438 776 58494 785
rect 58438 711 58494 720
<< via2 >>
rect 58438 59200 58494 59256
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 57518 57840 57574 57896
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 14186 55564 14188 55584
rect 14188 55564 14240 55584
rect 14240 55564 14242 55584
rect 14186 55528 14242 55564
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 11518 41692 11520 41712
rect 11520 41692 11572 41712
rect 11572 41692 11574 41712
rect 11518 41656 11574 41692
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4710 38936 4766 38992
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 2686 23060 2688 23080
rect 2688 23060 2740 23080
rect 2740 23060 2742 23080
rect 2686 23024 2742 23060
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 5538 33940 5540 33960
rect 5540 33940 5592 33960
rect 5592 33940 5594 33960
rect 5538 33904 5594 33940
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 5814 33904 5870 33960
rect 3054 23024 3110 23080
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1582 7928 1638 7984
rect 2778 8780 2780 8800
rect 2780 8780 2832 8800
rect 2832 8780 2834 8800
rect 2778 8744 2834 8780
rect 2134 3440 2190 3496
rect 2226 2896 2282 2952
rect 2778 5228 2834 5264
rect 2778 5208 2780 5228
rect 2780 5208 2832 5228
rect 2832 5208 2834 5228
rect 2962 2624 3018 2680
rect 3146 3984 3202 4040
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 6734 38956 6790 38992
rect 6734 38936 6736 38956
rect 6736 38936 6788 38956
rect 6788 38936 6790 38956
rect 4802 15308 4804 15328
rect 4804 15308 4856 15328
rect 4856 15308 4858 15328
rect 4802 15272 4858 15308
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3330 3340 3332 3360
rect 3332 3340 3384 3360
rect 3384 3340 3386 3360
rect 3330 3304 3386 3340
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4342 4684 4398 4720
rect 4342 4664 4344 4684
rect 4344 4664 4396 4684
rect 4396 4664 4398 4684
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 3974 3576 4030 3632
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1582 2216 1638 2272
rect 4250 2352 4306 2408
rect 4894 4256 4950 4312
rect 5630 7284 5632 7304
rect 5632 7284 5684 7304
rect 5684 7284 5686 7304
rect 5630 7248 5686 7284
rect 5262 4428 5264 4448
rect 5264 4428 5316 4448
rect 5316 4428 5318 4448
rect 5262 4392 5318 4428
rect 5262 4256 5318 4312
rect 5538 2352 5594 2408
rect 5814 2488 5870 2544
rect 6182 3596 6238 3632
rect 6182 3576 6184 3596
rect 6184 3576 6236 3596
rect 6236 3576 6238 3596
rect 7102 10784 7158 10840
rect 6826 8336 6882 8392
rect 8574 29180 8576 29200
rect 8576 29180 8628 29200
rect 8628 29180 8630 29200
rect 8574 29144 8630 29180
rect 8298 18828 8354 18864
rect 8298 18808 8300 18828
rect 8300 18808 8352 18828
rect 8352 18808 8354 18828
rect 8114 13776 8170 13832
rect 6458 3984 6514 4040
rect 7102 3984 7158 4040
rect 6826 3188 6882 3224
rect 6826 3168 6828 3188
rect 6828 3168 6880 3188
rect 6880 3168 6882 3188
rect 6918 2896 6974 2952
rect 7286 2896 7342 2952
rect 7654 2760 7710 2816
rect 7562 2624 7618 2680
rect 8390 7248 8446 7304
rect 7930 2896 7986 2952
rect 9586 29164 9642 29200
rect 9586 29144 9588 29164
rect 9588 29144 9640 29164
rect 9640 29144 9642 29164
rect 12898 41676 12954 41712
rect 12898 41656 12900 41676
rect 12900 41656 12952 41676
rect 12952 41656 12954 41676
rect 9862 19780 9918 19816
rect 9862 19760 9864 19780
rect 9864 19760 9916 19780
rect 9916 19760 9918 19780
rect 10046 15564 10102 15600
rect 10046 15544 10048 15564
rect 10048 15544 10100 15564
rect 10100 15544 10102 15564
rect 9678 11056 9734 11112
rect 9402 10376 9458 10432
rect 9402 9968 9458 10024
rect 8850 4392 8906 4448
rect 9586 8064 9642 8120
rect 9402 3984 9458 4040
rect 8482 2216 8538 2272
rect 9310 3848 9366 3904
rect 9218 3476 9220 3496
rect 9220 3476 9272 3496
rect 9272 3476 9274 3496
rect 9218 3440 9274 3476
rect 9218 2216 9274 2272
rect 9586 5208 9642 5264
rect 9678 3984 9734 4040
rect 9770 3732 9826 3768
rect 9770 3712 9772 3732
rect 9772 3712 9824 3732
rect 9824 3712 9826 3732
rect 12622 34584 12678 34640
rect 13174 33088 13230 33144
rect 10506 15408 10562 15464
rect 10782 15444 10784 15464
rect 10784 15444 10836 15464
rect 10836 15444 10838 15464
rect 10782 15408 10838 15444
rect 10598 10512 10654 10568
rect 12898 24148 12900 24168
rect 12900 24148 12952 24168
rect 12952 24148 12954 24168
rect 12898 24112 12954 24148
rect 14462 33532 14464 33552
rect 14464 33532 14516 33552
rect 14516 33532 14518 33552
rect 14462 33496 14518 33532
rect 14830 24148 14832 24168
rect 14832 24148 14884 24168
rect 14884 24148 14886 24168
rect 14830 24112 14886 24148
rect 12254 13232 12310 13288
rect 10414 2352 10470 2408
rect 10690 3304 10746 3360
rect 11886 7540 11942 7576
rect 11886 7520 11888 7540
rect 11888 7520 11940 7540
rect 11940 7520 11942 7540
rect 12990 15408 13046 15464
rect 12806 6296 12862 6352
rect 13542 6296 13598 6352
rect 13726 3068 13728 3088
rect 13728 3068 13780 3088
rect 13780 3068 13782 3088
rect 13726 3032 13782 3068
rect 14462 3984 14518 4040
rect 14554 2624 14610 2680
rect 14922 3168 14978 3224
rect 15198 19916 15254 19952
rect 15198 19896 15200 19916
rect 15200 19896 15252 19916
rect 15252 19896 15254 19916
rect 15474 3032 15530 3088
rect 16026 8236 16028 8256
rect 16028 8236 16080 8256
rect 16080 8236 16082 8256
rect 16026 8200 16082 8236
rect 16026 2352 16082 2408
rect 16578 55564 16580 55584
rect 16580 55564 16632 55584
rect 16632 55564 16634 55584
rect 16578 55528 16634 55564
rect 17222 55564 17224 55584
rect 17224 55564 17276 55584
rect 17276 55564 17278 55584
rect 17222 55528 17278 55564
rect 17406 33532 17408 33552
rect 17408 33532 17460 33552
rect 17460 33532 17462 33552
rect 17406 33496 17462 33532
rect 17222 23568 17278 23624
rect 16302 2624 16358 2680
rect 16762 8508 16764 8528
rect 16764 8508 16816 8528
rect 16816 8508 16818 8528
rect 16762 8472 16818 8508
rect 17682 8084 17738 8120
rect 17682 8064 17684 8084
rect 17684 8064 17736 8084
rect 17736 8064 17738 8084
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 18510 23604 18512 23624
rect 18512 23604 18564 23624
rect 18564 23604 18566 23624
rect 18510 23568 18566 23604
rect 18970 34620 18972 34640
rect 18972 34620 19024 34640
rect 19024 34620 19026 34640
rect 18970 34584 19026 34620
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 20350 56108 20352 56128
rect 20352 56108 20404 56128
rect 20404 56108 20406 56128
rect 20350 56072 20406 56108
rect 23110 56208 23166 56264
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19430 34584 19486 34640
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 17958 8492 18014 8528
rect 17958 8472 17960 8492
rect 17960 8472 18012 8492
rect 18012 8472 18014 8492
rect 17682 2644 17738 2680
rect 17682 2624 17684 2644
rect 17684 2624 17736 2644
rect 17736 2624 17738 2644
rect 18234 3188 18290 3224
rect 18234 3168 18236 3188
rect 18236 3168 18288 3188
rect 18288 3168 18290 3188
rect 18510 2524 18512 2544
rect 18512 2524 18564 2544
rect 18564 2524 18566 2544
rect 18510 2488 18566 2524
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19430 20576 19486 20632
rect 19430 20440 19486 20496
rect 19798 20304 19854 20360
rect 20166 20712 20222 20768
rect 20442 23044 20498 23080
rect 20442 23024 20444 23044
rect 20444 23024 20496 23044
rect 20496 23024 20498 23044
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20534 20476 20536 20496
rect 20536 20476 20588 20496
rect 20588 20476 20590 20496
rect 20534 20440 20590 20476
rect 21730 26324 21732 26344
rect 21732 26324 21784 26344
rect 21784 26324 21786 26344
rect 21730 26288 21786 26324
rect 21638 23704 21694 23760
rect 21822 20712 21878 20768
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 18878 3188 18934 3224
rect 18878 3168 18880 3188
rect 18880 3168 18932 3188
rect 18932 3168 18934 3188
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20442 5616 20498 5672
rect 20350 3984 20406 4040
rect 22466 26288 22522 26344
rect 22650 23740 22652 23760
rect 22652 23740 22704 23760
rect 22704 23740 22706 23760
rect 22650 23704 22706 23740
rect 22926 13232 22982 13288
rect 22742 12144 22798 12200
rect 21086 3188 21142 3224
rect 21086 3168 21088 3188
rect 21088 3168 21140 3188
rect 21140 3168 21142 3188
rect 21914 3732 21970 3768
rect 21914 3712 21916 3732
rect 21916 3712 21968 3732
rect 21968 3712 21970 3732
rect 27618 55700 27620 55720
rect 27620 55700 27672 55720
rect 27672 55700 27674 55720
rect 27618 55664 27674 55700
rect 23754 29144 23810 29200
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 30010 43696 30066 43752
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 33598 44784 33654 44840
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 32126 42336 32182 42392
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 24398 29144 24454 29200
rect 24030 15544 24086 15600
rect 23938 13776 23994 13832
rect 25502 29688 25558 29744
rect 26146 29028 26202 29064
rect 26146 29008 26148 29028
rect 26148 29008 26200 29028
rect 26200 29008 26202 29028
rect 26698 33940 26700 33960
rect 26700 33940 26752 33960
rect 26752 33940 26754 33960
rect 26698 33904 26754 33940
rect 27526 29008 27582 29064
rect 25594 19624 25650 19680
rect 25962 17176 26018 17232
rect 25502 12180 25504 12200
rect 25504 12180 25556 12200
rect 25556 12180 25558 12200
rect 25502 12144 25558 12180
rect 26974 19896 27030 19952
rect 26974 6316 27030 6352
rect 26974 6296 26976 6316
rect 26976 6296 27028 6316
rect 27028 6296 27030 6316
rect 26422 5244 26424 5264
rect 26424 5244 26476 5264
rect 26476 5244 26478 5264
rect 26422 5208 26478 5244
rect 28906 19624 28962 19680
rect 28538 10512 28594 10568
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 30654 37304 30710 37360
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 30838 21956 30894 21992
rect 30838 21936 30840 21956
rect 30840 21936 30892 21956
rect 30892 21936 30894 21956
rect 31482 29688 31538 29744
rect 30654 18844 30656 18864
rect 30656 18844 30708 18864
rect 30708 18844 30710 18864
rect 30654 18808 30710 18844
rect 30930 19760 30986 19816
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 31758 22500 31814 22536
rect 31758 22480 31760 22500
rect 31760 22480 31812 22500
rect 31812 22480 31814 22500
rect 32770 21972 32772 21992
rect 32772 21972 32824 21992
rect 32824 21972 32826 21992
rect 32770 21936 32826 21972
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34334 22500 34390 22536
rect 34334 22480 34336 22500
rect 34336 22480 34388 22500
rect 34388 22480 34390 22500
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 37278 15972 37334 16008
rect 37278 15952 37280 15972
rect 37280 15952 37332 15972
rect 37332 15952 37334 15972
rect 37278 8492 37334 8528
rect 37278 8472 37280 8492
rect 37280 8472 37332 8492
rect 37332 8472 37334 8492
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38842 8492 38898 8528
rect 38842 8472 38844 8492
rect 38844 8472 38896 8492
rect 38896 8472 38898 8492
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 45466 42200 45522 42256
rect 46110 42064 46166 42120
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 53378 2896 53434 2952
rect 53470 2760 53526 2816
rect 55310 2760 55366 2816
rect 57886 56480 57942 56536
rect 58162 55140 58218 55176
rect 58162 55120 58164 55140
rect 58164 55120 58216 55140
rect 58216 55120 58218 55140
rect 57886 53760 57942 53816
rect 57886 52436 57888 52456
rect 57888 52436 57940 52456
rect 57940 52436 57942 52456
rect 57886 52400 57942 52436
rect 58162 51040 58218 51096
rect 58162 49716 58164 49736
rect 58164 49716 58216 49736
rect 58216 49716 58218 49736
rect 58162 49680 58218 49716
rect 58162 48320 58218 48376
rect 58162 46996 58164 47016
rect 58164 46996 58216 47016
rect 58216 46996 58218 47016
rect 58162 46960 58218 46996
rect 58162 45600 58218 45656
rect 58162 44260 58218 44296
rect 58162 44240 58164 44260
rect 58164 44240 58216 44260
rect 58216 44240 58218 44260
rect 58162 42880 58218 42936
rect 58162 41556 58164 41576
rect 58164 41556 58216 41576
rect 58216 41556 58218 41576
rect 58162 41520 58218 41556
rect 58162 40160 58218 40216
rect 58162 38820 58218 38856
rect 58162 38800 58164 38820
rect 58164 38800 58216 38820
rect 58216 38800 58218 38820
rect 58162 37440 58218 37496
rect 58162 36116 58164 36136
rect 58164 36116 58216 36136
rect 58216 36116 58218 36136
rect 58162 36080 58218 36116
rect 58162 34720 58218 34776
rect 58162 33380 58218 33416
rect 58162 33360 58164 33380
rect 58164 33360 58216 33380
rect 58216 33360 58218 33380
rect 58162 32000 58218 32056
rect 58162 30676 58164 30696
rect 58164 30676 58216 30696
rect 58216 30676 58218 30696
rect 58162 30640 58218 30676
rect 58162 29280 58218 29336
rect 58162 27940 58218 27976
rect 58162 27920 58164 27940
rect 58164 27920 58216 27940
rect 58216 27920 58218 27940
rect 58162 26560 58218 26616
rect 58162 25236 58164 25256
rect 58164 25236 58216 25256
rect 58216 25236 58218 25256
rect 58162 25200 58218 25236
rect 58162 23840 58218 23896
rect 58162 22500 58218 22536
rect 58162 22480 58164 22500
rect 58164 22480 58216 22500
rect 58216 22480 58218 22500
rect 58162 21120 58218 21176
rect 58162 19796 58164 19816
rect 58164 19796 58216 19816
rect 58216 19796 58218 19816
rect 58162 19760 58218 19796
rect 58162 18400 58218 18456
rect 58162 17060 58218 17096
rect 58162 17040 58164 17060
rect 58164 17040 58216 17060
rect 58216 17040 58218 17060
rect 58162 15680 58218 15736
rect 58162 14356 58164 14376
rect 58164 14356 58216 14376
rect 58216 14356 58218 14376
rect 58162 14320 58218 14356
rect 58162 12960 58218 13016
rect 58162 11620 58218 11656
rect 58162 11600 58164 11620
rect 58164 11600 58216 11620
rect 58216 11600 58218 11620
rect 58162 10240 58218 10296
rect 58162 8916 58164 8936
rect 58164 8916 58216 8936
rect 58216 8916 58218 8936
rect 58162 8880 58218 8916
rect 58162 7520 58218 7576
rect 58162 6180 58218 6216
rect 58162 6160 58164 6180
rect 58164 6160 58216 6180
rect 58216 6160 58218 6180
rect 58162 4800 58218 4856
rect 58162 3476 58164 3496
rect 58164 3476 58216 3496
rect 58216 3476 58218 3496
rect 56598 2932 56600 2952
rect 56600 2932 56652 2952
rect 56652 2932 56654 2952
rect 56598 2896 56654 2932
rect 58162 3440 58218 3476
rect 57518 2080 57574 2136
rect 58438 720 58494 776
<< metal3 >>
rect 58433 59258 58499 59261
rect 59200 59258 60000 59288
rect 58433 59256 60000 59258
rect 58433 59200 58438 59256
rect 58494 59200 60000 59256
rect 58433 59198 60000 59200
rect 58433 59195 58499 59198
rect 59200 59168 60000 59198
rect 57513 57898 57579 57901
rect 59200 57898 60000 57928
rect 57513 57896 60000 57898
rect 57513 57840 57518 57896
rect 57574 57840 60000 57896
rect 57513 57838 60000 57840
rect 57513 57835 57579 57838
rect 59200 57808 60000 57838
rect 19570 57696 19886 57697
rect 0 57536 800 57656
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 57881 56538 57947 56541
rect 59200 56538 60000 56568
rect 57881 56536 60000 56538
rect 57881 56480 57886 56536
rect 57942 56480 60000 56536
rect 57881 56478 60000 56480
rect 57881 56475 57947 56478
rect 59200 56448 60000 56478
rect 23105 56266 23171 56269
rect 23238 56266 23244 56268
rect 23105 56264 23244 56266
rect 23105 56208 23110 56264
rect 23166 56208 23244 56264
rect 23105 56206 23244 56208
rect 23105 56203 23171 56206
rect 23238 56204 23244 56206
rect 23308 56204 23314 56268
rect 0 56040 800 56160
rect 20345 56130 20411 56133
rect 20478 56130 20484 56132
rect 20345 56128 20484 56130
rect 20345 56072 20350 56128
rect 20406 56072 20484 56128
rect 20345 56070 20484 56072
rect 20345 56067 20411 56070
rect 20478 56068 20484 56070
rect 20548 56068 20554 56132
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 23974 55660 23980 55724
rect 24044 55722 24050 55724
rect 27613 55722 27679 55725
rect 24044 55720 27679 55722
rect 24044 55664 27618 55720
rect 27674 55664 27679 55720
rect 24044 55662 27679 55664
rect 24044 55660 24050 55662
rect 27613 55659 27679 55662
rect 14181 55586 14247 55589
rect 14590 55586 14596 55588
rect 14181 55584 14596 55586
rect 14181 55528 14186 55584
rect 14242 55528 14596 55584
rect 14181 55526 14596 55528
rect 14181 55523 14247 55526
rect 14590 55524 14596 55526
rect 14660 55524 14666 55588
rect 15694 55524 15700 55588
rect 15764 55586 15770 55588
rect 16573 55586 16639 55589
rect 17217 55588 17283 55589
rect 15764 55584 16639 55586
rect 15764 55528 16578 55584
rect 16634 55528 16639 55584
rect 15764 55526 16639 55528
rect 15764 55524 15770 55526
rect 16573 55523 16639 55526
rect 17166 55524 17172 55588
rect 17236 55586 17283 55588
rect 17236 55584 17328 55586
rect 17278 55528 17328 55584
rect 17236 55526 17328 55528
rect 17236 55524 17283 55526
rect 17217 55523 17283 55524
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 58157 55178 58223 55181
rect 59200 55178 60000 55208
rect 58157 55176 60000 55178
rect 58157 55120 58162 55176
rect 58218 55120 60000 55176
rect 58157 55118 60000 55120
rect 58157 55115 58223 55118
rect 59200 55088 60000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 0 54544 800 54664
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 57881 53818 57947 53821
rect 59200 53818 60000 53848
rect 57881 53816 60000 53818
rect 57881 53760 57886 53816
rect 57942 53760 60000 53816
rect 57881 53758 60000 53760
rect 57881 53755 57947 53758
rect 59200 53728 60000 53758
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 0 53048 800 53168
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 57881 52458 57947 52461
rect 59200 52458 60000 52488
rect 57881 52456 60000 52458
rect 57881 52400 57886 52456
rect 57942 52400 60000 52456
rect 57881 52398 60000 52400
rect 57881 52395 57947 52398
rect 59200 52368 60000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51552 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 58157 51098 58223 51101
rect 59200 51098 60000 51128
rect 58157 51096 60000 51098
rect 58157 51040 58162 51096
rect 58218 51040 60000 51096
rect 58157 51038 60000 51040
rect 58157 51035 58223 51038
rect 59200 51008 60000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 0 50056 800 50176
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 58157 49738 58223 49741
rect 59200 49738 60000 49768
rect 58157 49736 60000 49738
rect 58157 49680 58162 49736
rect 58218 49680 60000 49736
rect 58157 49678 60000 49680
rect 58157 49675 58223 49678
rect 59200 49648 60000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48560 800 48680
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58157 48378 58223 48381
rect 59200 48378 60000 48408
rect 58157 48376 60000 48378
rect 58157 48320 58162 48376
rect 58218 48320 60000 48376
rect 58157 48318 60000 48320
rect 58157 48315 58223 48318
rect 59200 48288 60000 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 0 47064 800 47184
rect 58157 47018 58223 47021
rect 59200 47018 60000 47048
rect 58157 47016 60000 47018
rect 58157 46960 58162 47016
rect 58218 46960 60000 47016
rect 58157 46958 60000 46960
rect 58157 46955 58223 46958
rect 59200 46928 60000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 0 45568 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 58157 45658 58223 45661
rect 59200 45658 60000 45688
rect 58157 45656 60000 45658
rect 58157 45600 58162 45656
rect 58218 45600 60000 45656
rect 58157 45598 60000 45600
rect 58157 45595 58223 45598
rect 59200 45568 60000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 19006 44780 19012 44844
rect 19076 44842 19082 44844
rect 33593 44842 33659 44845
rect 19076 44840 33659 44842
rect 19076 44784 33598 44840
rect 33654 44784 33659 44840
rect 19076 44782 33659 44784
rect 19076 44780 19082 44782
rect 33593 44779 33659 44782
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 58157 44298 58223 44301
rect 59200 44298 60000 44328
rect 58157 44296 60000 44298
rect 58157 44240 58162 44296
rect 58218 44240 60000 44296
rect 58157 44238 60000 44240
rect 58157 44235 58223 44238
rect 59200 44208 60000 44238
rect 0 44072 800 44192
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 18270 43692 18276 43756
rect 18340 43754 18346 43756
rect 30005 43754 30071 43757
rect 18340 43752 30071 43754
rect 18340 43696 30010 43752
rect 30066 43696 30071 43752
rect 18340 43694 30071 43696
rect 18340 43692 18346 43694
rect 30005 43691 30071 43694
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 58157 42938 58223 42941
rect 59200 42938 60000 42968
rect 58157 42936 60000 42938
rect 58157 42880 58162 42936
rect 58218 42880 60000 42936
rect 58157 42878 60000 42880
rect 58157 42875 58223 42878
rect 59200 42848 60000 42878
rect 0 42576 800 42696
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 20110 42332 20116 42396
rect 20180 42394 20186 42396
rect 32121 42394 32187 42397
rect 20180 42392 32187 42394
rect 20180 42336 32126 42392
rect 32182 42336 32187 42392
rect 20180 42334 32187 42336
rect 20180 42332 20186 42334
rect 32121 42331 32187 42334
rect 21950 42196 21956 42260
rect 22020 42258 22026 42260
rect 45461 42258 45527 42261
rect 22020 42256 45527 42258
rect 22020 42200 45466 42256
rect 45522 42200 45527 42256
rect 22020 42198 45527 42200
rect 22020 42196 22026 42198
rect 45461 42195 45527 42198
rect 21214 42060 21220 42124
rect 21284 42122 21290 42124
rect 46105 42122 46171 42125
rect 21284 42120 46171 42122
rect 21284 42064 46110 42120
rect 46166 42064 46171 42120
rect 21284 42062 46171 42064
rect 21284 42060 21290 42062
rect 46105 42059 46171 42062
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 11513 41714 11579 41717
rect 12893 41714 12959 41717
rect 11513 41712 12959 41714
rect 11513 41656 11518 41712
rect 11574 41656 12898 41712
rect 12954 41656 12959 41712
rect 11513 41654 12959 41656
rect 11513 41651 11579 41654
rect 12893 41651 12959 41654
rect 58157 41578 58223 41581
rect 59200 41578 60000 41608
rect 58157 41576 60000 41578
rect 58157 41520 58162 41576
rect 58218 41520 60000 41576
rect 58157 41518 60000 41520
rect 58157 41515 58223 41518
rect 59200 41488 60000 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 0 41080 800 41200
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 58157 40218 58223 40221
rect 59200 40218 60000 40248
rect 58157 40216 60000 40218
rect 58157 40160 58162 40216
rect 58218 40160 60000 40216
rect 58157 40158 60000 40160
rect 58157 40155 58223 40158
rect 59200 40128 60000 40158
rect 4210 39744 4526 39745
rect 0 39584 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4705 38994 4771 38997
rect 6729 38994 6795 38997
rect 4705 38992 6795 38994
rect 4705 38936 4710 38992
rect 4766 38936 6734 38992
rect 6790 38936 6795 38992
rect 4705 38934 6795 38936
rect 4705 38931 4771 38934
rect 6729 38931 6795 38934
rect 58157 38858 58223 38861
rect 59200 38858 60000 38888
rect 58157 38856 60000 38858
rect 58157 38800 58162 38856
rect 58218 38800 60000 38856
rect 58157 38798 60000 38800
rect 58157 38795 58223 38798
rect 59200 38768 60000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 0 38088 800 38208
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 58157 37498 58223 37501
rect 59200 37498 60000 37528
rect 58157 37496 60000 37498
rect 58157 37440 58162 37496
rect 58218 37440 60000 37496
rect 58157 37438 60000 37440
rect 58157 37435 58223 37438
rect 59200 37408 60000 37438
rect 22686 37300 22692 37364
rect 22756 37362 22762 37364
rect 30649 37362 30715 37365
rect 22756 37360 30715 37362
rect 22756 37304 30654 37360
rect 30710 37304 30715 37360
rect 22756 37302 30715 37304
rect 22756 37300 22762 37302
rect 30649 37299 30715 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 0 36592 800 36712
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 58157 36138 58223 36141
rect 59200 36138 60000 36168
rect 58157 36136 60000 36138
rect 58157 36080 58162 36136
rect 58218 36080 60000 36136
rect 58157 36078 60000 36080
rect 58157 36075 58223 36078
rect 59200 36048 60000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 35096 800 35216
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 58157 34778 58223 34781
rect 59200 34778 60000 34808
rect 58157 34776 60000 34778
rect 58157 34720 58162 34776
rect 58218 34720 60000 34776
rect 58157 34718 60000 34720
rect 58157 34715 58223 34718
rect 59200 34688 60000 34718
rect 12617 34642 12683 34645
rect 18965 34642 19031 34645
rect 19425 34642 19491 34645
rect 12617 34640 19491 34642
rect 12617 34584 12622 34640
rect 12678 34584 18970 34640
rect 19026 34584 19430 34640
rect 19486 34584 19491 34640
rect 12617 34582 19491 34584
rect 12617 34579 12683 34582
rect 18965 34579 19031 34582
rect 19425 34579 19491 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 5533 33962 5599 33965
rect 5809 33962 5875 33965
rect 26693 33962 26759 33965
rect 5533 33960 26759 33962
rect 5533 33904 5538 33960
rect 5594 33904 5814 33960
rect 5870 33904 26698 33960
rect 26754 33904 26759 33960
rect 5533 33902 26759 33904
rect 5533 33899 5599 33902
rect 5809 33899 5875 33902
rect 26693 33899 26759 33902
rect 19570 33760 19886 33761
rect 0 33600 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 14457 33554 14523 33557
rect 17401 33554 17467 33557
rect 14457 33552 17467 33554
rect 14457 33496 14462 33552
rect 14518 33496 17406 33552
rect 17462 33496 17467 33552
rect 14457 33494 17467 33496
rect 14457 33491 14523 33494
rect 17401 33491 17467 33494
rect 58157 33418 58223 33421
rect 59200 33418 60000 33448
rect 58157 33416 60000 33418
rect 58157 33360 58162 33416
rect 58218 33360 60000 33416
rect 58157 33358 60000 33360
rect 58157 33355 58223 33358
rect 59200 33328 60000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 11830 33084 11836 33148
rect 11900 33146 11906 33148
rect 13169 33146 13235 33149
rect 11900 33144 13235 33146
rect 11900 33088 13174 33144
rect 13230 33088 13235 33144
rect 11900 33086 13235 33088
rect 11900 33084 11906 33086
rect 13169 33083 13235 33086
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32104 800 32224
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 58157 32058 58223 32061
rect 59200 32058 60000 32088
rect 58157 32056 60000 32058
rect 58157 32000 58162 32056
rect 58218 32000 60000 32056
rect 58157 31998 60000 32000
rect 58157 31995 58223 31998
rect 59200 31968 60000 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 0 30608 800 30728
rect 58157 30698 58223 30701
rect 59200 30698 60000 30728
rect 58157 30696 60000 30698
rect 58157 30640 58162 30696
rect 58218 30640 60000 30696
rect 58157 30638 60000 30640
rect 58157 30635 58223 30638
rect 59200 30608 60000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 25497 29746 25563 29749
rect 31477 29746 31543 29749
rect 25497 29744 31543 29746
rect 25497 29688 25502 29744
rect 25558 29688 31482 29744
rect 31538 29688 31543 29744
rect 25497 29686 31543 29688
rect 25497 29683 25563 29686
rect 31477 29683 31543 29686
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 58157 29338 58223 29341
rect 59200 29338 60000 29368
rect 58157 29336 60000 29338
rect 58157 29280 58162 29336
rect 58218 29280 60000 29336
rect 58157 29278 60000 29280
rect 58157 29275 58223 29278
rect 59200 29248 60000 29278
rect 0 29112 800 29232
rect 8569 29202 8635 29205
rect 9581 29202 9647 29205
rect 8569 29200 9647 29202
rect 8569 29144 8574 29200
rect 8630 29144 9586 29200
rect 9642 29144 9647 29200
rect 8569 29142 9647 29144
rect 8569 29139 8635 29142
rect 9581 29139 9647 29142
rect 23749 29202 23815 29205
rect 24393 29202 24459 29205
rect 23749 29200 24459 29202
rect 23749 29144 23754 29200
rect 23810 29144 24398 29200
rect 24454 29144 24459 29200
rect 23749 29142 24459 29144
rect 23749 29139 23815 29142
rect 24393 29139 24459 29142
rect 26141 29066 26207 29069
rect 27521 29066 27587 29069
rect 26141 29064 27587 29066
rect 26141 29008 26146 29064
rect 26202 29008 27526 29064
rect 27582 29008 27587 29064
rect 26141 29006 27587 29008
rect 26141 29003 26207 29006
rect 27521 29003 27587 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 58157 27978 58223 27981
rect 59200 27978 60000 28008
rect 58157 27976 60000 27978
rect 58157 27920 58162 27976
rect 58218 27920 60000 27976
rect 58157 27918 60000 27920
rect 58157 27915 58223 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 0 27616 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 58157 26618 58223 26621
rect 59200 26618 60000 26648
rect 58157 26616 60000 26618
rect 58157 26560 58162 26616
rect 58218 26560 60000 26616
rect 58157 26558 60000 26560
rect 58157 26555 58223 26558
rect 59200 26528 60000 26558
rect 21725 26346 21791 26349
rect 22461 26346 22527 26349
rect 21725 26344 22527 26346
rect 21725 26288 21730 26344
rect 21786 26288 22466 26344
rect 22522 26288 22527 26344
rect 21725 26286 22527 26288
rect 21725 26283 21791 26286
rect 22461 26283 22527 26286
rect 0 26120 800 26240
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 58157 25258 58223 25261
rect 59200 25258 60000 25288
rect 58157 25256 60000 25258
rect 58157 25200 58162 25256
rect 58218 25200 60000 25256
rect 58157 25198 60000 25200
rect 58157 25195 58223 25198
rect 59200 25168 60000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 0 24624 800 24744
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 12893 24170 12959 24173
rect 14825 24170 14891 24173
rect 12893 24168 14891 24170
rect 12893 24112 12898 24168
rect 12954 24112 14830 24168
rect 14886 24112 14891 24168
rect 12893 24110 14891 24112
rect 12893 24107 12959 24110
rect 14825 24107 14891 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 58157 23898 58223 23901
rect 59200 23898 60000 23928
rect 58157 23896 60000 23898
rect 58157 23840 58162 23896
rect 58218 23840 60000 23896
rect 58157 23838 60000 23840
rect 58157 23835 58223 23838
rect 59200 23808 60000 23838
rect 21633 23762 21699 23765
rect 22645 23762 22711 23765
rect 21633 23760 22711 23762
rect 21633 23704 21638 23760
rect 21694 23704 22650 23760
rect 22706 23704 22711 23760
rect 21633 23702 22711 23704
rect 21633 23699 21699 23702
rect 22645 23699 22711 23702
rect 17217 23626 17283 23629
rect 18505 23626 18571 23629
rect 17217 23624 18571 23626
rect 17217 23568 17222 23624
rect 17278 23568 18510 23624
rect 18566 23568 18571 23624
rect 17217 23566 18571 23568
rect 17217 23563 17283 23566
rect 18505 23563 18571 23566
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23128 800 23248
rect 2681 23082 2747 23085
rect 3049 23082 3115 23085
rect 2681 23080 3115 23082
rect 2681 23024 2686 23080
rect 2742 23024 3054 23080
rect 3110 23024 3115 23080
rect 2681 23022 3115 23024
rect 2681 23019 2747 23022
rect 3049 23019 3115 23022
rect 6678 23020 6684 23084
rect 6748 23082 6754 23084
rect 20437 23082 20503 23085
rect 6748 23080 20503 23082
rect 6748 23024 20442 23080
rect 20498 23024 20503 23080
rect 6748 23022 20503 23024
rect 6748 23020 6754 23022
rect 20437 23019 20503 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 31753 22538 31819 22541
rect 34329 22538 34395 22541
rect 31753 22536 34395 22538
rect 31753 22480 31758 22536
rect 31814 22480 34334 22536
rect 34390 22480 34395 22536
rect 31753 22478 34395 22480
rect 31753 22475 31819 22478
rect 34329 22475 34395 22478
rect 58157 22538 58223 22541
rect 59200 22538 60000 22568
rect 58157 22536 60000 22538
rect 58157 22480 58162 22536
rect 58218 22480 60000 22536
rect 58157 22478 60000 22480
rect 58157 22475 58223 22478
rect 59200 22448 60000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 30833 21994 30899 21997
rect 32765 21994 32831 21997
rect 30833 21992 32831 21994
rect 30833 21936 30838 21992
rect 30894 21936 32770 21992
rect 32826 21936 32831 21992
rect 30833 21934 32831 21936
rect 30833 21931 30899 21934
rect 32765 21931 32831 21934
rect 19570 21792 19886 21793
rect 0 21632 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 58157 21178 58223 21181
rect 59200 21178 60000 21208
rect 58157 21176 60000 21178
rect 58157 21120 58162 21176
rect 58218 21120 60000 21176
rect 58157 21118 60000 21120
rect 58157 21115 58223 21118
rect 59200 21088 60000 21118
rect 20161 20770 20227 20773
rect 21817 20770 21883 20773
rect 20161 20768 21883 20770
rect 20161 20712 20166 20768
rect 20222 20712 21822 20768
rect 21878 20712 21883 20768
rect 20161 20710 21883 20712
rect 20161 20707 20227 20710
rect 21817 20707 21883 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 19425 20634 19491 20637
rect 19290 20632 19491 20634
rect 19290 20576 19430 20632
rect 19486 20576 19491 20632
rect 19290 20574 19491 20576
rect 19290 20362 19350 20574
rect 19425 20571 19491 20574
rect 19425 20498 19491 20501
rect 20529 20498 20595 20501
rect 19425 20496 20595 20498
rect 19425 20440 19430 20496
rect 19486 20440 20534 20496
rect 20590 20440 20595 20496
rect 19425 20438 20595 20440
rect 19425 20435 19491 20438
rect 20529 20435 20595 20438
rect 19793 20362 19859 20365
rect 19290 20360 19859 20362
rect 19290 20304 19798 20360
rect 19854 20304 19859 20360
rect 19290 20302 19859 20304
rect 19793 20299 19859 20302
rect 0 20136 800 20256
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 15193 19954 15259 19957
rect 26969 19954 27035 19957
rect 15193 19952 27035 19954
rect 15193 19896 15198 19952
rect 15254 19896 26974 19952
rect 27030 19896 27035 19952
rect 15193 19894 27035 19896
rect 15193 19891 15259 19894
rect 26969 19891 27035 19894
rect 9857 19818 9923 19821
rect 30925 19818 30991 19821
rect 9857 19816 30991 19818
rect 9857 19760 9862 19816
rect 9918 19760 30930 19816
rect 30986 19760 30991 19816
rect 9857 19758 30991 19760
rect 9857 19755 9923 19758
rect 30925 19755 30991 19758
rect 58157 19818 58223 19821
rect 59200 19818 60000 19848
rect 58157 19816 60000 19818
rect 58157 19760 58162 19816
rect 58218 19760 60000 19816
rect 58157 19758 60000 19760
rect 58157 19755 58223 19758
rect 59200 19728 60000 19758
rect 25589 19682 25655 19685
rect 28901 19682 28967 19685
rect 25589 19680 28967 19682
rect 25589 19624 25594 19680
rect 25650 19624 28906 19680
rect 28962 19624 28967 19680
rect 25589 19622 28967 19624
rect 25589 19619 25655 19622
rect 28901 19619 28967 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 8293 18866 8359 18869
rect 30649 18866 30715 18869
rect 8293 18864 30715 18866
rect 8293 18808 8298 18864
rect 8354 18808 30654 18864
rect 30710 18808 30715 18864
rect 8293 18806 30715 18808
rect 8293 18803 8359 18806
rect 30649 18803 30715 18806
rect 0 18640 800 18760
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 58157 18458 58223 18461
rect 59200 18458 60000 18488
rect 58157 18456 60000 18458
rect 58157 18400 58162 18456
rect 58218 18400 60000 18456
rect 58157 18398 60000 18400
rect 58157 18395 58223 18398
rect 59200 18368 60000 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 17144 800 17264
rect 25957 17234 26023 17237
rect 37222 17234 37228 17236
rect 25957 17232 37228 17234
rect 25957 17176 25962 17232
rect 26018 17176 37228 17232
rect 25957 17174 37228 17176
rect 25957 17171 26023 17174
rect 37222 17172 37228 17174
rect 37292 17172 37298 17236
rect 58157 17098 58223 17101
rect 59200 17098 60000 17128
rect 58157 17096 60000 17098
rect 58157 17040 58162 17096
rect 58218 17040 60000 17096
rect 58157 17038 60000 17040
rect 58157 17035 58223 17038
rect 59200 17008 60000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 37273 16012 37339 16013
rect 37222 15948 37228 16012
rect 37292 16010 37339 16012
rect 37292 16008 37384 16010
rect 37334 15952 37384 16008
rect 37292 15950 37384 15952
rect 37292 15948 37339 15950
rect 37273 15947 37339 15948
rect 4210 15808 4526 15809
rect 0 15648 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 58157 15738 58223 15741
rect 59200 15738 60000 15768
rect 58157 15736 60000 15738
rect 58157 15680 58162 15736
rect 58218 15680 60000 15736
rect 58157 15678 60000 15680
rect 58157 15675 58223 15678
rect 59200 15648 60000 15678
rect 10041 15602 10107 15605
rect 24025 15602 24091 15605
rect 10041 15600 24091 15602
rect 10041 15544 10046 15600
rect 10102 15544 24030 15600
rect 24086 15544 24091 15600
rect 10041 15542 24091 15544
rect 10041 15539 10107 15542
rect 24025 15539 24091 15542
rect 10501 15466 10567 15469
rect 10777 15466 10843 15469
rect 12985 15466 13051 15469
rect 10501 15464 13051 15466
rect 10501 15408 10506 15464
rect 10562 15408 10782 15464
rect 10838 15408 12990 15464
rect 13046 15408 13051 15464
rect 10501 15406 13051 15408
rect 10501 15403 10567 15406
rect 10777 15403 10843 15406
rect 12985 15403 13051 15406
rect 4797 15332 4863 15333
rect 4797 15330 4844 15332
rect 4752 15328 4844 15330
rect 4752 15272 4802 15328
rect 4752 15270 4844 15272
rect 4797 15268 4844 15270
rect 4908 15268 4914 15332
rect 4797 15267 4863 15268
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 58157 14378 58223 14381
rect 59200 14378 60000 14408
rect 58157 14376 60000 14378
rect 58157 14320 58162 14376
rect 58218 14320 60000 14376
rect 58157 14318 60000 14320
rect 58157 14315 58223 14318
rect 59200 14288 60000 14318
rect 0 14152 800 14272
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 8109 13834 8175 13837
rect 23933 13834 23999 13837
rect 8109 13832 23999 13834
rect 8109 13776 8114 13832
rect 8170 13776 23938 13832
rect 23994 13776 23999 13832
rect 8109 13774 23999 13776
rect 8109 13771 8175 13774
rect 23933 13771 23999 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 12249 13290 12315 13293
rect 22921 13290 22987 13293
rect 12249 13288 22987 13290
rect 12249 13232 12254 13288
rect 12310 13232 22926 13288
rect 22982 13232 22987 13288
rect 12249 13230 22987 13232
rect 12249 13227 12315 13230
rect 22921 13227 22987 13230
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 58157 13018 58223 13021
rect 59200 13018 60000 13048
rect 58157 13016 60000 13018
rect 58157 12960 58162 13016
rect 58218 12960 60000 13016
rect 58157 12958 60000 12960
rect 58157 12955 58223 12958
rect 59200 12928 60000 12958
rect 0 12656 800 12776
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 22737 12202 22803 12205
rect 25497 12202 25563 12205
rect 22737 12200 25563 12202
rect 22737 12144 22742 12200
rect 22798 12144 25502 12200
rect 25558 12144 25563 12200
rect 22737 12142 25563 12144
rect 22737 12139 22803 12142
rect 25497 12139 25563 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 58157 11658 58223 11661
rect 59200 11658 60000 11688
rect 58157 11656 60000 11658
rect 58157 11600 58162 11656
rect 58218 11600 60000 11656
rect 58157 11598 60000 11600
rect 58157 11595 58223 11598
rect 59200 11568 60000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 11160 800 11280
rect 5942 11052 5948 11116
rect 6012 11114 6018 11116
rect 9673 11114 9739 11117
rect 6012 11112 9739 11114
rect 6012 11056 9678 11112
rect 9734 11056 9739 11112
rect 6012 11054 9739 11056
rect 6012 11052 6018 11054
rect 9673 11051 9739 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 7097 10842 7163 10845
rect 8334 10842 8340 10844
rect 7097 10840 8340 10842
rect 7097 10784 7102 10840
rect 7158 10784 8340 10840
rect 7097 10782 8340 10784
rect 7097 10779 7163 10782
rect 8334 10780 8340 10782
rect 8404 10780 8410 10844
rect 10358 10508 10364 10572
rect 10428 10570 10434 10572
rect 10593 10570 10659 10573
rect 28533 10570 28599 10573
rect 10428 10568 10659 10570
rect 10428 10512 10598 10568
rect 10654 10512 10659 10568
rect 10428 10510 10659 10512
rect 10428 10508 10434 10510
rect 10593 10507 10659 10510
rect 12390 10568 28599 10570
rect 12390 10512 28538 10568
rect 28594 10512 28599 10568
rect 12390 10510 28599 10512
rect 9397 10434 9463 10437
rect 12390 10434 12450 10510
rect 28533 10507 28599 10510
rect 9397 10432 12450 10434
rect 9397 10376 9402 10432
rect 9458 10376 12450 10432
rect 9397 10374 12450 10376
rect 9397 10371 9463 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 58157 10298 58223 10301
rect 59200 10298 60000 10328
rect 58157 10296 60000 10298
rect 58157 10240 58162 10296
rect 58218 10240 60000 10296
rect 58157 10238 60000 10240
rect 58157 10235 58223 10238
rect 59200 10208 60000 10238
rect 9397 10026 9463 10029
rect 9622 10026 9628 10028
rect 9397 10024 9628 10026
rect 9397 9968 9402 10024
rect 9458 9968 9628 10024
rect 9397 9966 9628 9968
rect 9397 9963 9463 9966
rect 9622 9964 9628 9966
rect 9692 9964 9698 10028
rect 19570 9824 19886 9825
rect 0 9664 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 58157 8938 58223 8941
rect 59200 8938 60000 8968
rect 58157 8936 60000 8938
rect 58157 8880 58162 8936
rect 58218 8880 60000 8936
rect 58157 8878 60000 8880
rect 58157 8875 58223 8878
rect 59200 8848 60000 8878
rect 2773 8802 2839 8805
rect 8518 8802 8524 8804
rect 2773 8800 8524 8802
rect 2773 8744 2778 8800
rect 2834 8744 8524 8800
rect 2773 8742 8524 8744
rect 2773 8739 2839 8742
rect 8518 8740 8524 8742
rect 8588 8740 8594 8804
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 16757 8530 16823 8533
rect 17953 8530 18019 8533
rect 16757 8528 18019 8530
rect 16757 8472 16762 8528
rect 16818 8472 17958 8528
rect 18014 8472 18019 8528
rect 16757 8470 18019 8472
rect 16757 8467 16823 8470
rect 17953 8467 18019 8470
rect 37273 8530 37339 8533
rect 38837 8530 38903 8533
rect 37273 8528 38903 8530
rect 37273 8472 37278 8528
rect 37334 8472 38842 8528
rect 38898 8472 38903 8528
rect 37273 8470 38903 8472
rect 37273 8467 37339 8470
rect 38837 8467 38903 8470
rect 6821 8396 6887 8397
rect 6821 8392 6868 8396
rect 6932 8394 6938 8396
rect 6821 8336 6826 8392
rect 6821 8332 6868 8336
rect 6932 8334 6978 8394
rect 6932 8332 6938 8334
rect 6821 8331 6887 8332
rect 0 8168 800 8288
rect 9438 8196 9444 8260
rect 9508 8258 9514 8260
rect 16021 8258 16087 8261
rect 9508 8256 16087 8258
rect 9508 8200 16026 8256
rect 16082 8200 16087 8256
rect 9508 8198 16087 8200
rect 9508 8196 9514 8198
rect 16021 8195 16087 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 9581 8122 9647 8125
rect 9806 8122 9812 8124
rect 9581 8120 9812 8122
rect 9581 8064 9586 8120
rect 9642 8064 9812 8120
rect 9581 8062 9812 8064
rect 9581 8059 9647 8062
rect 9806 8060 9812 8062
rect 9876 8122 9882 8124
rect 17677 8122 17743 8125
rect 9876 8120 17743 8122
rect 9876 8064 17682 8120
rect 17738 8064 17743 8120
rect 9876 8062 17743 8064
rect 9876 8060 9882 8062
rect 17677 8059 17743 8062
rect 1577 7986 1643 7989
rect 2814 7986 2820 7988
rect 1577 7984 2820 7986
rect 1577 7928 1582 7984
rect 1638 7928 2820 7984
rect 1577 7926 2820 7928
rect 1577 7923 1643 7926
rect 2814 7924 2820 7926
rect 2884 7924 2890 7988
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 11881 7580 11947 7581
rect 11830 7516 11836 7580
rect 11900 7578 11947 7580
rect 58157 7578 58223 7581
rect 59200 7578 60000 7608
rect 11900 7576 11992 7578
rect 11942 7520 11992 7576
rect 11900 7518 11992 7520
rect 58157 7576 60000 7578
rect 58157 7520 58162 7576
rect 58218 7520 60000 7576
rect 58157 7518 60000 7520
rect 11900 7516 11947 7518
rect 11881 7515 11947 7516
rect 58157 7515 58223 7518
rect 59200 7488 60000 7518
rect 4654 7244 4660 7308
rect 4724 7306 4730 7308
rect 5625 7306 5691 7309
rect 8385 7306 8451 7309
rect 4724 7304 8451 7306
rect 4724 7248 5630 7304
rect 5686 7248 8390 7304
rect 8446 7248 8451 7304
rect 4724 7246 8451 7248
rect 4724 7244 4730 7246
rect 5625 7243 5691 7246
rect 8385 7243 8451 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6672 800 6792
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 12801 6354 12867 6357
rect 13537 6354 13603 6357
rect 26969 6354 27035 6357
rect 12801 6352 27035 6354
rect 12801 6296 12806 6352
rect 12862 6296 13542 6352
rect 13598 6296 26974 6352
rect 27030 6296 27035 6352
rect 12801 6294 27035 6296
rect 12801 6291 12867 6294
rect 13537 6291 13603 6294
rect 26969 6291 27035 6294
rect 58157 6218 58223 6221
rect 59200 6218 60000 6248
rect 58157 6216 60000 6218
rect 58157 6160 58162 6216
rect 58218 6160 60000 6216
rect 58157 6158 60000 6160
rect 58157 6155 58223 6158
rect 59200 6128 60000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 20437 5674 20503 5677
rect 23974 5674 23980 5676
rect 20437 5672 23980 5674
rect 20437 5616 20442 5672
rect 20498 5616 23980 5672
rect 20437 5614 23980 5616
rect 20437 5611 20503 5614
rect 23974 5612 23980 5614
rect 24044 5612 24050 5676
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 8518 5340 8524 5404
rect 8588 5402 8594 5404
rect 8588 5342 9690 5402
rect 8588 5340 8594 5342
rect 0 5176 800 5296
rect 9630 5269 9690 5342
rect 2773 5266 2839 5269
rect 9438 5266 9444 5268
rect 2773 5264 9444 5266
rect 2773 5208 2778 5264
rect 2834 5208 9444 5264
rect 2773 5206 9444 5208
rect 2773 5203 2839 5206
rect 9438 5204 9444 5206
rect 9508 5204 9514 5268
rect 9581 5266 9690 5269
rect 26417 5266 26483 5269
rect 9581 5264 26483 5266
rect 9581 5208 9586 5264
rect 9642 5208 26422 5264
rect 26478 5208 26483 5264
rect 9581 5206 26483 5208
rect 9581 5203 9647 5206
rect 26417 5203 26483 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 58157 4858 58223 4861
rect 59200 4858 60000 4888
rect 58157 4856 60000 4858
rect 58157 4800 58162 4856
rect 58218 4800 60000 4856
rect 58157 4798 60000 4800
rect 58157 4795 58223 4798
rect 59200 4768 60000 4798
rect 4337 4722 4403 4725
rect 4654 4722 4660 4724
rect 4337 4720 4660 4722
rect 4337 4664 4342 4720
rect 4398 4664 4660 4720
rect 4337 4662 4660 4664
rect 4337 4659 4403 4662
rect 4654 4660 4660 4662
rect 4724 4660 4730 4724
rect 5257 4450 5323 4453
rect 8845 4450 8911 4453
rect 5257 4448 8911 4450
rect 5257 4392 5262 4448
rect 5318 4392 8850 4448
rect 8906 4392 8911 4448
rect 5257 4390 8911 4392
rect 5257 4387 5323 4390
rect 8845 4387 8911 4390
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4889 4314 4955 4317
rect 5257 4314 5323 4317
rect 4889 4312 5323 4314
rect 4889 4256 4894 4312
rect 4950 4256 5262 4312
rect 5318 4256 5323 4312
rect 4889 4254 5323 4256
rect 4889 4251 4955 4254
rect 5257 4251 5323 4254
rect 3141 4042 3207 4045
rect 6453 4042 6519 4045
rect 3141 4040 6519 4042
rect 3141 3984 3146 4040
rect 3202 3984 6458 4040
rect 6514 3984 6519 4040
rect 3141 3982 6519 3984
rect 3141 3979 3207 3982
rect 6453 3979 6519 3982
rect 6862 3980 6868 4044
rect 6932 4042 6938 4044
rect 7097 4042 7163 4045
rect 6932 4040 7163 4042
rect 6932 3984 7102 4040
rect 7158 3984 7163 4040
rect 6932 3982 7163 3984
rect 6932 3980 6938 3982
rect 7097 3979 7163 3982
rect 8334 3980 8340 4044
rect 8404 4042 8410 4044
rect 9397 4042 9463 4045
rect 9673 4044 9739 4045
rect 9622 4042 9628 4044
rect 8404 4040 9463 4042
rect 8404 3984 9402 4040
rect 9458 3984 9463 4040
rect 8404 3982 9463 3984
rect 9582 3982 9628 4042
rect 9692 4040 9739 4044
rect 9734 3984 9739 4040
rect 8404 3980 8410 3982
rect 9397 3979 9463 3982
rect 9622 3980 9628 3982
rect 9692 3980 9739 3984
rect 9673 3979 9739 3980
rect 14457 4042 14523 4045
rect 14590 4042 14596 4044
rect 14457 4040 14596 4042
rect 14457 3984 14462 4040
rect 14518 3984 14596 4040
rect 14457 3982 14596 3984
rect 14457 3979 14523 3982
rect 14590 3980 14596 3982
rect 14660 3980 14666 4044
rect 20345 4042 20411 4045
rect 20478 4042 20484 4044
rect 20345 4040 20484 4042
rect 20345 3984 20350 4040
rect 20406 3984 20484 4040
rect 20345 3982 20484 3984
rect 20345 3979 20411 3982
rect 20478 3980 20484 3982
rect 20548 3980 20554 4044
rect 9305 3906 9371 3909
rect 9438 3906 9444 3908
rect 9305 3904 9444 3906
rect 9305 3848 9310 3904
rect 9366 3848 9444 3904
rect 9305 3846 9444 3848
rect 9305 3843 9371 3846
rect 9438 3844 9444 3846
rect 9508 3844 9514 3908
rect 4210 3840 4526 3841
rect 0 3680 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 9765 3772 9831 3773
rect 21909 3772 21975 3773
rect 9765 3770 9812 3772
rect 9720 3768 9812 3770
rect 9720 3712 9770 3768
rect 9720 3710 9812 3712
rect 9765 3708 9812 3710
rect 9876 3708 9882 3772
rect 21909 3770 21956 3772
rect 21864 3768 21956 3770
rect 21864 3712 21914 3768
rect 21864 3710 21956 3712
rect 21909 3708 21956 3710
rect 22020 3708 22026 3772
rect 9765 3707 9831 3708
rect 21909 3707 21975 3708
rect 3969 3634 4035 3637
rect 6177 3634 6243 3637
rect 3969 3632 6243 3634
rect 3969 3576 3974 3632
rect 4030 3576 6182 3632
rect 6238 3576 6243 3632
rect 3969 3574 6243 3576
rect 3969 3571 4035 3574
rect 6177 3571 6243 3574
rect 2129 3498 2195 3501
rect 9213 3498 9279 3501
rect 2129 3496 9279 3498
rect 2129 3440 2134 3496
rect 2190 3440 9218 3496
rect 9274 3440 9279 3496
rect 2129 3438 9279 3440
rect 2129 3435 2195 3438
rect 9213 3435 9279 3438
rect 58157 3498 58223 3501
rect 59200 3498 60000 3528
rect 58157 3496 60000 3498
rect 58157 3440 58162 3496
rect 58218 3440 60000 3496
rect 58157 3438 60000 3440
rect 58157 3435 58223 3438
rect 59200 3408 60000 3438
rect 3325 3362 3391 3365
rect 10685 3362 10751 3365
rect 3325 3360 10751 3362
rect 3325 3304 3330 3360
rect 3386 3304 10690 3360
rect 10746 3304 10751 3360
rect 3325 3302 10751 3304
rect 3325 3299 3391 3302
rect 10685 3299 10751 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 6821 3226 6887 3229
rect 14917 3226 14983 3229
rect 18229 3228 18295 3229
rect 18229 3226 18276 3228
rect 6821 3224 14983 3226
rect 6821 3168 6826 3224
rect 6882 3168 14922 3224
rect 14978 3168 14983 3224
rect 6821 3166 14983 3168
rect 18184 3224 18276 3226
rect 18184 3168 18234 3224
rect 18184 3166 18276 3168
rect 6821 3163 6887 3166
rect 14917 3163 14983 3166
rect 18229 3164 18276 3166
rect 18340 3164 18346 3228
rect 18873 3226 18939 3229
rect 19006 3226 19012 3228
rect 18873 3224 19012 3226
rect 18873 3168 18878 3224
rect 18934 3168 19012 3224
rect 18873 3166 19012 3168
rect 18229 3163 18295 3164
rect 18873 3163 18939 3166
rect 19006 3164 19012 3166
rect 19076 3164 19082 3228
rect 21081 3226 21147 3229
rect 21214 3226 21220 3228
rect 21081 3224 21220 3226
rect 21081 3168 21086 3224
rect 21142 3168 21220 3224
rect 21081 3166 21220 3168
rect 21081 3163 21147 3166
rect 21214 3164 21220 3166
rect 21284 3164 21290 3228
rect 13721 3090 13787 3093
rect 15469 3090 15535 3093
rect 13721 3088 15535 3090
rect 13721 3032 13726 3088
rect 13782 3032 15474 3088
rect 15530 3032 15535 3088
rect 13721 3030 15535 3032
rect 13721 3027 13787 3030
rect 15469 3027 15535 3030
rect 2221 2954 2287 2957
rect 6913 2954 6979 2957
rect 2221 2952 6979 2954
rect 2221 2896 2226 2952
rect 2282 2896 6918 2952
rect 6974 2896 6979 2952
rect 2221 2894 6979 2896
rect 2221 2891 2287 2894
rect 6913 2891 6979 2894
rect 7281 2954 7347 2957
rect 7925 2954 7991 2957
rect 7281 2952 7482 2954
rect 7281 2896 7286 2952
rect 7342 2896 7482 2952
rect 7281 2894 7482 2896
rect 7281 2891 7347 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 2814 2620 2820 2684
rect 2884 2682 2890 2684
rect 2957 2682 3023 2685
rect 2884 2680 3023 2682
rect 2884 2624 2962 2680
rect 3018 2624 3023 2680
rect 2884 2622 3023 2624
rect 7422 2682 7482 2894
rect 7790 2952 7991 2954
rect 7790 2896 7930 2952
rect 7986 2896 7991 2952
rect 7790 2894 7991 2896
rect 7649 2818 7715 2821
rect 7790 2818 7850 2894
rect 7925 2891 7991 2894
rect 53373 2954 53439 2957
rect 56593 2954 56659 2957
rect 53373 2952 56659 2954
rect 53373 2896 53378 2952
rect 53434 2896 56598 2952
rect 56654 2896 56659 2952
rect 53373 2894 56659 2896
rect 53373 2891 53439 2894
rect 56593 2891 56659 2894
rect 7649 2816 7850 2818
rect 7649 2760 7654 2816
rect 7710 2760 7850 2816
rect 7649 2758 7850 2760
rect 53465 2818 53531 2821
rect 55305 2818 55371 2821
rect 53465 2816 55371 2818
rect 53465 2760 53470 2816
rect 53526 2760 55310 2816
rect 55366 2760 55371 2816
rect 53465 2758 55371 2760
rect 7649 2755 7715 2758
rect 53465 2755 53531 2758
rect 55305 2755 55371 2758
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 7557 2682 7623 2685
rect 7422 2680 7623 2682
rect 7422 2624 7562 2680
rect 7618 2624 7623 2680
rect 7422 2622 7623 2624
rect 2884 2620 2890 2622
rect 2957 2619 3023 2622
rect 7557 2619 7623 2622
rect 14549 2682 14615 2685
rect 15694 2682 15700 2684
rect 14549 2680 15700 2682
rect 14549 2624 14554 2680
rect 14610 2624 15700 2680
rect 14549 2622 15700 2624
rect 14549 2619 14615 2622
rect 15694 2620 15700 2622
rect 15764 2620 15770 2684
rect 16297 2682 16363 2685
rect 17166 2682 17172 2684
rect 16297 2680 17172 2682
rect 16297 2624 16302 2680
rect 16358 2624 17172 2680
rect 16297 2622 17172 2624
rect 16297 2619 16363 2622
rect 17166 2620 17172 2622
rect 17236 2620 17242 2684
rect 17677 2682 17743 2685
rect 20110 2682 20116 2684
rect 17677 2680 20116 2682
rect 17677 2624 17682 2680
rect 17738 2624 20116 2680
rect 17677 2622 20116 2624
rect 17677 2619 17743 2622
rect 20110 2620 20116 2622
rect 20180 2620 20186 2684
rect 5809 2546 5875 2549
rect 5942 2546 5948 2548
rect 5809 2544 5948 2546
rect 5809 2488 5814 2544
rect 5870 2488 5948 2544
rect 5809 2486 5948 2488
rect 5809 2483 5875 2486
rect 5942 2484 5948 2486
rect 6012 2484 6018 2548
rect 18505 2546 18571 2549
rect 22686 2546 22692 2548
rect 18505 2544 22692 2546
rect 18505 2488 18510 2544
rect 18566 2488 22692 2544
rect 18505 2486 22692 2488
rect 18505 2483 18571 2486
rect 22686 2484 22692 2486
rect 22756 2484 22762 2548
rect 4245 2410 4311 2413
rect 4838 2410 4844 2412
rect 4245 2408 4844 2410
rect 4245 2352 4250 2408
rect 4306 2352 4844 2408
rect 4245 2350 4844 2352
rect 4245 2347 4311 2350
rect 4838 2348 4844 2350
rect 4908 2348 4914 2412
rect 5533 2410 5599 2413
rect 10409 2412 10475 2413
rect 6678 2410 6684 2412
rect 5533 2408 6684 2410
rect 5533 2352 5538 2408
rect 5594 2352 6684 2408
rect 5533 2350 6684 2352
rect 5533 2347 5599 2350
rect 6678 2348 6684 2350
rect 6748 2348 6754 2412
rect 10358 2410 10364 2412
rect 10318 2350 10364 2410
rect 10428 2408 10475 2412
rect 10470 2352 10475 2408
rect 10358 2348 10364 2350
rect 10428 2348 10475 2352
rect 10409 2347 10475 2348
rect 16021 2410 16087 2413
rect 23238 2410 23244 2412
rect 16021 2408 23244 2410
rect 16021 2352 16026 2408
rect 16082 2352 23244 2408
rect 16021 2350 23244 2352
rect 16021 2347 16087 2350
rect 23238 2348 23244 2350
rect 23308 2348 23314 2412
rect 0 2184 800 2304
rect 1577 2274 1643 2277
rect 8477 2274 8543 2277
rect 9213 2274 9279 2277
rect 1577 2272 9279 2274
rect 1577 2216 1582 2272
rect 1638 2216 8482 2272
rect 8538 2216 9218 2272
rect 9274 2216 9279 2272
rect 1577 2214 9279 2216
rect 1577 2211 1643 2214
rect 8477 2211 8543 2214
rect 9213 2211 9279 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 57513 2138 57579 2141
rect 59200 2138 60000 2168
rect 57513 2136 60000 2138
rect 57513 2080 57518 2136
rect 57574 2080 60000 2136
rect 57513 2078 60000 2080
rect 57513 2075 57579 2078
rect 59200 2048 60000 2078
rect 58433 778 58499 781
rect 59200 778 60000 808
rect 58433 776 60000 778
rect 58433 720 58438 776
rect 58494 720 60000 776
rect 58433 718 60000 720
rect 58433 715 58499 718
rect 59200 688 60000 718
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 23244 56204 23308 56268
rect 20484 56068 20548 56132
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 23980 55660 24044 55724
rect 14596 55524 14660 55588
rect 15700 55524 15764 55588
rect 17172 55584 17236 55588
rect 17172 55528 17222 55584
rect 17222 55528 17236 55584
rect 17172 55524 17236 55528
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19012 44780 19076 44844
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 18276 43692 18340 43756
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 20116 42332 20180 42396
rect 21956 42196 22020 42260
rect 21220 42060 21284 42124
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 22692 37300 22756 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 11836 33084 11900 33148
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 6684 23020 6748 23084
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 37228 17172 37292 17236
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 37228 16008 37292 16012
rect 37228 15952 37278 16008
rect 37278 15952 37292 16008
rect 37228 15948 37292 15952
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4844 15328 4908 15332
rect 4844 15272 4858 15328
rect 4858 15272 4908 15328
rect 4844 15268 4908 15272
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 5948 11052 6012 11116
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 8340 10780 8404 10844
rect 10364 10508 10428 10572
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 9628 9964 9692 10028
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 8524 8740 8588 8804
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 6868 8392 6932 8396
rect 6868 8336 6882 8392
rect 6882 8336 6932 8392
rect 6868 8332 6932 8336
rect 9444 8196 9508 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 9812 8060 9876 8124
rect 2820 7924 2884 7988
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 11836 7576 11900 7580
rect 11836 7520 11886 7576
rect 11886 7520 11900 7576
rect 11836 7516 11900 7520
rect 4660 7244 4724 7308
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 23980 5612 24044 5676
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 8524 5340 8588 5404
rect 9444 5204 9508 5268
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4660 4660 4724 4724
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 6868 3980 6932 4044
rect 8340 3980 8404 4044
rect 9628 4040 9692 4044
rect 9628 3984 9678 4040
rect 9678 3984 9692 4040
rect 9628 3980 9692 3984
rect 14596 3980 14660 4044
rect 20484 3980 20548 4044
rect 9444 3844 9508 3908
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 9812 3768 9876 3772
rect 9812 3712 9826 3768
rect 9826 3712 9876 3768
rect 9812 3708 9876 3712
rect 21956 3768 22020 3772
rect 21956 3712 21970 3768
rect 21970 3712 22020 3768
rect 21956 3708 22020 3712
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 18276 3224 18340 3228
rect 18276 3168 18290 3224
rect 18290 3168 18340 3224
rect 18276 3164 18340 3168
rect 19012 3164 19076 3228
rect 21220 3164 21284 3228
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 2820 2620 2884 2684
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 15700 2620 15764 2684
rect 17172 2620 17236 2684
rect 20116 2620 20180 2684
rect 5948 2484 6012 2548
rect 22692 2484 22756 2548
rect 4844 2348 4908 2412
rect 6684 2348 6748 2412
rect 10364 2408 10428 2412
rect 10364 2352 10414 2408
rect 10414 2352 10428 2408
rect 10364 2348 10428 2352
rect 23244 2348 23308 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 14595 55588 14661 55589
rect 14595 55524 14596 55588
rect 14660 55524 14661 55588
rect 14595 55523 14661 55524
rect 15699 55588 15765 55589
rect 15699 55524 15700 55588
rect 15764 55524 15765 55588
rect 15699 55523 15765 55524
rect 17171 55588 17237 55589
rect 17171 55524 17172 55588
rect 17236 55524 17237 55588
rect 17171 55523 17237 55524
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 11835 33148 11901 33149
rect 11835 33084 11836 33148
rect 11900 33084 11901 33148
rect 11835 33083 11901 33084
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 6683 23084 6749 23085
rect 6683 23020 6684 23084
rect 6748 23020 6749 23084
rect 6683 23019 6749 23020
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4843 15332 4909 15333
rect 4843 15268 4844 15332
rect 4908 15268 4909 15332
rect 4843 15267 4909 15268
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 2819 7988 2885 7989
rect 2819 7924 2820 7988
rect 2884 7924 2885 7988
rect 2819 7923 2885 7924
rect 2822 2685 2882 7923
rect 4208 7104 4528 8128
rect 4659 7308 4725 7309
rect 4659 7244 4660 7308
rect 4724 7244 4725 7308
rect 4659 7243 4725 7244
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4662 4725 4722 7243
rect 4659 4724 4725 4725
rect 4659 4660 4660 4724
rect 4724 4660 4725 4724
rect 4659 4659 4725 4660
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 2819 2684 2885 2685
rect 2819 2620 2820 2684
rect 2884 2620 2885 2684
rect 2819 2619 2885 2620
rect 4208 2128 4528 2688
rect 4846 2413 4906 15267
rect 5947 11116 6013 11117
rect 5947 11052 5948 11116
rect 6012 11052 6013 11116
rect 5947 11051 6013 11052
rect 5950 2549 6010 11051
rect 5947 2548 6013 2549
rect 5947 2484 5948 2548
rect 6012 2484 6013 2548
rect 5947 2483 6013 2484
rect 6686 2413 6746 23019
rect 8339 10844 8405 10845
rect 8339 10780 8340 10844
rect 8404 10780 8405 10844
rect 8339 10779 8405 10780
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 6870 4045 6930 8331
rect 8342 4045 8402 10779
rect 10363 10572 10429 10573
rect 10363 10508 10364 10572
rect 10428 10508 10429 10572
rect 10363 10507 10429 10508
rect 9627 10028 9693 10029
rect 9627 9964 9628 10028
rect 9692 9964 9693 10028
rect 9627 9963 9693 9964
rect 8523 8804 8589 8805
rect 8523 8740 8524 8804
rect 8588 8740 8589 8804
rect 8523 8739 8589 8740
rect 8526 5405 8586 8739
rect 9443 8260 9509 8261
rect 9443 8196 9444 8260
rect 9508 8196 9509 8260
rect 9443 8195 9509 8196
rect 8523 5404 8589 5405
rect 8523 5340 8524 5404
rect 8588 5340 8589 5404
rect 8523 5339 8589 5340
rect 9446 5269 9506 8195
rect 9443 5268 9509 5269
rect 9443 5204 9444 5268
rect 9508 5204 9509 5268
rect 9443 5203 9509 5204
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 8339 4044 8405 4045
rect 8339 3980 8340 4044
rect 8404 3980 8405 4044
rect 8339 3979 8405 3980
rect 9446 3909 9506 5203
rect 9630 4045 9690 9963
rect 9811 8124 9877 8125
rect 9811 8060 9812 8124
rect 9876 8060 9877 8124
rect 9811 8059 9877 8060
rect 9627 4044 9693 4045
rect 9627 3980 9628 4044
rect 9692 3980 9693 4044
rect 9627 3979 9693 3980
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 9814 3773 9874 8059
rect 9811 3772 9877 3773
rect 9811 3708 9812 3772
rect 9876 3708 9877 3772
rect 9811 3707 9877 3708
rect 10366 2413 10426 10507
rect 11838 7581 11898 33083
rect 11835 7580 11901 7581
rect 11835 7516 11836 7580
rect 11900 7516 11901 7580
rect 11835 7515 11901 7516
rect 14598 4045 14658 55523
rect 14595 4044 14661 4045
rect 14595 3980 14596 4044
rect 14660 3980 14661 4044
rect 14595 3979 14661 3980
rect 15702 2685 15762 55523
rect 17174 2685 17234 55523
rect 19568 55520 19888 56544
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 23243 56268 23309 56269
rect 23243 56204 23244 56268
rect 23308 56204 23309 56268
rect 23243 56203 23309 56204
rect 20483 56132 20549 56133
rect 20483 56068 20484 56132
rect 20548 56068 20549 56132
rect 20483 56067 20549 56068
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19011 44844 19077 44845
rect 19011 44780 19012 44844
rect 19076 44780 19077 44844
rect 19011 44779 19077 44780
rect 18275 43756 18341 43757
rect 18275 43692 18276 43756
rect 18340 43692 18341 43756
rect 18275 43691 18341 43692
rect 18278 3229 18338 43691
rect 19014 3229 19074 44779
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 20115 42396 20181 42397
rect 20115 42332 20116 42396
rect 20180 42332 20181 42396
rect 20115 42331 20181 42332
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 18275 3228 18341 3229
rect 18275 3164 18276 3228
rect 18340 3164 18341 3228
rect 18275 3163 18341 3164
rect 19011 3228 19077 3229
rect 19011 3164 19012 3228
rect 19076 3164 19077 3228
rect 19011 3163 19077 3164
rect 15699 2684 15765 2685
rect 15699 2620 15700 2684
rect 15764 2620 15765 2684
rect 15699 2619 15765 2620
rect 17171 2684 17237 2685
rect 17171 2620 17172 2684
rect 17236 2620 17237 2684
rect 17171 2619 17237 2620
rect 4843 2412 4909 2413
rect 4843 2348 4844 2412
rect 4908 2348 4909 2412
rect 4843 2347 4909 2348
rect 6683 2412 6749 2413
rect 6683 2348 6684 2412
rect 6748 2348 6749 2412
rect 6683 2347 6749 2348
rect 10363 2412 10429 2413
rect 10363 2348 10364 2412
rect 10428 2348 10429 2412
rect 10363 2347 10429 2348
rect 19568 2208 19888 3232
rect 20118 2685 20178 42331
rect 20486 4045 20546 56067
rect 21955 42260 22021 42261
rect 21955 42196 21956 42260
rect 22020 42196 22021 42260
rect 21955 42195 22021 42196
rect 21219 42124 21285 42125
rect 21219 42060 21220 42124
rect 21284 42060 21285 42124
rect 21219 42059 21285 42060
rect 20483 4044 20549 4045
rect 20483 3980 20484 4044
rect 20548 3980 20549 4044
rect 20483 3979 20549 3980
rect 21222 3229 21282 42059
rect 21958 3773 22018 42195
rect 22691 37364 22757 37365
rect 22691 37300 22692 37364
rect 22756 37300 22757 37364
rect 22691 37299 22757 37300
rect 21955 3772 22021 3773
rect 21955 3708 21956 3772
rect 22020 3708 22021 3772
rect 21955 3707 22021 3708
rect 21219 3228 21285 3229
rect 21219 3164 21220 3228
rect 21284 3164 21285 3228
rect 21219 3163 21285 3164
rect 20115 2684 20181 2685
rect 20115 2620 20116 2684
rect 20180 2620 20181 2684
rect 20115 2619 20181 2620
rect 22694 2549 22754 37299
rect 22691 2548 22757 2549
rect 22691 2484 22692 2548
rect 22756 2484 22757 2548
rect 22691 2483 22757 2484
rect 23246 2413 23306 56203
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 23979 55724 24045 55725
rect 23979 55660 23980 55724
rect 24044 55660 24045 55724
rect 23979 55659 24045 55660
rect 23982 5677 24042 55659
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 37227 17236 37293 17237
rect 37227 17172 37228 17236
rect 37292 17172 37293 17236
rect 37227 17171 37293 17172
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 37230 16013 37290 17171
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 37227 16012 37293 16013
rect 37227 15948 37228 16012
rect 37292 15948 37293 16012
rect 37227 15947 37293 15948
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 23979 5676 24045 5677
rect 23979 5612 23980 5676
rect 24044 5612 24045 5676
rect 23979 5611 24045 5612
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 23243 2412 23309 2413
rect 23243 2348 23244 2412
rect 23308 2348 23309 2412
rect 23243 2347 23309 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B
timestamp 1649977179
transform 1 0 9016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A0
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A0
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A0
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A0
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A0
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A0
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A0
timestamp 1649977179
transform 1 0 6808 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A0
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A0
timestamp 1649977179
transform -1 0 2024 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A0
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A0
timestamp 1649977179
transform -1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A0
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1649977179
transform 1 0 8280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1649977179
transform 1 0 5796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1649977179
transform 1 0 17664 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1649977179
transform 1 0 12420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B
timestamp 1649977179
transform -1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1649977179
transform -1 0 8004 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1649977179
transform -1 0 12144 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1649977179
transform 1 0 7544 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1649977179
transform -1 0 5060 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1649977179
transform -1 0 5888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1649977179
transform 1 0 3772 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1649977179
transform -1 0 6808 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1649977179
transform -1 0 4784 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1649977179
transform -1 0 9660 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1649977179
transform -1 0 5704 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1649977179
transform 1 0 22908 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1649977179
transform -1 0 12236 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1649977179
transform -1 0 13616 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1649977179
transform -1 0 24840 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A1
timestamp 1649977179
transform -1 0 15916 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1649977179
transform -1 0 23368 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp 1649977179
transform -1 0 17204 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1649977179
transform 1 0 26036 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1649977179
transform 1 0 15824 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1649977179
transform 1 0 24564 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1649977179
transform 1 0 13432 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1649977179
transform 1 0 15824 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1649977179
transform -1 0 14628 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1649977179
transform -1 0 14260 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C1
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1649977179
transform 1 0 13248 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1649977179
transform 1 0 13800 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__C1
timestamp 1649977179
transform 1 0 14352 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1649977179
transform -1 0 20240 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1649977179
transform -1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1649977179
transform 1 0 28888 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1649977179
transform -1 0 32016 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1649977179
transform 1 0 29440 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1649977179
transform 1 0 27784 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__C1
timestamp 1649977179
transform -1 0 28152 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1649977179
transform 1 0 27508 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__C1
timestamp 1649977179
transform 1 0 27048 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1649977179
transform 1 0 26680 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__C1
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1649977179
transform 1 0 30084 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1649977179
transform 1 0 29532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform 1 0 29716 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1
timestamp 1649977179
transform 1 0 35788 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp 1649977179
transform -1 0 37444 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1
timestamp 1649977179
transform 1 0 35236 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1649977179
transform 1 0 36616 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A1
timestamp 1649977179
transform -1 0 37444 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1649977179
transform 1 0 33672 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1649977179
transform 1 0 31464 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B
timestamp 1649977179
transform -1 0 17940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1649977179
transform -1 0 29072 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1649977179
transform 1 0 31464 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1649977179
transform 1 0 31188 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1649977179
transform -1 0 30544 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1
timestamp 1649977179
transform 1 0 26312 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1649977179
transform 1 0 27324 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A1
timestamp 1649977179
transform -1 0 30452 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A1
timestamp 1649977179
transform 1 0 29992 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A1
timestamp 1649977179
transform 1 0 33488 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1649977179
transform 1 0 31464 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1649977179
transform 1 0 32936 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A1
timestamp 1649977179
transform 1 0 33764 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A1
timestamp 1649977179
transform 1 0 34684 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A1
timestamp 1649977179
transform 1 0 34040 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A1
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1649977179
transform 1 0 29440 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1649977179
transform -1 0 30452 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C1
timestamp 1649977179
transform 1 0 29716 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1649977179
transform 1 0 10856 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1649977179
transform -1 0 10212 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1649977179
transform 1 0 16560 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1649977179
transform 1 0 5152 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__C1
timestamp 1649977179
transform 1 0 5704 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A1
timestamp 1649977179
transform -1 0 2208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__C1
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1649977179
transform 1 0 5428 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C1
timestamp 1649977179
transform -1 0 5060 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1649977179
transform 1 0 8188 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__C1
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1649977179
transform -1 0 23000 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1649977179
transform -1 0 18032 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1649977179
transform 1 0 7820 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__C1
timestamp 1649977179
transform 1 0 8096 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__C1
timestamp 1649977179
transform 1 0 19780 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__C1
timestamp 1649977179
transform -1 0 18768 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1649977179
transform 1 0 20148 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__C1
timestamp 1649977179
transform 1 0 17756 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1649977179
transform 1 0 20792 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__C1
timestamp 1649977179
transform -1 0 19872 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1649977179
transform 1 0 19504 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A1
timestamp 1649977179
transform 1 0 19136 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1649977179
transform 1 0 15824 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1649977179
transform 1 0 17204 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B
timestamp 1649977179
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1649977179
transform -1 0 15548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1649977179
transform 1 0 8924 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1649977179
transform 1 0 9016 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1649977179
transform 1 0 22724 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1649977179
transform 1 0 11592 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1649977179
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A1
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__C1
timestamp 1649977179
transform 1 0 13064 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1649977179
transform 1 0 13616 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__C1
timestamp 1649977179
transform -1 0 15180 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A1
timestamp 1649977179
transform 1 0 23920 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__C1
timestamp 1649977179
transform -1 0 23920 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1649977179
transform 1 0 23736 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__C1
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1649977179
transform 1 0 23736 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A1
timestamp 1649977179
transform 1 0 23736 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A1
timestamp 1649977179
transform 1 0 25760 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1649977179
transform 1 0 24656 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1649977179
transform 1 0 23736 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A1
timestamp 1649977179
transform 1 0 23736 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1649977179
transform -1 0 21988 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1649977179
transform -1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1649977179
transform -1 0 23368 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1649977179
transform -1 0 24840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A1
timestamp 1649977179
transform -1 0 24288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A1
timestamp 1649977179
transform 1 0 23368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1649977179
transform 1 0 18032 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1
timestamp 1649977179
transform -1 0 25024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A
timestamp 1649977179
transform -1 0 19412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A1
timestamp 1649977179
transform -1 0 25208 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1649977179
transform 1 0 28336 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1649977179
transform -1 0 33764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A1
timestamp 1649977179
transform -1 0 29716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1649977179
transform -1 0 31464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1649977179
transform 1 0 31924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform 1 0 28888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1649977179
transform 1 0 30544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1649977179
transform -1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A1
timestamp 1649977179
transform -1 0 33396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1649977179
transform 1 0 27140 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A1
timestamp 1649977179
transform -1 0 30636 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1649977179
transform 1 0 22448 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A1
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B
timestamp 1649977179
transform 1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1649977179
transform 1 0 18768 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A1
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A1
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A1
timestamp 1649977179
transform -1 0 18216 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__C1
timestamp 1649977179
transform -1 0 18768 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A1
timestamp 1649977179
transform 1 0 19320 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__C1
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1
timestamp 1649977179
transform -1 0 28704 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__C1
timestamp 1649977179
transform 1 0 28704 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A1
timestamp 1649977179
transform -1 0 31188 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__C1
timestamp 1649977179
transform -1 0 29900 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1
timestamp 1649977179
transform 1 0 31464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__C1
timestamp 1649977179
transform 1 0 30176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A1
timestamp 1649977179
transform -1 0 27508 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__C1
timestamp 1649977179
transform 1 0 28980 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__C1
timestamp 1649977179
transform 1 0 26312 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1649977179
transform -1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__C1
timestamp 1649977179
transform 1 0 23000 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1649977179
transform -1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__C1
timestamp 1649977179
transform 1 0 22264 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1649977179
transform 1 0 22080 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B
timestamp 1649977179
transform -1 0 25668 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1649977179
transform 1 0 35512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1649977179
transform -1 0 37352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1649977179
transform 1 0 33948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__C1
timestamp 1649977179
transform -1 0 34684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A1
timestamp 1649977179
transform -1 0 40020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__C1
timestamp 1649977179
transform 1 0 37904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A1
timestamp 1649977179
transform -1 0 36708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__C1
timestamp 1649977179
transform 1 0 35972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A1
timestamp 1649977179
transform 1 0 36616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__C1
timestamp 1649977179
transform -1 0 39836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 1649977179
transform 1 0 37536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__C1
timestamp 1649977179
transform 1 0 38088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A1
timestamp 1649977179
transform 1 0 37904 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__C1
timestamp 1649977179
transform -1 0 37536 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1649977179
transform 1 0 32752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A1
timestamp 1649977179
transform 1 0 39928 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1
timestamp 1649977179
transform -1 0 41860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1
timestamp 1649977179
transform -1 0 41584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A1
timestamp 1649977179
transform -1 0 41400 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A1
timestamp 1649977179
transform -1 0 41124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A1
timestamp 1649977179
transform 1 0 35880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A
timestamp 1649977179
transform 1 0 34960 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1
timestamp 1649977179
transform -1 0 34960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A1
timestamp 1649977179
transform 1 0 34040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A1
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1
timestamp 1649977179
transform 1 0 37260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1
timestamp 1649977179
transform 1 0 38364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1649977179
transform -1 0 37536 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A1
timestamp 1649977179
transform 1 0 39192 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__A1
timestamp 1649977179
transform 1 0 40756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A1
timestamp 1649977179
transform 1 0 37904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1649977179
transform 1 0 40388 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1649977179
transform 1 0 38272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1649977179
transform 1 0 35144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1649977179
transform -1 0 24564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B
timestamp 1649977179
transform -1 0 23000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1649977179
transform -1 0 25852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A
timestamp 1649977179
transform 1 0 26312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A1
timestamp 1649977179
transform 1 0 26312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A1
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A1
timestamp 1649977179
transform -1 0 29716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1649977179
transform 1 0 29440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1649977179
transform -1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1
timestamp 1649977179
transform 1 0 34592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A1
timestamp 1649977179
transform 1 0 33212 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1649977179
transform -1 0 23920 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A1
timestamp 1649977179
transform 1 0 32200 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A1
timestamp 1649977179
transform 1 0 32384 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A1
timestamp 1649977179
transform 1 0 31464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A1
timestamp 1649977179
transform 1 0 27140 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1649977179
transform 1 0 5612 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1649977179
transform 1 0 19044 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1649977179
transform 1 0 16008 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1649977179
transform 1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1649977179
transform 1 0 8096 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A
timestamp 1649977179
transform -1 0 16836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A
timestamp 1649977179
transform 1 0 8096 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A1
timestamp 1649977179
transform 1 0 4324 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A1
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1649977179
transform 1 0 2852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A
timestamp 1649977179
transform 1 0 6348 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A1
timestamp 1649977179
transform 1 0 5888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1649977179
transform 1 0 8464 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A1
timestamp 1649977179
transform 1 0 8096 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1649977179
transform -1 0 21896 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1649977179
transform 1 0 20700 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A
timestamp 1649977179
transform 1 0 19688 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1649977179
transform -1 0 21160 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1649977179
transform 1 0 21896 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A1
timestamp 1649977179
transform -1 0 23828 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A1
timestamp 1649977179
transform -1 0 23552 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A
timestamp 1649977179
transform 1 0 16836 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1649977179
transform 1 0 21160 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 1649977179
transform -1 0 17020 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A1
timestamp 1649977179
transform -1 0 21252 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A
timestamp 1649977179
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__B
timestamp 1649977179
transform 1 0 17756 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A
timestamp 1649977179
transform 1 0 17940 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A1
timestamp 1649977179
transform 1 0 17664 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A2
timestamp 1649977179
transform -1 0 17664 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 1649977179
transform 1 0 10120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__B
timestamp 1649977179
transform -1 0 21436 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1649977179
transform -1 0 19320 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A2
timestamp 1649977179
transform 1 0 19320 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A
timestamp 1649977179
transform -1 0 21528 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__B
timestamp 1649977179
transform 1 0 22172 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1649977179
transform -1 0 22540 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1649977179
transform -1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1649977179
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A1
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 1649977179
transform 1 0 18400 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1649977179
transform 1 0 16928 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A1
timestamp 1649977179
transform -1 0 19872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A1
timestamp 1649977179
transform -1 0 24564 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A1
timestamp 1649977179
transform -1 0 26312 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A1
timestamp 1649977179
transform -1 0 27140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1649977179
transform -1 0 13248 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A1
timestamp 1649977179
transform 1 0 24472 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__C1
timestamp 1649977179
transform -1 0 24840 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__A1
timestamp 1649977179
transform -1 0 25116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__C1
timestamp 1649977179
transform 1 0 24380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A1
timestamp 1649977179
transform 1 0 21804 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__C1
timestamp 1649977179
transform -1 0 22172 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__A1
timestamp 1649977179
transform 1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__C1
timestamp 1649977179
transform 1 0 22172 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1649977179
transform -1 0 10856 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__B
timestamp 1649977179
transform -1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 1649977179
transform -1 0 8464 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A
timestamp 1649977179
transform 1 0 12880 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A1
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__C1
timestamp 1649977179
transform 1 0 8004 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A1
timestamp 1649977179
transform -1 0 2208 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__C1
timestamp 1649977179
transform -1 0 3956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1649977179
transform 1 0 2576 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__C1
timestamp 1649977179
transform 1 0 3956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A1
timestamp 1649977179
transform 1 0 4968 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__C1
timestamp 1649977179
transform 1 0 5520 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A1
timestamp 1649977179
transform 1 0 7820 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__C1
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A1
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__C1
timestamp 1649977179
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A1
timestamp 1649977179
transform 1 0 16192 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A1
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A1
timestamp 1649977179
transform 1 0 18032 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A1
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A1
timestamp 1649977179
transform -1 0 12512 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A1
timestamp 1649977179
transform 1 0 10764 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A
timestamp 1649977179
transform -1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__B
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A
timestamp 1649977179
transform 1 0 8740 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A
timestamp 1649977179
transform 1 0 9292 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A1
timestamp 1649977179
transform 1 0 3864 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A1
timestamp 1649977179
transform -1 0 3956 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A1
timestamp 1649977179
transform 1 0 2852 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A1
timestamp 1649977179
transform 1 0 5428 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1649977179
transform -1 0 8372 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A1
timestamp 1649977179
transform -1 0 9844 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A1
timestamp 1649977179
transform 1 0 10856 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A1
timestamp 1649977179
transform -1 0 11040 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__A1
timestamp 1649977179
transform 1 0 10856 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A
timestamp 1649977179
transform 1 0 11684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A1
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__C1
timestamp 1649977179
transform 1 0 11040 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__A1
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__C1
timestamp 1649977179
transform 1 0 9936 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A1
timestamp 1649977179
transform 1 0 9936 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__C1
timestamp 1649977179
transform 1 0 10488 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A
timestamp 1649977179
transform -1 0 15088 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__B
timestamp 1649977179
transform 1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__A
timestamp 1649977179
transform -1 0 14628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A
timestamp 1649977179
transform 1 0 15732 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__A1
timestamp 1649977179
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__C1
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A1
timestamp 1649977179
transform 1 0 9292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__C1
timestamp 1649977179
transform -1 0 12512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A
timestamp 1649977179
transform 1 0 14260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__A1
timestamp 1649977179
transform -1 0 11776 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A1
timestamp 1649977179
transform -1 0 13340 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A1
timestamp 1649977179
transform 1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A1
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__A1
timestamp 1649977179
transform -1 0 20148 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__A
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A1
timestamp 1649977179
transform -1 0 20516 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__A1
timestamp 1649977179
transform 1 0 21160 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A1
timestamp 1649977179
transform 1 0 16928 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A1
timestamp 1649977179
transform 1 0 17848 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A1
timestamp 1649977179
transform 1 0 18216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__A
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__A
timestamp 1649977179
transform 1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__A
timestamp 1649977179
transform -1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__A
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A1
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A1
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__A1
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A1
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A1
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__A
timestamp 1649977179
transform -1 0 25576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__A1
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__A1
timestamp 1649977179
transform 1 0 29624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A1
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A1
timestamp 1649977179
transform 1 0 26312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__A1
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__A1
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__C1
timestamp 1649977179
transform 1 0 16744 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A1
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__C1
timestamp 1649977179
transform -1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__D
timestamp 1649977179
transform -1 0 25116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__C1
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__D
timestamp 1649977179
transform -1 0 25024 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1551__A
timestamp 1649977179
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__C1
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__A
timestamp 1649977179
transform 1 0 24104 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__D
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__C1
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__A
timestamp 1649977179
transform 1 0 30452 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__A
timestamp 1649977179
transform -1 0 32292 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__A2
timestamp 1649977179
transform -1 0 14996 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__B1
timestamp 1649977179
transform -1 0 14996 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__A
timestamp 1649977179
transform -1 0 8648 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1604__A1
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__A2
timestamp 1649977179
transform -1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__B1
timestamp 1649977179
transform 1 0 15272 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__A
timestamp 1649977179
transform -1 0 9936 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__A2
timestamp 1649977179
transform -1 0 24564 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__B1
timestamp 1649977179
transform -1 0 23828 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1633__B1
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__A2
timestamp 1649977179
transform 1 0 23092 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__B1
timestamp 1649977179
transform 1 0 23460 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1646__B1
timestamp 1649977179
transform -1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__A2
timestamp 1649977179
transform -1 0 23552 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__B1
timestamp 1649977179
transform 1 0 22172 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1671__B1
timestamp 1649977179
transform -1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__B1
timestamp 1649977179
transform -1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1707__B1
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1708__A
timestamp 1649977179
transform -1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2167__A
timestamp 1649977179
transform 1 0 42688 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2168__A
timestamp 1649977179
transform -1 0 45172 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2169__A
timestamp 1649977179
transform 1 0 43976 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2170__A
timestamp 1649977179
transform 1 0 21896 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2171__A
timestamp 1649977179
transform -1 0 20424 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2172__A
timestamp 1649977179
transform -1 0 29716 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2173__A
timestamp 1649977179
transform 1 0 43332 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2174__A
timestamp 1649977179
transform 1 0 45908 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2175__A
timestamp 1649977179
transform -1 0 45448 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2176__A
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2177__A
timestamp 1649977179
transform 1 0 15088 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2178__A
timestamp 1649977179
transform -1 0 16192 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2179__A
timestamp 1649977179
transform 1 0 16468 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2180__A
timestamp 1649977179
transform 1 0 17112 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2181__A
timestamp 1649977179
transform 1 0 18400 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2182__A
timestamp 1649977179
transform -1 0 20608 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2183__A
timestamp 1649977179
transform -1 0 23920 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2184__A
timestamp 1649977179
transform 1 0 17756 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2185__A
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2186__A
timestamp 1649977179
transform 1 0 27048 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2187__A
timestamp 1649977179
transform -1 0 28244 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2188__A
timestamp 1649977179
transform 1 0 29992 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2189__A
timestamp 1649977179
transform -1 0 32936 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2190__A
timestamp 1649977179
transform -1 0 34408 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2191__A
timestamp 1649977179
transform 1 0 30820 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2192__A
timestamp 1649977179
transform -1 0 36616 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2193__A
timestamp 1649977179
transform -1 0 28428 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2194__A
timestamp 1649977179
transform 1 0 46552 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2195__A
timestamp 1649977179
transform -1 0 43976 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2196__A
timestamp 1649977179
transform -1 0 57132 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 20608 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_wb_clk_i_A
timestamp 1649977179
transform -1 0 12420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 12604 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 27232 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1649977179
transform -1 0 16008 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1649977179
transform 1 0 6716 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1649977179
transform 1 0 7084 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1649977179
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1649977179
transform 1 0 17388 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1649977179
transform 1 0 16376 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1649977179
transform 1 0 23276 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1649977179
transform 1 0 29716 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1649977179
transform 1 0 25944 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1649977179
transform -1 0 29900 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1649977179
transform 1 0 32292 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1649977179
transform 1 0 38180 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1649977179
transform 1 0 31464 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1649977179
transform 1 0 28612 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1649977179
transform 1 0 30544 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1649977179
transform -1 0 37536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1649977179
transform 1 0 36616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1649977179
transform 1 0 37352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1649977179
transform -1 0 32384 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_wb_clk_i_A
timestamp 1649977179
transform 1 0 27048 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_wb_clk_i_A
timestamp 1649977179
transform 1 0 28152 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_wb_clk_i_A
timestamp 1649977179
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_28_wb_clk_i_A
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_29_wb_clk_i_A
timestamp 1649977179
transform 1 0 16836 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_30_wb_clk_i_A
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_31_wb_clk_i_A
timestamp 1649977179
transform -1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_32_wb_clk_i_A
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_33_wb_clk_i_A
timestamp 1649977179
transform -1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 11316 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 12972 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 17664 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 23368 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 25668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 21344 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 19504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 20332 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 20884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 20792 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 22264 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 21712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 22816 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 23460 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 25116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 22632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 14996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 14444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 12972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 24012 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 11868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 13892 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 6900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 6072 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 9016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 6992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 1564 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 4968 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 1656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 2024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 5520 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 1840 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 3312 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1649977179
transform 1 0 40756 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1649977179
transform 1 0 42320 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform 1 0 56028 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36
timestamp 1649977179
transform 1 0 4416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9476 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1649977179
transform 1 0 17296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_184
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1649977179
transform 1 0 19872 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1649977179
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1649977179
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_255
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_283
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1649977179
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_323
timestamp 1649977179
transform 1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1649977179
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_340
timestamp 1649977179
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1649977179
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1649977179
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10
timestamp 1649977179
transform 1 0 2024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_38
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_43
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1649977179
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1649977179
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_212
timestamp 1649977179
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1649977179
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1649977179
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_244
timestamp 1649977179
transform 1 0 23552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1649977179
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_303
timestamp 1649977179
transform 1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1649977179
transform 1 0 29624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_324 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_340
timestamp 1649977179
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_354
timestamp 1649977179
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1649977179
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1649977179
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1649977179
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1649977179
transform 1 0 58512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_89
timestamp 1649977179
transform 1 0 9292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp 1649977179
transform 1 0 11960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1649977179
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_183
timestamp 1649977179
transform 1 0 17940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1649977179
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1649977179
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_214
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_223
timestamp 1649977179
transform 1 0 21620 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1649977179
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1649977179
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1649977179
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_257
timestamp 1649977179
transform 1 0 24748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_261
timestamp 1649977179
transform 1 0 25116 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_270
timestamp 1649977179
transform 1 0 25944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_278
timestamp 1649977179
transform 1 0 26680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_282
timestamp 1649977179
transform 1 0 27048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_291
timestamp 1649977179
transform 1 0 27876 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_299
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1649977179
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_340
timestamp 1649977179
transform 1 0 32384 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_352
timestamp 1649977179
transform 1 0 33488 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1649977179
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_376
timestamp 1649977179
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1649977179
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_390
timestamp 1649977179
transform 1 0 36984 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_399
timestamp 1649977179
transform 1 0 37812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_407
timestamp 1649977179
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1649977179
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1649977179
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_440
timestamp 1649977179
transform 1 0 41584 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_448
timestamp 1649977179
transform 1 0 42320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1649977179
transform 1 0 42780 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_460
timestamp 1649977179
transform 1 0 43424 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1649977179
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1649977179
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1649977179
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1649977179
transform 1 0 46552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_510
timestamp 1649977179
transform 1 0 48024 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_517
timestamp 1649977179
transform 1 0 48668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_529
timestamp 1649977179
transform 1 0 49772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_537
timestamp 1649977179
transform 1 0 50508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_544
timestamp 1649977179
transform 1 0 51152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_551
timestamp 1649977179
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_558
timestamp 1649977179
transform 1 0 52440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1649977179
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_610
timestamp 1649977179
transform 1 0 57224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_614
timestamp 1649977179
transform 1 0 57592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1649977179
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1649977179
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_19
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_43
timestamp 1649977179
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_63
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_84
timestamp 1649977179
transform 1 0 8832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_92
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_96
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1649977179
transform 1 0 12420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1649977179
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_196
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1649977179
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1649977179
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1649977179
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_246
timestamp 1649977179
transform 1 0 23736 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_255
timestamp 1649977179
transform 1 0 24564 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_267
timestamp 1649977179
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_297
timestamp 1649977179
transform 1 0 28428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_309
timestamp 1649977179
transform 1 0 29532 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_321
timestamp 1649977179
transform 1 0 30636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp 1649977179
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_380
timestamp 1649977179
transform 1 0 36064 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_547
timestamp 1649977179
transform 1 0 51428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_554
timestamp 1649977179
transform 1 0 52072 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_564
timestamp 1649977179
transform 1 0 52992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1649977179
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_578
timestamp 1649977179
transform 1 0 54280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_592
timestamp 1649977179
transform 1 0 55568 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_599
timestamp 1649977179
transform 1 0 56212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_611
timestamp 1649977179
transform 1 0 57316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1649977179
transform 1 0 58236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_8
timestamp 1649977179
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_14
timestamp 1649977179
transform 1 0 2392 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1649977179
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_57
timestamp 1649977179
transform 1 0 6348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_92
timestamp 1649977179
transform 1 0 9568 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_107
timestamp 1649977179
transform 1 0 10948 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_111
timestamp 1649977179
transform 1 0 11316 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1649977179
transform 1 0 11684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_122
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_143
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_150
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1649977179
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1649977179
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1649977179
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1649977179
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_269
timestamp 1649977179
transform 1 0 25852 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_281
timestamp 1649977179
transform 1 0 26956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_293
timestamp 1649977179
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 1649977179
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_341
timestamp 1649977179
transform 1 0 32476 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_353
timestamp 1649977179
transform 1 0 33580 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 1649977179
transform 1 0 34316 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_553
timestamp 1649977179
transform 1 0 51980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_558
timestamp 1649977179
transform 1 0 52440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_565
timestamp 1649977179
transform 1 0 53084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_572
timestamp 1649977179
transform 1 0 53728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_579
timestamp 1649977179
transform 1 0 54372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_592
timestamp 1649977179
transform 1 0 55568 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_599
timestamp 1649977179
transform 1 0 56212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_611
timestamp 1649977179
transform 1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1649977179
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_10
timestamp 1649977179
transform 1 0 2024 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_23
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_62
timestamp 1649977179
transform 1 0 6808 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_80
timestamp 1649977179
transform 1 0 8464 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_87
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1649977179
transform 1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1649977179
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_121
timestamp 1649977179
transform 1 0 12236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_142
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1649977179
transform 1 0 15180 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_174
timestamp 1649977179
transform 1 0 17112 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_182
timestamp 1649977179
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_194
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_203
timestamp 1649977179
transform 1 0 19780 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_210
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1649977179
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_228
timestamp 1649977179
transform 1 0 22080 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1649977179
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_266
timestamp 1649977179
transform 1 0 25576 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1649977179
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_289
timestamp 1649977179
transform 1 0 27692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_301
timestamp 1649977179
transform 1 0 28796 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_309
timestamp 1649977179
transform 1 0 29532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_312
timestamp 1649977179
transform 1 0 29808 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_324
timestamp 1649977179
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_340
timestamp 1649977179
transform 1 0 32384 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_352
timestamp 1649977179
transform 1 0 33488 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_364
timestamp 1649977179
transform 1 0 34592 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_376
timestamp 1649977179
transform 1 0 35696 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1649977179
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_409
timestamp 1649977179
transform 1 0 38732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_421
timestamp 1649977179
transform 1 0 39836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_433
timestamp 1649977179
transform 1 0 40940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1649977179
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_569
timestamp 1649977179
transform 1 0 53452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_575
timestamp 1649977179
transform 1 0 54004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_582
timestamp 1649977179
transform 1 0 54648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_589
timestamp 1649977179
transform 1 0 55292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_601
timestamp 1649977179
transform 1 0 56396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_613
timestamp 1649977179
transform 1 0 57500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1649977179
transform 1 0 58236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_39
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_50
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1649977179
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_64
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_95
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_104
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_111
timestamp 1649977179
transform 1 0 11316 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_118
timestamp 1649977179
transform 1 0 11960 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_127
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_179
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_183
timestamp 1649977179
transform 1 0 17940 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_224
timestamp 1649977179
transform 1 0 21712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1649977179
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_236
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_242
timestamp 1649977179
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1649977179
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_258
timestamp 1649977179
transform 1 0 24840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_276
timestamp 1649977179
transform 1 0 26496 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_284
timestamp 1649977179
transform 1 0 27232 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_290
timestamp 1649977179
transform 1 0 27784 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1649977179
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_311
timestamp 1649977179
transform 1 0 29716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1649977179
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_332
timestamp 1649977179
transform 1 0 31648 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_360
timestamp 1649977179
transform 1 0 34224 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_373
timestamp 1649977179
transform 1 0 35420 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_384
timestamp 1649977179
transform 1 0 36432 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_396
timestamp 1649977179
transform 1 0 37536 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_408
timestamp 1649977179
transform 1 0 38640 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_13
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_19
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_64
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_68
timestamp 1649977179
transform 1 0 7360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_82
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_86
timestamp 1649977179
transform 1 0 9016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1649977179
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1649977179
transform 1 0 12420 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_135
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_155
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_206
timestamp 1649977179
transform 1 0 20056 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_209
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_215
timestamp 1649977179
transform 1 0 20884 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1649977179
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_246
timestamp 1649977179
transform 1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_252
timestamp 1649977179
transform 1 0 24288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_283
timestamp 1649977179
transform 1 0 27140 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_295
timestamp 1649977179
transform 1 0 28244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_303
timestamp 1649977179
transform 1 0 28980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_307
timestamp 1649977179
transform 1 0 29348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_319
timestamp 1649977179
transform 1 0 30452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_328
timestamp 1649977179
transform 1 0 31280 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_381
timestamp 1649977179
transform 1 0 36156 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_387
timestamp 1649977179
transform 1 0 36708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_401
timestamp 1649977179
transform 1 0 37996 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_420
timestamp 1649977179
transform 1 0 39744 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_432
timestamp 1649977179
transform 1 0 40848 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_444
timestamp 1649977179
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1649977179
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_16
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_50
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_8_61
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1649977179
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_111
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_131
timestamp 1649977179
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_145
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_151
timestamp 1649977179
transform 1 0 14996 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_173
timestamp 1649977179
transform 1 0 17020 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_200
timestamp 1649977179
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_214
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_220
timestamp 1649977179
transform 1 0 21344 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_236
timestamp 1649977179
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_261
timestamp 1649977179
transform 1 0 25116 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_267
timestamp 1649977179
transform 1 0 25668 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_278
timestamp 1649977179
transform 1 0 26680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_284
timestamp 1649977179
transform 1 0 27232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_304
timestamp 1649977179
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_313
timestamp 1649977179
transform 1 0 29900 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_330
timestamp 1649977179
transform 1 0 31464 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_342
timestamp 1649977179
transform 1 0 32568 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_354
timestamp 1649977179
transform 1 0 33672 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1649977179
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_373
timestamp 1649977179
transform 1 0 35420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_385
timestamp 1649977179
transform 1 0 36524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_394
timestamp 1649977179
transform 1 0 37352 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_402
timestamp 1649977179
transform 1 0 38088 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_414
timestamp 1649977179
transform 1 0 39192 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_423
timestamp 1649977179
transform 1 0 40020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_435
timestamp 1649977179
transform 1 0 41124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_447
timestamp 1649977179
transform 1 0 42228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_459
timestamp 1649977179
transform 1 0 43332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_471
timestamp 1649977179
transform 1 0 44436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_8
timestamp 1649977179
transform 1 0 1840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_14
timestamp 1649977179
transform 1 0 2392 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_20
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_26
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_32
timestamp 1649977179
transform 1 0 4048 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_68
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_102
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1649977179
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_124
timestamp 1649977179
transform 1 0 12512 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_130
timestamp 1649977179
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_133
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_145
timestamp 1649977179
transform 1 0 14444 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_155
timestamp 1649977179
transform 1 0 15364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1649977179
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_180
timestamp 1649977179
transform 1 0 17664 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_194
timestamp 1649977179
transform 1 0 18952 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_201
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_238
timestamp 1649977179
transform 1 0 23000 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1649977179
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_253
timestamp 1649977179
transform 1 0 24380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_257
timestamp 1649977179
transform 1 0 24748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_260
timestamp 1649977179
transform 1 0 25024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1649977179
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_284
timestamp 1649977179
transform 1 0 27232 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_292
timestamp 1649977179
transform 1 0 27968 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_298
timestamp 1649977179
transform 1 0 28520 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_310
timestamp 1649977179
transform 1 0 29624 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_323
timestamp 1649977179
transform 1 0 30820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_357
timestamp 1649977179
transform 1 0 33948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_363
timestamp 1649977179
transform 1 0 34500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_375
timestamp 1649977179
transform 1 0 35604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_386
timestamp 1649977179
transform 1 0 36616 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_413
timestamp 1649977179
transform 1 0 39100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_425
timestamp 1649977179
transform 1 0 40204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_437
timestamp 1649977179
transform 1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1649977179
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_6
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_12
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_18
timestamp 1649977179
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_42
timestamp 1649977179
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_48
timestamp 1649977179
transform 1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_54
timestamp 1649977179
transform 1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_74
timestamp 1649977179
transform 1 0 7912 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_93
timestamp 1649977179
transform 1 0 9660 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_128
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_132
timestamp 1649977179
transform 1 0 13248 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_149
timestamp 1649977179
transform 1 0 14812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_173
timestamp 1649977179
transform 1 0 17020 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_179
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_182
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_188
timestamp 1649977179
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_202
timestamp 1649977179
transform 1 0 19688 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_214
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_225
timestamp 1649977179
transform 1 0 21804 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_241
timestamp 1649977179
transform 1 0 23276 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_249
timestamp 1649977179
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_258
timestamp 1649977179
transform 1 0 24840 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_266
timestamp 1649977179
transform 1 0 25576 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_283
timestamp 1649977179
transform 1 0 27140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_295
timestamp 1649977179
transform 1 0 28244 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_315
timestamp 1649977179
transform 1 0 30084 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_332
timestamp 1649977179
transform 1 0 31648 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_344
timestamp 1649977179
transform 1 0 32752 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_356
timestamp 1649977179
transform 1 0 33856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_375
timestamp 1649977179
transform 1 0 35604 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_381
timestamp 1649977179
transform 1 0 36156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1649977179
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_399
timestamp 1649977179
transform 1 0 37812 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1649977179
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_617
timestamp 1649977179
transform 1 0 57868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1649977179
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_5
timestamp 1649977179
transform 1 0 1564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_11
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_31
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_92
timestamp 1649977179
transform 1 0 9568 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_154
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1649977179
transform 1 0 16928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1649977179
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_303
timestamp 1649977179
transform 1 0 28980 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_327
timestamp 1649977179
transform 1 0 31188 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_339
timestamp 1649977179
transform 1 0 32292 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_351
timestamp 1649977179
transform 1 0 33396 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_363
timestamp 1649977179
transform 1 0 34500 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_368
timestamp 1649977179
transform 1 0 34960 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_380
timestamp 1649977179
transform 1 0 36064 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1649977179
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1649977179
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_415
timestamp 1649977179
transform 1 0 39284 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_421
timestamp 1649977179
transform 1 0 39836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_433
timestamp 1649977179
transform 1 0 40940 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_445
timestamp 1649977179
transform 1 0 42044 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_10
timestamp 1649977179
transform 1 0 2024 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1649977179
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_35
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_48
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_55
timestamp 1649977179
transform 1 0 6164 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_68
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_74
timestamp 1649977179
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1649977179
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_118
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_130
timestamp 1649977179
transform 1 0 13064 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_164
timestamp 1649977179
transform 1 0 16192 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_170
timestamp 1649977179
transform 1 0 16744 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_213
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_220
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_236
timestamp 1649977179
transform 1 0 22816 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_248
timestamp 1649977179
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_255
timestamp 1649977179
transform 1 0 24564 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_267
timestamp 1649977179
transform 1 0 25668 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_279
timestamp 1649977179
transform 1 0 26772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_290
timestamp 1649977179
transform 1 0 27784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_316
timestamp 1649977179
transform 1 0 30176 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_344
timestamp 1649977179
transform 1 0 32752 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_356
timestamp 1649977179
transform 1 0 33856 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_376
timestamp 1649977179
transform 1 0 35696 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_384
timestamp 1649977179
transform 1 0 36432 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_392
timestamp 1649977179
transform 1 0 37168 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_416
timestamp 1649977179
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_617
timestamp 1649977179
transform 1 0 57868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1649977179
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_6
timestamp 1649977179
transform 1 0 1656 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_26
timestamp 1649977179
transform 1 0 3496 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_38
timestamp 1649977179
transform 1 0 4600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_65
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_71
timestamp 1649977179
transform 1 0 7636 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_84
timestamp 1649977179
transform 1 0 8832 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_116
timestamp 1649977179
transform 1 0 11776 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_120
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_123
timestamp 1649977179
transform 1 0 12420 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_144
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_194
timestamp 1649977179
transform 1 0 18952 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_206
timestamp 1649977179
transform 1 0 20056 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_212
timestamp 1649977179
transform 1 0 20608 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_235
timestamp 1649977179
transform 1 0 22724 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_246
timestamp 1649977179
transform 1 0 23736 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_258
timestamp 1649977179
transform 1 0 24840 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1649977179
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1649977179
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_314
timestamp 1649977179
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_318
timestamp 1649977179
transform 1 0 30360 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_321
timestamp 1649977179
transform 1 0 30636 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1649977179
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_345
timestamp 1649977179
transform 1 0 32844 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_351
timestamp 1649977179
transform 1 0 33396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_363
timestamp 1649977179
transform 1 0 34500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_367
timestamp 1649977179
transform 1 0 34868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_384
timestamp 1649977179
transform 1 0 36432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_396
timestamp 1649977179
transform 1 0 37536 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_404
timestamp 1649977179
transform 1 0 38272 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_421
timestamp 1649977179
transform 1 0 39836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_433
timestamp 1649977179
transform 1 0 40940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1649977179
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_16
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_35
timestamp 1649977179
transform 1 0 4324 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_40
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_52
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_63
timestamp 1649977179
transform 1 0 6900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1649977179
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_145
timestamp 1649977179
transform 1 0 14444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_151
timestamp 1649977179
transform 1 0 14996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_167
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_173
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_185
timestamp 1649977179
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1649977179
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_259
timestamp 1649977179
transform 1 0 24932 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_262
timestamp 1649977179
transform 1 0 25208 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_266
timestamp 1649977179
transform 1 0 25576 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_272
timestamp 1649977179
transform 1 0 26128 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_284
timestamp 1649977179
transform 1 0 27232 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_296
timestamp 1649977179
transform 1 0 28336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_319
timestamp 1649977179
transform 1 0 30452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_331
timestamp 1649977179
transform 1 0 31556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_337
timestamp 1649977179
transform 1 0 32108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_371
timestamp 1649977179
transform 1 0 35236 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_410
timestamp 1649977179
transform 1 0 38824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_418
timestamp 1649977179
transform 1 0 39560 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_67
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_79
timestamp 1649977179
transform 1 0 8372 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_91
timestamp 1649977179
transform 1 0 9476 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_115
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_127
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_139
timestamp 1649977179
transform 1 0 13892 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_151
timestamp 1649977179
transform 1 0 14996 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_199
timestamp 1649977179
transform 1 0 19412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_211
timestamp 1649977179
transform 1 0 20516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 1649977179
transform 1 0 22172 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_235
timestamp 1649977179
transform 1 0 22724 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_239
timestamp 1649977179
transform 1 0 23092 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_242
timestamp 1649977179
transform 1 0 23368 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_250
timestamp 1649977179
transform 1 0 24104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_258
timestamp 1649977179
transform 1 0 24840 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_270
timestamp 1649977179
transform 1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_278
timestamp 1649977179
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_284
timestamp 1649977179
transform 1 0 27232 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1649977179
transform 1 0 28244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_319
timestamp 1649977179
transform 1 0 30452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1649977179
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_359
timestamp 1649977179
transform 1 0 34132 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_365
timestamp 1649977179
transform 1 0 34684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_377
timestamp 1649977179
transform 1 0 35788 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_386
timestamp 1649977179
transform 1 0 36616 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_425
timestamp 1649977179
transform 1 0 40204 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_437
timestamp 1649977179
transform 1 0 41308 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_445
timestamp 1649977179
transform 1 0 42044 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1649977179
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1649977179
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_87
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_99
timestamp 1649977179
transform 1 0 10212 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_115
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_186
timestamp 1649977179
transform 1 0 18216 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_200
timestamp 1649977179
transform 1 0 19504 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_208
timestamp 1649977179
transform 1 0 20240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_212
timestamp 1649977179
transform 1 0 20608 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_220
timestamp 1649977179
transform 1 0 21344 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_238
timestamp 1649977179
transform 1 0 23000 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_247
timestamp 1649977179
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_264
timestamp 1649977179
transform 1 0 25392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_286
timestamp 1649977179
transform 1 0 27416 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_294
timestamp 1649977179
transform 1 0 28152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_299
timestamp 1649977179
transform 1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_315
timestamp 1649977179
transform 1 0 30084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_332
timestamp 1649977179
transform 1 0 31648 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_346
timestamp 1649977179
transform 1 0 32936 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1649977179
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_383
timestamp 1649977179
transform 1 0 36340 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_395
timestamp 1649977179
transform 1 0 37444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_398
timestamp 1649977179
transform 1 0 37720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_404
timestamp 1649977179
transform 1 0 38272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1649977179
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_426
timestamp 1649977179
transform 1 0 40296 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_438
timestamp 1649977179
transform 1 0 41400 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_450
timestamp 1649977179
transform 1 0 42504 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_462
timestamp 1649977179
transform 1 0 43608 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_474
timestamp 1649977179
transform 1 0 44712 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_22
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_40
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_66
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_100
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_197
timestamp 1649977179
transform 1 0 19228 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_236
timestamp 1649977179
transform 1 0 22816 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_243
timestamp 1649977179
transform 1 0 23460 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_257
timestamp 1649977179
transform 1 0 24748 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1649977179
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_299
timestamp 1649977179
transform 1 0 28612 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_307
timestamp 1649977179
transform 1 0 29348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_311
timestamp 1649977179
transform 1 0 29716 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_323
timestamp 1649977179
transform 1 0 30820 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_342
timestamp 1649977179
transform 1 0 32568 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_354
timestamp 1649977179
transform 1 0 33672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_366
timestamp 1649977179
transform 1 0 34776 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_377
timestamp 1649977179
transform 1 0 35788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_389
timestamp 1649977179
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_397
timestamp 1649977179
transform 1 0 37628 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_408
timestamp 1649977179
transform 1 0 38640 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_414
timestamp 1649977179
transform 1 0 39192 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_419
timestamp 1649977179
transform 1 0 39652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_431
timestamp 1649977179
transform 1 0 40756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_443
timestamp 1649977179
transform 1 0 41860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1649977179
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1649977179
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1649977179
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_58
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_64
timestamp 1649977179
transform 1 0 6992 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_79
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_127
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_173
timestamp 1649977179
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_179
timestamp 1649977179
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1649977179
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_199
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1649977179
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_228
timestamp 1649977179
transform 1 0 22080 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1649977179
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_240
timestamp 1649977179
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1649977179
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_267
timestamp 1649977179
transform 1 0 25668 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_279
timestamp 1649977179
transform 1 0 26772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_285
timestamp 1649977179
transform 1 0 27324 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_290
timestamp 1649977179
transform 1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_298
timestamp 1649977179
transform 1 0 28520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_306
timestamp 1649977179
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_317
timestamp 1649977179
transform 1 0 30268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_322
timestamp 1649977179
transform 1 0 30728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_334
timestamp 1649977179
transform 1 0 31832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_354
timestamp 1649977179
transform 1 0 33672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1649977179
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_380
timestamp 1649977179
transform 1 0 36064 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_404
timestamp 1649977179
transform 1 0 38272 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_416
timestamp 1649977179
transform 1 0 39376 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1649977179
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1649977179
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1649977179
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_9
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_33
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_59
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_63
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_88
timestamp 1649977179
transform 1 0 9200 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1649977179
transform 1 0 10120 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_138
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_186
timestamp 1649977179
transform 1 0 18216 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_198
timestamp 1649977179
transform 1 0 19320 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_206
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_227
timestamp 1649977179
transform 1 0 21988 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_235
timestamp 1649977179
transform 1 0 22724 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_238
timestamp 1649977179
transform 1 0 23000 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_246
timestamp 1649977179
transform 1 0 23736 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_252
timestamp 1649977179
transform 1 0 24288 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_258
timestamp 1649977179
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_270
timestamp 1649977179
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1649977179
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_283
timestamp 1649977179
transform 1 0 27140 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_295
timestamp 1649977179
transform 1 0 28244 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_307
timestamp 1649977179
transform 1 0 29348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_319
timestamp 1649977179
transform 1 0 30452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_331
timestamp 1649977179
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_344
timestamp 1649977179
transform 1 0 32752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_358
timestamp 1649977179
transform 1 0 34040 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_366
timestamp 1649977179
transform 1 0 34776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_370
timestamp 1649977179
transform 1 0 35144 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_376
timestamp 1649977179
transform 1 0 35696 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1649977179
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_398
timestamp 1649977179
transform 1 0 37720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_406
timestamp 1649977179
transform 1 0 38456 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_424
timestamp 1649977179
transform 1 0 40112 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_436
timestamp 1649977179
transform 1 0 41216 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_16
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_37
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1649977179
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_59
timestamp 1649977179
transform 1 0 6532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_95
timestamp 1649977179
transform 1 0 9844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_107
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_115
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_120
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_159
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_171
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_183
timestamp 1649977179
transform 1 0 17940 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_199
timestamp 1649977179
transform 1 0 19412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_207
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_227
timestamp 1649977179
transform 1 0 21988 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_230
timestamp 1649977179
transform 1 0 22264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1649977179
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_281
timestamp 1649977179
transform 1 0 26956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_290
timestamp 1649977179
transform 1 0 27784 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_296
timestamp 1649977179
transform 1 0 28336 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_325
timestamp 1649977179
transform 1 0 31004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_337
timestamp 1649977179
transform 1 0 32108 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_349
timestamp 1649977179
transform 1 0 33212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_355
timestamp 1649977179
transform 1 0 33764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_369
timestamp 1649977179
transform 1 0 35052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_380
timestamp 1649977179
transform 1 0 36064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_384
timestamp 1649977179
transform 1 0 36432 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_388
timestamp 1649977179
transform 1 0 36800 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_394
timestamp 1649977179
transform 1 0 37352 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_398
timestamp 1649977179
transform 1 0 37720 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_404
timestamp 1649977179
transform 1 0 38272 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_416
timestamp 1649977179
transform 1 0 39376 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1649977179
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1649977179
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_617
timestamp 1649977179
transform 1 0 57868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1649977179
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_65
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_77
timestamp 1649977179
transform 1 0 8188 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_82
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_94
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_148
timestamp 1649977179
transform 1 0 14720 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_160
timestamp 1649977179
transform 1 0 15824 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1649977179
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_200
timestamp 1649977179
transform 1 0 19504 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_209
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_216
timestamp 1649977179
transform 1 0 20976 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_231
timestamp 1649977179
transform 1 0 22356 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_244
timestamp 1649977179
transform 1 0 23552 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1649977179
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_260
timestamp 1649977179
transform 1 0 25024 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_272
timestamp 1649977179
transform 1 0 26128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_292
timestamp 1649977179
transform 1 0 27968 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_298
timestamp 1649977179
transform 1 0 28520 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_304
timestamp 1649977179
transform 1 0 29072 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_316
timestamp 1649977179
transform 1 0 30176 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_324
timestamp 1649977179
transform 1 0 30912 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1649977179
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_366
timestamp 1649977179
transform 1 0 34776 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_375
timestamp 1649977179
transform 1 0 35604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_379
timestamp 1649977179
transform 1 0 35972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1649977179
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_415
timestamp 1649977179
transform 1 0 39284 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_423
timestamp 1649977179
transform 1 0 40020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_435
timestamp 1649977179
transform 1 0 41124 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_32
timestamp 1649977179
transform 1 0 4048 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_44
timestamp 1649977179
transform 1 0 5152 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_70
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_98
timestamp 1649977179
transform 1 0 10120 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_110
timestamp 1649977179
transform 1 0 11224 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_127
timestamp 1649977179
transform 1 0 12788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_184
timestamp 1649977179
transform 1 0 18032 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_217
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_223
timestamp 1649977179
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1649977179
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_255
timestamp 1649977179
transform 1 0 24564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_297
timestamp 1649977179
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_305
timestamp 1649977179
transform 1 0 29164 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_311
timestamp 1649977179
transform 1 0 29716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_319
timestamp 1649977179
transform 1 0 30452 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_322
timestamp 1649977179
transform 1 0 30728 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_346
timestamp 1649977179
transform 1 0 32936 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_358
timestamp 1649977179
transform 1 0 34040 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_376
timestamp 1649977179
transform 1 0 35696 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_380
timestamp 1649977179
transform 1 0 36064 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_407
timestamp 1649977179
transform 1 0 38548 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1649977179
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_421
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_429
timestamp 1649977179
transform 1 0 40572 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_441
timestamp 1649977179
transform 1 0 41676 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_453
timestamp 1649977179
transform 1 0 42780 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_465
timestamp 1649977179
transform 1 0 43884 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_473
timestamp 1649977179
transform 1 0 44620 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_617
timestamp 1649977179
transform 1 0 57868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1649977179
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1649977179
transform 1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_41
timestamp 1649977179
transform 1 0 4876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_53
timestamp 1649977179
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_68
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_77
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_89
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1649977179
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_102
timestamp 1649977179
transform 1 0 10488 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_131
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_141
timestamp 1649977179
transform 1 0 14076 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_153
timestamp 1649977179
transform 1 0 15180 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_172
timestamp 1649977179
transform 1 0 16928 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_180
timestamp 1649977179
transform 1 0 17664 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_200
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_206
timestamp 1649977179
transform 1 0 20056 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_211
timestamp 1649977179
transform 1 0 20516 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_218
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_229
timestamp 1649977179
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_233
timestamp 1649977179
transform 1 0 22540 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1649977179
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_248
timestamp 1649977179
transform 1 0 23920 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_255
timestamp 1649977179
transform 1 0 24564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_267
timestamp 1649977179
transform 1 0 25668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_290
timestamp 1649977179
transform 1 0 27784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_302
timestamp 1649977179
transform 1 0 28888 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_310
timestamp 1649977179
transform 1 0 29624 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_322
timestamp 1649977179
transform 1 0 30728 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1649977179
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_343
timestamp 1649977179
transform 1 0 32660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_354
timestamp 1649977179
transform 1 0 33672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_362
timestamp 1649977179
transform 1 0 34408 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_374
timestamp 1649977179
transform 1 0 35512 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_381
timestamp 1649977179
transform 1 0 36156 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_387
timestamp 1649977179
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_401
timestamp 1649977179
transform 1 0 37996 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_409
timestamp 1649977179
transform 1 0 38732 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_426
timestamp 1649977179
transform 1 0 40296 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_438
timestamp 1649977179
transform 1 0 41400 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1649977179
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_16
timestamp 1649977179
transform 1 0 2576 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_37
timestamp 1649977179
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_40
timestamp 1649977179
transform 1 0 4784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_52
timestamp 1649977179
transform 1 0 5888 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_60
timestamp 1649977179
transform 1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1649977179
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_93
timestamp 1649977179
transform 1 0 9660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_111
timestamp 1649977179
transform 1 0 11316 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_146
timestamp 1649977179
transform 1 0 14536 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_152
timestamp 1649977179
transform 1 0 15088 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_164
timestamp 1649977179
transform 1 0 16192 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_167
timestamp 1649977179
transform 1 0 16468 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_183
timestamp 1649977179
transform 1 0 17940 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_205
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_212
timestamp 1649977179
transform 1 0 20608 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_222
timestamp 1649977179
transform 1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_229
timestamp 1649977179
transform 1 0 22172 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_236
timestamp 1649977179
transform 1 0 22816 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1649977179
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_255
timestamp 1649977179
transform 1 0 24564 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_269
timestamp 1649977179
transform 1 0 25852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_276
timestamp 1649977179
transform 1 0 26496 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_285
timestamp 1649977179
transform 1 0 27324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_297
timestamp 1649977179
transform 1 0 28428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1649977179
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_325
timestamp 1649977179
transform 1 0 31004 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_337
timestamp 1649977179
transform 1 0 32108 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_343
timestamp 1649977179
transform 1 0 32660 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_346
timestamp 1649977179
transform 1 0 32936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1649977179
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_371
timestamp 1649977179
transform 1 0 35236 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_382
timestamp 1649977179
transform 1 0 36248 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_388
timestamp 1649977179
transform 1 0 36800 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_399
timestamp 1649977179
transform 1 0 37812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_411
timestamp 1649977179
transform 1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_429
timestamp 1649977179
transform 1 0 40572 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_435
timestamp 1649977179
transform 1 0 41124 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_447
timestamp 1649977179
transform 1 0 42228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_459
timestamp 1649977179
transform 1 0 43332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_471
timestamp 1649977179
transform 1 0 44436 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_25
timestamp 1649977179
transform 1 0 3404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_38
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_50
timestamp 1649977179
transform 1 0 5704 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_70
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_76
timestamp 1649977179
transform 1 0 8096 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_80
timestamp 1649977179
transform 1 0 8464 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_96
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_155
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_173
timestamp 1649977179
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_182
timestamp 1649977179
transform 1 0 17848 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_206
timestamp 1649977179
transform 1 0 20056 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_239
timestamp 1649977179
transform 1 0 23092 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_253
timestamp 1649977179
transform 1 0 24380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_265
timestamp 1649977179
transform 1 0 25484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_286
timestamp 1649977179
transform 1 0 27416 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_292
timestamp 1649977179
transform 1 0 27968 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1649977179
transform 1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_310
timestamp 1649977179
transform 1 0 29624 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1649977179
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_345
timestamp 1649977179
transform 1 0 32844 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_362
timestamp 1649977179
transform 1 0 34408 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1649977179
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_400
timestamp 1649977179
transform 1 0 37904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_406
timestamp 1649977179
transform 1 0 38456 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_426
timestamp 1649977179
transform 1 0 40296 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_440
timestamp 1649977179
transform 1 0 41584 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1649977179
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_48
timestamp 1649977179
transform 1 0 5520 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_60
timestamp 1649977179
transform 1 0 6624 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1649977179
transform 1 0 9660 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_100
timestamp 1649977179
transform 1 0 10304 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_106
timestamp 1649977179
transform 1 0 10856 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_114
timestamp 1649977179
transform 1 0 11592 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_126
timestamp 1649977179
transform 1 0 12696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1649977179
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1649977179
transform 1 0 17572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1649977179
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_202
timestamp 1649977179
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_208
timestamp 1649977179
transform 1 0 20240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_214
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_226
timestamp 1649977179
transform 1 0 21896 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_232
timestamp 1649977179
transform 1 0 22448 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_238
timestamp 1649977179
transform 1 0 23000 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1649977179
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_267
timestamp 1649977179
transform 1 0 25668 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_273
timestamp 1649977179
transform 1 0 26220 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_279
timestamp 1649977179
transform 1 0 26772 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_285
timestamp 1649977179
transform 1 0 27324 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_297
timestamp 1649977179
transform 1 0 28428 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_302
timestamp 1649977179
transform 1 0 28888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_323
timestamp 1649977179
transform 1 0 30820 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_335
timestamp 1649977179
transform 1 0 31924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_347
timestamp 1649977179
transform 1 0 33028 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_351
timestamp 1649977179
transform 1 0 33396 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_369
timestamp 1649977179
transform 1 0 35052 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_372
timestamp 1649977179
transform 1 0 35328 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_384
timestamp 1649977179
transform 1 0 36432 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_395
timestamp 1649977179
transform 1 0 37444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_407
timestamp 1649977179
transform 1 0 38548 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_426
timestamp 1649977179
transform 1 0 40296 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_438
timestamp 1649977179
transform 1 0 41400 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_450
timestamp 1649977179
transform 1 0 42504 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_462
timestamp 1649977179
transform 1 0 43608 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_474
timestamp 1649977179
transform 1 0 44712 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_32
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_40
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_45
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_65
timestamp 1649977179
transform 1 0 7084 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_77
timestamp 1649977179
transform 1 0 8188 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_89
timestamp 1649977179
transform 1 0 9292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_101
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_116
timestamp 1649977179
transform 1 0 11776 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_133
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_185
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_210
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_230
timestamp 1649977179
transform 1 0 22264 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_234
timestamp 1649977179
transform 1 0 22632 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1649977179
transform 1 0 23644 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_259
timestamp 1649977179
transform 1 0 24932 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_275
timestamp 1649977179
transform 1 0 26404 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_289
timestamp 1649977179
transform 1 0 27692 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_301
timestamp 1649977179
transform 1 0 28796 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_313
timestamp 1649977179
transform 1 0 29900 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_319
timestamp 1649977179
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1649977179
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_347
timestamp 1649977179
transform 1 0 33028 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_359
timestamp 1649977179
transform 1 0 34132 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_371
timestamp 1649977179
transform 1 0 35236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1649977179
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_417
timestamp 1649977179
transform 1 0 39468 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_425
timestamp 1649977179
transform 1 0 40204 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_437
timestamp 1649977179
transform 1 0 41308 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_445
timestamp 1649977179
transform 1 0 42044 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1649977179
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_31
timestamp 1649977179
transform 1 0 3956 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_47
timestamp 1649977179
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_59
timestamp 1649977179
transform 1 0 6532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1649977179
transform 1 0 7268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_73
timestamp 1649977179
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1649977179
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_112
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_124
timestamp 1649977179
transform 1 0 12512 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_167
timestamp 1649977179
transform 1 0 16468 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_179
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_217
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_236
timestamp 1649977179
transform 1 0 22816 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1649977179
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_270
timestamp 1649977179
transform 1 0 25944 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1649977179
transform 1 0 26496 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_293
timestamp 1649977179
transform 1 0 28060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1649977179
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_328
timestamp 1649977179
transform 1 0 31280 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_340
timestamp 1649977179
transform 1 0 32384 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_348
timestamp 1649977179
transform 1 0 33120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_385
timestamp 1649977179
transform 1 0 36524 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_409
timestamp 1649977179
transform 1 0 38732 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1649977179
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_429
timestamp 1649977179
transform 1 0 40572 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_441
timestamp 1649977179
transform 1 0 41676 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_453
timestamp 1649977179
transform 1 0 42780 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_465
timestamp 1649977179
transform 1 0 43884 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_473
timestamp 1649977179
transform 1 0 44620 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_16
timestamp 1649977179
transform 1 0 2576 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_23
timestamp 1649977179
transform 1 0 3220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_38
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_46
timestamp 1649977179
transform 1 0 5336 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1649977179
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_71
timestamp 1649977179
transform 1 0 7636 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_79
timestamp 1649977179
transform 1 0 8372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_82
timestamp 1649977179
transform 1 0 8648 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_90
timestamp 1649977179
transform 1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_146
timestamp 1649977179
transform 1 0 14536 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_158
timestamp 1649977179
transform 1 0 15640 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_189
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_204
timestamp 1649977179
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_216
timestamp 1649977179
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_230
timestamp 1649977179
transform 1 0 22264 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_262
timestamp 1649977179
transform 1 0 25208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1649977179
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_285
timestamp 1649977179
transform 1 0 27324 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_297
timestamp 1649977179
transform 1 0 28428 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_309
timestamp 1649977179
transform 1 0 29532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_321
timestamp 1649977179
transform 1 0 30636 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1649977179
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_348
timestamp 1649977179
transform 1 0 33120 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_360
timestamp 1649977179
transform 1 0 34224 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_366
timestamp 1649977179
transform 1 0 34776 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_378
timestamp 1649977179
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1649977179
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_403
timestamp 1649977179
transform 1 0 38180 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_425
timestamp 1649977179
transform 1 0 40204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_437
timestamp 1649977179
transform 1 0 41308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_445
timestamp 1649977179
transform 1 0 42044 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1649977179
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_49
timestamp 1649977179
transform 1 0 5612 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_60
timestamp 1649977179
transform 1 0 6624 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_68
timestamp 1649977179
transform 1 0 7360 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_74
timestamp 1649977179
transform 1 0 7912 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_80
timestamp 1649977179
transform 1 0 8464 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_91
timestamp 1649977179
transform 1 0 9476 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_130
timestamp 1649977179
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_147
timestamp 1649977179
transform 1 0 14628 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_159
timestamp 1649977179
transform 1 0 15732 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1649977179
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_174
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_186
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_230
timestamp 1649977179
transform 1 0 22264 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_236
timestamp 1649977179
transform 1 0 22816 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_241
timestamp 1649977179
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1649977179
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_263
timestamp 1649977179
transform 1 0 25300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_267
timestamp 1649977179
transform 1 0 25668 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_273
timestamp 1649977179
transform 1 0 26220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_279
timestamp 1649977179
transform 1 0 26772 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_317
timestamp 1649977179
transform 1 0 30268 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_327
timestamp 1649977179
transform 1 0 31188 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_340
timestamp 1649977179
transform 1 0 32384 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1649977179
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_385
timestamp 1649977179
transform 1 0 36524 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_400
timestamp 1649977179
transform 1 0 37904 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_412
timestamp 1649977179
transform 1 0 39008 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_427
timestamp 1649977179
transform 1 0 40388 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_439
timestamp 1649977179
transform 1 0 41492 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_451
timestamp 1649977179
transform 1 0 42596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_463
timestamp 1649977179
transform 1 0 43700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_617
timestamp 1649977179
transform 1 0 57868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1649977179
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_25
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_76
timestamp 1649977179
transform 1 0 8096 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_82
timestamp 1649977179
transform 1 0 8648 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1649977179
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1649977179
transform 1 0 11960 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_124
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_136
timestamp 1649977179
transform 1 0 13616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_145
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp 1649977179
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_232
timestamp 1649977179
transform 1 0 22448 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_238
timestamp 1649977179
transform 1 0 23000 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_250
timestamp 1649977179
transform 1 0 24104 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_269
timestamp 1649977179
transform 1 0 25852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1649977179
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_287
timestamp 1649977179
transform 1 0 27508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_306
timestamp 1649977179
transform 1 0 29256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_320
timestamp 1649977179
transform 1 0 30544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_330
timestamp 1649977179
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_359
timestamp 1649977179
transform 1 0 34132 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_371
timestamp 1649977179
transform 1 0 35236 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1649977179
transform 1 0 36432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_403
timestamp 1649977179
transform 1 0 38180 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_425
timestamp 1649977179
transform 1 0 40204 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_434
timestamp 1649977179
transform 1 0 41032 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_446
timestamp 1649977179
transform 1 0 42136 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_16
timestamp 1649977179
transform 1 0 2576 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_39
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_43
timestamp 1649977179
transform 1 0 5060 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_46
timestamp 1649977179
transform 1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_52
timestamp 1649977179
transform 1 0 5888 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_62
timestamp 1649977179
transform 1 0 6808 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_72
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_90
timestamp 1649977179
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_96
timestamp 1649977179
transform 1 0 9936 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_108
timestamp 1649977179
transform 1 0 11040 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1649977179
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_119
timestamp 1649977179
transform 1 0 12052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1649977179
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_146
timestamp 1649977179
transform 1 0 14536 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_155
timestamp 1649977179
transform 1 0 15364 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_173
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_185
timestamp 1649977179
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1649977179
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_227
timestamp 1649977179
transform 1 0 21988 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_276
timestamp 1649977179
transform 1 0 26496 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_285
timestamp 1649977179
transform 1 0 27324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_291
timestamp 1649977179
transform 1 0 27876 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1649977179
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_322
timestamp 1649977179
transform 1 0 30728 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_334
timestamp 1649977179
transform 1 0 31832 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_342
timestamp 1649977179
transform 1 0 32568 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_351
timestamp 1649977179
transform 1 0 33396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_395
timestamp 1649977179
transform 1 0 37444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1649977179
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_425
timestamp 1649977179
transform 1 0 40204 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_434
timestamp 1649977179
transform 1 0 41032 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_440
timestamp 1649977179
transform 1 0 41584 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_452
timestamp 1649977179
transform 1 0 42688 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_464
timestamp 1649977179
transform 1 0 43792 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_617
timestamp 1649977179
transform 1 0 57868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1649977179
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_43
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_61
timestamp 1649977179
transform 1 0 6716 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_68
timestamp 1649977179
transform 1 0 7360 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_78
timestamp 1649977179
transform 1 0 8280 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_90
timestamp 1649977179
transform 1 0 9384 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_188
timestamp 1649977179
transform 1 0 18400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_229
timestamp 1649977179
transform 1 0 22172 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_254
timestamp 1649977179
transform 1 0 24472 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1649977179
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_289
timestamp 1649977179
transform 1 0 27692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_297
timestamp 1649977179
transform 1 0 28428 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_302
timestamp 1649977179
transform 1 0 28888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_313
timestamp 1649977179
transform 1 0 29900 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_323
timestamp 1649977179
transform 1 0 30820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_341
timestamp 1649977179
transform 1 0 32476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_350
timestamp 1649977179
transform 1 0 33304 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_370
timestamp 1649977179
transform 1 0 35144 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_382
timestamp 1649977179
transform 1 0 36248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1649977179
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_400
timestamp 1649977179
transform 1 0 37904 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_408
timestamp 1649977179
transform 1 0 38640 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_426
timestamp 1649977179
transform 1 0 40296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_438
timestamp 1649977179
transform 1 0 41400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1649977179
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1649977179
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_37
timestamp 1649977179
transform 1 0 4508 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_49
timestamp 1649977179
transform 1 0 5612 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_54
timestamp 1649977179
transform 1 0 6072 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_62
timestamp 1649977179
transform 1 0 6808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_74
timestamp 1649977179
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1649977179
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_93
timestamp 1649977179
transform 1 0 9660 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_103
timestamp 1649977179
transform 1 0 10580 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_111
timestamp 1649977179
transform 1 0 11316 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_117
timestamp 1649977179
transform 1 0 11868 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1649977179
transform 1 0 12604 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1649977179
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_149
timestamp 1649977179
transform 1 0 14812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_162
timestamp 1649977179
transform 1 0 16008 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_182
timestamp 1649977179
transform 1 0 17848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1649977179
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_203
timestamp 1649977179
transform 1 0 19780 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_212
timestamp 1649977179
transform 1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_220
timestamp 1649977179
transform 1 0 21344 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_224
timestamp 1649977179
transform 1 0 21712 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_227
timestamp 1649977179
transform 1 0 21988 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_239
timestamp 1649977179
transform 1 0 23092 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1649977179
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_287
timestamp 1649977179
transform 1 0 27508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_295
timestamp 1649977179
transform 1 0 28244 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_298
timestamp 1649977179
transform 1 0 28520 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1649977179
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_317
timestamp 1649977179
transform 1 0 30268 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_329
timestamp 1649977179
transform 1 0 31372 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_341
timestamp 1649977179
transform 1 0 32476 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_353
timestamp 1649977179
transform 1 0 33580 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_361
timestamp 1649977179
transform 1 0 34316 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_393
timestamp 1649977179
transform 1 0 37260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_396
timestamp 1649977179
transform 1 0 37536 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_408
timestamp 1649977179
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_432
timestamp 1649977179
transform 1 0 40848 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_438
timestamp 1649977179
transform 1 0 41400 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_450
timestamp 1649977179
transform 1 0 42504 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_462
timestamp 1649977179
transform 1 0 43608 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_474
timestamp 1649977179
transform 1 0 44712 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_19
timestamp 1649977179
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_35
timestamp 1649977179
transform 1 0 4324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_43
timestamp 1649977179
transform 1 0 5060 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1649977179
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_73
timestamp 1649977179
transform 1 0 7820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_85
timestamp 1649977179
transform 1 0 8924 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1649977179
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1649977179
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_145
timestamp 1649977179
transform 1 0 14444 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_151
timestamp 1649977179
transform 1 0 14996 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1649977179
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_184
timestamp 1649977179
transform 1 0 18032 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_196
timestamp 1649977179
transform 1 0 19136 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_204
timestamp 1649977179
transform 1 0 19872 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_207
timestamp 1649977179
transform 1 0 20148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_215
timestamp 1649977179
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_231
timestamp 1649977179
transform 1 0 22356 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_251
timestamp 1649977179
transform 1 0 24196 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_260
timestamp 1649977179
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1649977179
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_287
timestamp 1649977179
transform 1 0 27508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_299
timestamp 1649977179
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_315
timestamp 1649977179
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1649977179
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_343
timestamp 1649977179
transform 1 0 32660 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_399
timestamp 1649977179
transform 1 0 37812 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_402
timestamp 1649977179
transform 1 0 38088 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_414
timestamp 1649977179
transform 1 0 39192 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_426
timestamp 1649977179
transform 1 0 40296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 1649977179
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1649977179
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_621
timestamp 1649977179
transform 1 0 58236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_45
timestamp 1649977179
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 1649977179
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_72
timestamp 1649977179
transform 1 0 7728 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_78
timestamp 1649977179
transform 1 0 8280 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_36_87
timestamp 1649977179
transform 1 0 9108 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_102
timestamp 1649977179
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1649977179
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_119
timestamp 1649977179
transform 1 0 12052 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_131
timestamp 1649977179
transform 1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1649977179
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1649977179
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_151
timestamp 1649977179
transform 1 0 14996 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_160
timestamp 1649977179
transform 1 0 15824 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_174
timestamp 1649977179
transform 1 0 17112 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_186
timestamp 1649977179
transform 1 0 18216 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1649977179
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1649977179
transform 1 0 20700 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_219
timestamp 1649977179
transform 1 0 21252 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_229
timestamp 1649977179
transform 1 0 22172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_241
timestamp 1649977179
transform 1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1649977179
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_285
timestamp 1649977179
transform 1 0 27324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1649977179
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_340
timestamp 1649977179
transform 1 0 32384 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_351
timestamp 1649977179
transform 1 0 33396 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_395
timestamp 1649977179
transform 1 0 37444 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_412
timestamp 1649977179
transform 1 0 39008 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1649977179
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1649977179
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1649977179
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1649977179
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1649977179
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_10
timestamp 1649977179
transform 1 0 2024 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_30
timestamp 1649977179
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_75
timestamp 1649977179
transform 1 0 8004 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_82
timestamp 1649977179
transform 1 0 8648 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_94
timestamp 1649977179
transform 1 0 9752 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_100
timestamp 1649977179
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1649977179
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_141
timestamp 1649977179
transform 1 0 14076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_153
timestamp 1649977179
transform 1 0 15180 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_156
timestamp 1649977179
transform 1 0 15456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_162
timestamp 1649977179
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_171
timestamp 1649977179
transform 1 0 16836 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_199
timestamp 1649977179
transform 1 0 19412 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_208
timestamp 1649977179
transform 1 0 20240 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_219
timestamp 1649977179
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_245
timestamp 1649977179
transform 1 0 23644 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_248
timestamp 1649977179
transform 1 0 23920 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1649977179
transform 1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1649977179
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1649977179
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_286
timestamp 1649977179
transform 1 0 27416 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_294
timestamp 1649977179
transform 1 0 28152 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_300
timestamp 1649977179
transform 1 0 28704 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_312
timestamp 1649977179
transform 1 0 29808 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_324
timestamp 1649977179
transform 1 0 30912 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_340
timestamp 1649977179
transform 1 0 32384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_352
timestamp 1649977179
transform 1 0 33488 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_362
timestamp 1649977179
transform 1 0 34408 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_374
timestamp 1649977179
transform 1 0 35512 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_382
timestamp 1649977179
transform 1 0 36248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_390
timestamp 1649977179
transform 1 0 36984 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_398
timestamp 1649977179
transform 1 0 37720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_402
timestamp 1649977179
transform 1 0 38088 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_408
timestamp 1649977179
transform 1 0 38640 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_420
timestamp 1649977179
transform 1 0 39744 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_424
timestamp 1649977179
transform 1 0 40112 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_436
timestamp 1649977179
transform 1 0 41216 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_621
timestamp 1649977179
transform 1 0 58236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1649977179
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1649977179
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_31
timestamp 1649977179
transform 1 0 3956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_43
timestamp 1649977179
transform 1 0 5060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_55
timestamp 1649977179
transform 1 0 6164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_61
timestamp 1649977179
transform 1 0 6716 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_72
timestamp 1649977179
transform 1 0 7728 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_78
timestamp 1649977179
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_101
timestamp 1649977179
transform 1 0 10396 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_123
timestamp 1649977179
transform 1 0 12420 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1649977179
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_145
timestamp 1649977179
transform 1 0 14444 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_156
timestamp 1649977179
transform 1 0 15456 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_182
timestamp 1649977179
transform 1 0 17848 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1649977179
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_212
timestamp 1649977179
transform 1 0 20608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_236
timestamp 1649977179
transform 1 0 22816 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_246
timestamp 1649977179
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_263
timestamp 1649977179
transform 1 0 25300 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_285
timestamp 1649977179
transform 1 0 27324 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_297
timestamp 1649977179
transform 1 0 28428 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1649977179
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_341
timestamp 1649977179
transform 1 0 32476 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1649977179
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_374
timestamp 1649977179
transform 1 0 35512 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_394
timestamp 1649977179
transform 1 0 37352 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_406
timestamp 1649977179
transform 1 0 38456 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1649977179
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_432
timestamp 1649977179
transform 1 0 40848 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_444
timestamp 1649977179
transform 1 0 41952 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_456
timestamp 1649977179
transform 1 0 43056 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_468
timestamp 1649977179
transform 1 0 44160 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_11
timestamp 1649977179
transform 1 0 2116 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_17
timestamp 1649977179
transform 1 0 2668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 1649977179
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_41
timestamp 1649977179
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1649977179
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1649977179
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_72
timestamp 1649977179
transform 1 0 7728 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_78
timestamp 1649977179
transform 1 0 8280 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_84
timestamp 1649977179
transform 1 0 8832 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_87
timestamp 1649977179
transform 1 0 9108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_99
timestamp 1649977179
transform 1 0 10212 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1649977179
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_120
timestamp 1649977179
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_124
timestamp 1649977179
transform 1 0 12512 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_127
timestamp 1649977179
transform 1 0 12788 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_147
timestamp 1649977179
transform 1 0 14628 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_153
timestamp 1649977179
transform 1 0 15180 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_159
timestamp 1649977179
transform 1 0 15732 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1649977179
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_178
timestamp 1649977179
transform 1 0 17480 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_190
timestamp 1649977179
transform 1 0 18584 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_202
timestamp 1649977179
transform 1 0 19688 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_214
timestamp 1649977179
transform 1 0 20792 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1649977179
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_239
timestamp 1649977179
transform 1 0 23092 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_251
timestamp 1649977179
transform 1 0 24196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1649977179
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_297
timestamp 1649977179
transform 1 0 28428 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_300
timestamp 1649977179
transform 1 0 28704 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_312
timestamp 1649977179
transform 1 0 29808 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_318
timestamp 1649977179
transform 1 0 30360 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_330
timestamp 1649977179
transform 1 0 31464 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_347
timestamp 1649977179
transform 1 0 33028 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_357
timestamp 1649977179
transform 1 0 33948 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_369
timestamp 1649977179
transform 1 0 35052 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_382
timestamp 1649977179
transform 1 0 36248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1649977179
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_396
timestamp 1649977179
transform 1 0 37536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_402
timestamp 1649977179
transform 1 0 38088 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_408
timestamp 1649977179
transform 1 0 38640 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_425
timestamp 1649977179
transform 1 0 40204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_437
timestamp 1649977179
transform 1 0 41308 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_443
timestamp 1649977179
transform 1 0 41860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_31
timestamp 1649977179
transform 1 0 3956 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_43
timestamp 1649977179
transform 1 0 5060 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_55
timestamp 1649977179
transform 1 0 6164 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_67
timestamp 1649977179
transform 1 0 7268 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_79
timestamp 1649977179
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_101
timestamp 1649977179
transform 1 0 10396 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_110
timestamp 1649977179
transform 1 0 11224 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1649977179
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1649977179
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_149
timestamp 1649977179
transform 1 0 14812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_158
timestamp 1649977179
transform 1 0 15640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_166
timestamp 1649977179
transform 1 0 16376 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_174
timestamp 1649977179
transform 1 0 17112 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1649977179
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1649977179
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_202
timestamp 1649977179
transform 1 0 19688 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_214
timestamp 1649977179
transform 1 0 20792 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_218
timestamp 1649977179
transform 1 0 21160 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_227
timestamp 1649977179
transform 1 0 21988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_239
timestamp 1649977179
transform 1 0 23092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_261
timestamp 1649977179
transform 1 0 25116 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_281
timestamp 1649977179
transform 1 0 26956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_293
timestamp 1649977179
transform 1 0 28060 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1649977179
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_325
timestamp 1649977179
transform 1 0 31004 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_337
timestamp 1649977179
transform 1 0 32108 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_349
timestamp 1649977179
transform 1 0 33212 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1649977179
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_430
timestamp 1649977179
transform 1 0 40664 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_439
timestamp 1649977179
transform 1 0 41492 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_451
timestamp 1649977179
transform 1 0 42596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_463
timestamp 1649977179
transform 1 0 43700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1649977179
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_617
timestamp 1649977179
transform 1 0 57868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1649977179
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_32
timestamp 1649977179
transform 1 0 4048 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1649977179
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_59
timestamp 1649977179
transform 1 0 6532 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_71
timestamp 1649977179
transform 1 0 7636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_83
timestamp 1649977179
transform 1 0 8740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_88
timestamp 1649977179
transform 1 0 9200 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_100
timestamp 1649977179
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_116
timestamp 1649977179
transform 1 0 11776 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1649977179
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_132
timestamp 1649977179
transform 1 0 13248 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_138
timestamp 1649977179
transform 1 0 13800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1649977179
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1649977179
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_191
timestamp 1649977179
transform 1 0 18676 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_211
timestamp 1649977179
transform 1 0 20516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_229
timestamp 1649977179
transform 1 0 22172 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_238
timestamp 1649977179
transform 1 0 23000 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_250
timestamp 1649977179
transform 1 0 24104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_255
timestamp 1649977179
transform 1 0 24564 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_267
timestamp 1649977179
transform 1 0 25668 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_297
timestamp 1649977179
transform 1 0 28428 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_314
timestamp 1649977179
transform 1 0 29992 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_326
timestamp 1649977179
transform 1 0 31096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1649977179
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_344
timestamp 1649977179
transform 1 0 32752 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_356
timestamp 1649977179
transform 1 0 33856 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_368
timestamp 1649977179
transform 1 0 34960 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_380
timestamp 1649977179
transform 1 0 36064 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_398
timestamp 1649977179
transform 1 0 37720 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_406
timestamp 1649977179
transform 1 0 38456 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_425
timestamp 1649977179
transform 1 0 40204 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_433
timestamp 1649977179
transform 1 0 40940 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_445
timestamp 1649977179
transform 1 0 42044 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_9
timestamp 1649977179
transform 1 0 1932 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_12
timestamp 1649977179
transform 1 0 2208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1649977179
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_73
timestamp 1649977179
transform 1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1649977179
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1649977179
transform 1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_115
timestamp 1649977179
transform 1 0 11684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_127
timestamp 1649977179
transform 1 0 12788 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_131
timestamp 1649977179
transform 1 0 13156 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1649977179
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_147
timestamp 1649977179
transform 1 0 14628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_161
timestamp 1649977179
transform 1 0 15916 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_167
timestamp 1649977179
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_171
timestamp 1649977179
transform 1 0 16836 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_174
timestamp 1649977179
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_188
timestamp 1649977179
transform 1 0 18400 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_199
timestamp 1649977179
transform 1 0 19412 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_207
timestamp 1649977179
transform 1 0 20148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_219
timestamp 1649977179
transform 1 0 21252 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_230
timestamp 1649977179
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 1649977179
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1649977179
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_273
timestamp 1649977179
transform 1 0 26220 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1649977179
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_313
timestamp 1649977179
transform 1 0 29900 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1649977179
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_373
timestamp 1649977179
transform 1 0 35420 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_392
timestamp 1649977179
transform 1 0 37168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_404
timestamp 1649977179
transform 1 0 38272 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_412
timestamp 1649977179
transform 1 0 39008 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1649977179
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_429
timestamp 1649977179
transform 1 0 40572 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_441
timestamp 1649977179
transform 1 0 41676 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_453
timestamp 1649977179
transform 1 0 42780 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_465
timestamp 1649977179
transform 1 0 43884 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_473
timestamp 1649977179
transform 1 0 44620 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_617
timestamp 1649977179
transform 1 0 57868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1649977179
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_32
timestamp 1649977179
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_44
timestamp 1649977179
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1649977179
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_59
timestamp 1649977179
transform 1 0 6532 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_71
timestamp 1649977179
transform 1 0 7636 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_77
timestamp 1649977179
transform 1 0 8188 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1649977179
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_127
timestamp 1649977179
transform 1 0 12788 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_133
timestamp 1649977179
transform 1 0 13340 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_138
timestamp 1649977179
transform 1 0 13800 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_146
timestamp 1649977179
transform 1 0 14536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1649977179
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_172
timestamp 1649977179
transform 1 0 16928 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_184
timestamp 1649977179
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_188
timestamp 1649977179
transform 1 0 18400 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_194
timestamp 1649977179
transform 1 0 18952 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_203
timestamp 1649977179
transform 1 0 19780 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_211
timestamp 1649977179
transform 1 0 20516 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1649977179
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_241
timestamp 1649977179
transform 1 0 23276 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_253
timestamp 1649977179
transform 1 0 24380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_265
timestamp 1649977179
transform 1 0 25484 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_274
timestamp 1649977179
transform 1 0 26312 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_283
timestamp 1649977179
transform 1 0 27140 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_295
timestamp 1649977179
transform 1 0 28244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_304
timestamp 1649977179
transform 1 0 29072 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_327
timestamp 1649977179
transform 1 0 31188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_343
timestamp 1649977179
transform 1 0 32660 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_360
timestamp 1649977179
transform 1 0 34224 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_372
timestamp 1649977179
transform 1 0 35328 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_384
timestamp 1649977179
transform 1 0 36432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_396
timestamp 1649977179
transform 1 0 37536 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_402
timestamp 1649977179
transform 1 0 38088 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1649977179
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1649977179
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1649977179
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_34
timestamp 1649977179
transform 1 0 4232 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_44
timestamp 1649977179
transform 1 0 5152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_50
timestamp 1649977179
transform 1 0 5704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_62
timestamp 1649977179
transform 1 0 6808 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_66
timestamp 1649977179
transform 1 0 7176 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1649977179
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_113
timestamp 1649977179
transform 1 0 11500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_118
timestamp 1649977179
transform 1 0 11960 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_126
timestamp 1649977179
transform 1 0 12696 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1649977179
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_185
timestamp 1649977179
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1649977179
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_205
timestamp 1649977179
transform 1 0 19964 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_218
timestamp 1649977179
transform 1 0 21160 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_230
timestamp 1649977179
transform 1 0 22264 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_239
timestamp 1649977179
transform 1 0 23092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_263
timestamp 1649977179
transform 1 0 25300 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_283
timestamp 1649977179
transform 1 0 27140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_292
timestamp 1649977179
transform 1 0 27968 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_298
timestamp 1649977179
transform 1 0 28520 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_329
timestamp 1649977179
transform 1 0 31372 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_332
timestamp 1649977179
transform 1 0 31648 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1649977179
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_381
timestamp 1649977179
transform 1 0 36156 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_393
timestamp 1649977179
transform 1 0 37260 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_405
timestamp 1649977179
transform 1 0 38364 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1649977179
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_426
timestamp 1649977179
transform 1 0 40296 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_438
timestamp 1649977179
transform 1 0 41400 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_450
timestamp 1649977179
transform 1 0 42504 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_462
timestamp 1649977179
transform 1 0 43608 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_474
timestamp 1649977179
transform 1 0 44712 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_18
timestamp 1649977179
transform 1 0 2760 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_33
timestamp 1649977179
transform 1 0 4140 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_48
timestamp 1649977179
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_73
timestamp 1649977179
transform 1 0 7820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_85
timestamp 1649977179
transform 1 0 8924 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_99
timestamp 1649977179
transform 1 0 10212 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_103
timestamp 1649977179
transform 1 0 10580 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1649977179
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_115
timestamp 1649977179
transform 1 0 11684 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_129
timestamp 1649977179
transform 1 0 12972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_141
timestamp 1649977179
transform 1 0 14076 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_153
timestamp 1649977179
transform 1 0 15180 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_157
timestamp 1649977179
transform 1 0 15548 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1649977179
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_174
timestamp 1649977179
transform 1 0 17112 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_184
timestamp 1649977179
transform 1 0 18032 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_190
timestamp 1649977179
transform 1 0 18584 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_194
timestamp 1649977179
transform 1 0 18952 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_211
timestamp 1649977179
transform 1 0 20516 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1649977179
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_245
timestamp 1649977179
transform 1 0 23644 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_253
timestamp 1649977179
transform 1 0 24380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_256
timestamp 1649977179
transform 1 0 24656 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_268
timestamp 1649977179
transform 1 0 25760 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1649977179
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_310
timestamp 1649977179
transform 1 0 29624 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_322
timestamp 1649977179
transform 1 0 30728 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1649977179
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_348
timestamp 1649977179
transform 1 0 33120 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_356
timestamp 1649977179
transform 1 0 33856 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_368
timestamp 1649977179
transform 1 0 34960 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_380
timestamp 1649977179
transform 1 0 36064 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_423
timestamp 1649977179
transform 1 0 40020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_435
timestamp 1649977179
transform 1 0 41124 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1649977179
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1649977179
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_49
timestamp 1649977179
transform 1 0 5612 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_61
timestamp 1649977179
transform 1 0 6716 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_70
timestamp 1649977179
transform 1 0 7544 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1649977179
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1649977179
transform 1 0 9200 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_102
timestamp 1649977179
transform 1 0 10488 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_116
timestamp 1649977179
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1649977179
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_167
timestamp 1649977179
transform 1 0 16468 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_173
timestamp 1649977179
transform 1 0 17020 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_179
timestamp 1649977179
transform 1 0 17572 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_182
timestamp 1649977179
transform 1 0 17848 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_190
timestamp 1649977179
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_201
timestamp 1649977179
transform 1 0 19596 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1649977179
transform 1 0 20700 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1649977179
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1649977179
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_258
timestamp 1649977179
transform 1 0 24840 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_266
timestamp 1649977179
transform 1 0 25576 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_273
timestamp 1649977179
transform 1 0 26220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_293
timestamp 1649977179
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_299
timestamp 1649977179
transform 1 0 28612 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1649977179
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_311
timestamp 1649977179
transform 1 0 29716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_335
timestamp 1649977179
transform 1 0 31924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_346
timestamp 1649977179
transform 1 0 32936 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_370
timestamp 1649977179
transform 1 0 35144 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_382
timestamp 1649977179
transform 1 0 36248 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_394
timestamp 1649977179
transform 1 0 37352 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_406
timestamp 1649977179
transform 1 0 38456 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_418
timestamp 1649977179
transform 1 0 39560 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1649977179
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1649977179
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_65
timestamp 1649977179
transform 1 0 7084 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_77
timestamp 1649977179
transform 1 0 8188 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_85
timestamp 1649977179
transform 1 0 8924 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_92
timestamp 1649977179
transform 1 0 9568 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_98
timestamp 1649977179
transform 1 0 10120 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_104
timestamp 1649977179
transform 1 0 10672 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_118
timestamp 1649977179
transform 1 0 11960 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_131
timestamp 1649977179
transform 1 0 13156 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_140
timestamp 1649977179
transform 1 0 13984 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_148
timestamp 1649977179
transform 1 0 14720 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_151
timestamp 1649977179
transform 1 0 14996 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1649977179
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_177
timestamp 1649977179
transform 1 0 17388 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1649977179
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_197
timestamp 1649977179
transform 1 0 19228 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_201
timestamp 1649977179
transform 1 0 19596 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_212
timestamp 1649977179
transform 1 0 20608 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_257
timestamp 1649977179
transform 1 0 24748 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_269
timestamp 1649977179
transform 1 0 25852 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_276
timestamp 1649977179
transform 1 0 26496 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_285
timestamp 1649977179
transform 1 0 27324 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_297
timestamp 1649977179
transform 1 0 28428 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_301
timestamp 1649977179
transform 1 0 28796 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_304
timestamp 1649977179
transform 1 0 29072 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_318
timestamp 1649977179
transform 1 0 30360 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_339
timestamp 1649977179
transform 1 0 32292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_351
timestamp 1649977179
transform 1 0 33396 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_364
timestamp 1649977179
transform 1 0 34592 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_376
timestamp 1649977179
transform 1 0 35696 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1649977179
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_423
timestamp 1649977179
transform 1 0 40020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_435
timestamp 1649977179
transform 1 0 41124 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_621
timestamp 1649977179
transform 1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1649977179
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_34
timestamp 1649977179
transform 1 0 4232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_38
timestamp 1649977179
transform 1 0 4600 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_46
timestamp 1649977179
transform 1 0 5336 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_58
timestamp 1649977179
transform 1 0 6440 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_66
timestamp 1649977179
transform 1 0 7176 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_73
timestamp 1649977179
transform 1 0 7820 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_81
timestamp 1649977179
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_101
timestamp 1649977179
transform 1 0 10396 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_107
timestamp 1649977179
transform 1 0 10948 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_115
timestamp 1649977179
transform 1 0 11684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_120
timestamp 1649977179
transform 1 0 12144 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1649977179
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_149
timestamp 1649977179
transform 1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_169
timestamp 1649977179
transform 1 0 16652 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_224
timestamp 1649977179
transform 1 0 21712 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_232
timestamp 1649977179
transform 1 0 22448 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_237
timestamp 1649977179
transform 1 0 22908 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1649977179
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_263
timestamp 1649977179
transform 1 0 25300 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_275
timestamp 1649977179
transform 1 0 26404 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_287
timestamp 1649977179
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_299
timestamp 1649977179
transform 1 0 28612 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_323
timestamp 1649977179
transform 1 0 30820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_330
timestamp 1649977179
transform 1 0 31464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_336
timestamp 1649977179
transform 1 0 32016 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_344
timestamp 1649977179
transform 1 0 32752 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1649977179
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_372
timestamp 1649977179
transform 1 0 35328 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_385
timestamp 1649977179
transform 1 0 36524 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_409
timestamp 1649977179
transform 1 0 38732 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_417
timestamp 1649977179
transform 1 0 39468 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_26
timestamp 1649977179
transform 1 0 3496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_32
timestamp 1649977179
transform 1 0 4048 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_36
timestamp 1649977179
transform 1 0 4416 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_44
timestamp 1649977179
transform 1 0 5152 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_65
timestamp 1649977179
transform 1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_73
timestamp 1649977179
transform 1 0 7820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_82
timestamp 1649977179
transform 1 0 8648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_94
timestamp 1649977179
transform 1 0 9752 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1649977179
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_118
timestamp 1649977179
transform 1 0 11960 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_130
timestamp 1649977179
transform 1 0 13064 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_140
timestamp 1649977179
transform 1 0 13984 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_146
timestamp 1649977179
transform 1 0 14536 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_154
timestamp 1649977179
transform 1 0 15272 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_173
timestamp 1649977179
transform 1 0 17020 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_185
timestamp 1649977179
transform 1 0 18124 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_201
timestamp 1649977179
transform 1 0 19596 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_209
timestamp 1649977179
transform 1 0 20332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_221
timestamp 1649977179
transform 1 0 21436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1649977179
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_236
timestamp 1649977179
transform 1 0 22816 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_247
timestamp 1649977179
transform 1 0 23828 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_259
timestamp 1649977179
transform 1 0 24932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_267
timestamp 1649977179
transform 1 0 25668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_310
timestamp 1649977179
transform 1 0 29624 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_319
timestamp 1649977179
transform 1 0 30452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_326
timestamp 1649977179
transform 1 0 31096 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1649977179
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_355
timestamp 1649977179
transform 1 0 33764 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_367
timestamp 1649977179
transform 1 0 34868 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_376
timestamp 1649977179
transform 1 0 35696 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1649977179
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_395
timestamp 1649977179
transform 1 0 37444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_401
timestamp 1649977179
transform 1 0 37996 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_418
timestamp 1649977179
transform 1 0 39560 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_430
timestamp 1649977179
transform 1 0 40664 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_442
timestamp 1649977179
transform 1 0 41768 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_11
timestamp 1649977179
transform 1 0 2116 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_20
timestamp 1649977179
transform 1 0 2944 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_31
timestamp 1649977179
transform 1 0 3956 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_42
timestamp 1649977179
transform 1 0 4968 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_54
timestamp 1649977179
transform 1 0 6072 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_66
timestamp 1649977179
transform 1 0 7176 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_72
timestamp 1649977179
transform 1 0 7728 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_75
timestamp 1649977179
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_90
timestamp 1649977179
transform 1 0 9384 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_98
timestamp 1649977179
transform 1 0 10120 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_118
timestamp 1649977179
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_130
timestamp 1649977179
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1649977179
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_170
timestamp 1649977179
transform 1 0 16744 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_178
timestamp 1649977179
transform 1 0 17480 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_183
timestamp 1649977179
transform 1 0 17940 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_200
timestamp 1649977179
transform 1 0 19504 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_215
timestamp 1649977179
transform 1 0 20884 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_236
timestamp 1649977179
transform 1 0 22816 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_242
timestamp 1649977179
transform 1 0 23368 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1649977179
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_257
timestamp 1649977179
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_261
timestamp 1649977179
transform 1 0 25116 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_278
timestamp 1649977179
transform 1 0 26680 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_290
timestamp 1649977179
transform 1 0 27784 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_302
timestamp 1649977179
transform 1 0 28888 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_313
timestamp 1649977179
transform 1 0 29900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_319
timestamp 1649977179
transform 1 0 30452 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_331
timestamp 1649977179
transform 1 0 31556 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_351
timestamp 1649977179
transform 1 0 33396 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1649977179
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_368
timestamp 1649977179
transform 1 0 34960 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_384
timestamp 1649977179
transform 1 0 36432 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_396
timestamp 1649977179
transform 1 0 37536 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_408
timestamp 1649977179
transform 1 0 38640 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_617
timestamp 1649977179
transform 1 0 57868 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_621
timestamp 1649977179
transform 1 0 58236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_11
timestamp 1649977179
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_30
timestamp 1649977179
transform 1 0 3864 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_42
timestamp 1649977179
transform 1 0 4968 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1649977179
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_91
timestamp 1649977179
transform 1 0 9476 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_103
timestamp 1649977179
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_115
timestamp 1649977179
transform 1 0 11684 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_124
timestamp 1649977179
transform 1 0 12512 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_130
timestamp 1649977179
transform 1 0 13064 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_142
timestamp 1649977179
transform 1 0 14168 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_156
timestamp 1649977179
transform 1 0 15456 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_162
timestamp 1649977179
transform 1 0 16008 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_175
timestamp 1649977179
transform 1 0 17204 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1649977179
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_211
timestamp 1649977179
transform 1 0 20516 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1649977179
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_236
timestamp 1649977179
transform 1 0 22816 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_244
timestamp 1649977179
transform 1 0 23552 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_250
timestamp 1649977179
transform 1 0 24104 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_254
timestamp 1649977179
transform 1 0 24472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_263
timestamp 1649977179
transform 1 0 25300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_271
timestamp 1649977179
transform 1 0 26036 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_283
timestamp 1649977179
transform 1 0 27140 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_291
timestamp 1649977179
transform 1 0 27876 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_309
timestamp 1649977179
transform 1 0 29532 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_320
timestamp 1649977179
transform 1 0 30544 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_326
timestamp 1649977179
transform 1 0 31096 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_347
timestamp 1649977179
transform 1 0 33028 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_358
timestamp 1649977179
transform 1 0 34040 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_370
timestamp 1649977179
transform 1 0 35144 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_379
timestamp 1649977179
transform 1 0 35972 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1649977179
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1649977179
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1649977179
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1649977179
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1649977179
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_45
timestamp 1649977179
transform 1 0 5244 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_62
timestamp 1649977179
transform 1 0 6808 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_71
timestamp 1649977179
transform 1 0 7636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_127
timestamp 1649977179
transform 1 0 12788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_143
timestamp 1649977179
transform 1 0 14260 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_147
timestamp 1649977179
transform 1 0 14628 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_164
timestamp 1649977179
transform 1 0 16192 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_176
timestamp 1649977179
transform 1 0 17296 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_180
timestamp 1649977179
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1649977179
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_213
timestamp 1649977179
transform 1 0 20700 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_238
timestamp 1649977179
transform 1 0 23000 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1649977179
transform 1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_263
timestamp 1649977179
transform 1 0 25300 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_283
timestamp 1649977179
transform 1 0 27140 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_291
timestamp 1649977179
transform 1 0 27876 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1649977179
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_325
timestamp 1649977179
transform 1 0 31004 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_334
timestamp 1649977179
transform 1 0 31832 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_353
timestamp 1649977179
transform 1 0 33580 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1649977179
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_373
timestamp 1649977179
transform 1 0 35420 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_385
timestamp 1649977179
transform 1 0 36524 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_397
timestamp 1649977179
transform 1 0 37628 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1649977179
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_617
timestamp 1649977179
transform 1 0 57868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_621
timestamp 1649977179
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_19
timestamp 1649977179
transform 1 0 2852 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_28
timestamp 1649977179
transform 1 0 3680 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_40
timestamp 1649977179
transform 1 0 4784 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_46
timestamp 1649977179
transform 1 0 5336 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1649977179
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1649977179
transform 1 0 7820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_79
timestamp 1649977179
transform 1 0 8372 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_97
timestamp 1649977179
transform 1 0 10028 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_106
timestamp 1649977179
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_126
timestamp 1649977179
transform 1 0 12696 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_138
timestamp 1649977179
transform 1 0 13800 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_154
timestamp 1649977179
transform 1 0 15272 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1649977179
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_177
timestamp 1649977179
transform 1 0 17388 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_182
timestamp 1649977179
transform 1 0 17848 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_194
timestamp 1649977179
transform 1 0 18952 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_198
timestamp 1649977179
transform 1 0 19320 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_204
timestamp 1649977179
transform 1 0 19872 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_218
timestamp 1649977179
transform 1 0 21160 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_234
timestamp 1649977179
transform 1 0 22632 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_243
timestamp 1649977179
transform 1 0 23460 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_252
timestamp 1649977179
transform 1 0 24288 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_258
timestamp 1649977179
transform 1 0 24840 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1649977179
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1649977179
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_286
timestamp 1649977179
transform 1 0 27416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_295
timestamp 1649977179
transform 1 0 28244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_319
timestamp 1649977179
transform 1 0 30452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_330
timestamp 1649977179
transform 1 0 31464 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_339
timestamp 1649977179
transform 1 0 32292 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_351
timestamp 1649977179
transform 1 0 33396 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_363
timestamp 1649977179
transform 1 0 34500 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_374
timestamp 1649977179
transform 1 0 35512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_386
timestamp 1649977179
transform 1 0 36616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_395
timestamp 1649977179
transform 1 0 37444 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_7
timestamp 1649977179
transform 1 0 1748 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1649977179
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_50
timestamp 1649977179
transform 1 0 5704 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_54
timestamp 1649977179
transform 1 0 6072 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_63
timestamp 1649977179
transform 1 0 6900 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_69
timestamp 1649977179
transform 1 0 7452 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1649977179
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_91
timestamp 1649977179
transform 1 0 9476 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_108
timestamp 1649977179
transform 1 0 11040 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_116
timestamp 1649977179
transform 1 0 11776 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_143
timestamp 1649977179
transform 1 0 14260 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_155
timestamp 1649977179
transform 1 0 15364 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_163
timestamp 1649977179
transform 1 0 16100 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_168
timestamp 1649977179
transform 1 0 16560 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1649977179
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_215
timestamp 1649977179
transform 1 0 20884 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_218
timestamp 1649977179
transform 1 0 21160 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_232
timestamp 1649977179
transform 1 0 22448 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_236
timestamp 1649977179
transform 1 0 22816 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_239
timestamp 1649977179
transform 1 0 23092 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1649977179
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_281
timestamp 1649977179
transform 1 0 26956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_302
timestamp 1649977179
transform 1 0 28888 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_313
timestamp 1649977179
transform 1 0 29900 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_317
timestamp 1649977179
transform 1 0 30268 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_329
timestamp 1649977179
transform 1 0 31372 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_337
timestamp 1649977179
transform 1 0 32108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_346
timestamp 1649977179
transform 1 0 32936 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_358
timestamp 1649977179
transform 1 0 34040 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_369
timestamp 1649977179
transform 1 0 35052 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_375
timestamp 1649977179
transform 1 0 35604 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_387
timestamp 1649977179
transform 1 0 36708 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_399
timestamp 1649977179
transform 1 0 37812 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_411
timestamp 1649977179
transform 1 0 38916 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1649977179
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_43
timestamp 1649977179
transform 1 0 5060 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_46
timestamp 1649977179
transform 1 0 5336 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1649977179
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_59
timestamp 1649977179
transform 1 0 6532 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_79
timestamp 1649977179
transform 1 0 8372 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_88
timestamp 1649977179
transform 1 0 9200 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1649977179
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_131
timestamp 1649977179
transform 1 0 13156 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_142
timestamp 1649977179
transform 1 0 14168 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_154
timestamp 1649977179
transform 1 0 15272 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1649977179
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_174
timestamp 1649977179
transform 1 0 17112 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_188
timestamp 1649977179
transform 1 0 18400 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_196
timestamp 1649977179
transform 1 0 19136 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_202
timestamp 1649977179
transform 1 0 19688 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1649977179
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1649977179
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_230
timestamp 1649977179
transform 1 0 22264 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_234
timestamp 1649977179
transform 1 0 22632 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_245
timestamp 1649977179
transform 1 0 23644 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_255
timestamp 1649977179
transform 1 0 24564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1649977179
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_296
timestamp 1649977179
transform 1 0 28336 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_307
timestamp 1649977179
transform 1 0 29348 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_313
timestamp 1649977179
transform 1 0 29900 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_322
timestamp 1649977179
transform 1 0 30728 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1649977179
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_341
timestamp 1649977179
transform 1 0 32476 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_358
timestamp 1649977179
transform 1 0 34040 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_370
timestamp 1649977179
transform 1 0 35144 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_376
timestamp 1649977179
transform 1 0 35696 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_379
timestamp 1649977179
transform 1 0 35972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_411
timestamp 1649977179
transform 1 0 38916 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_423
timestamp 1649977179
transform 1 0 40020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_435
timestamp 1649977179
transform 1 0 41124 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_621
timestamp 1649977179
transform 1 0 58236 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_31
timestamp 1649977179
transform 1 0 3956 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_39
timestamp 1649977179
transform 1 0 4692 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_61
timestamp 1649977179
transform 1 0 6716 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_73
timestamp 1649977179
transform 1 0 7820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_79
timestamp 1649977179
transform 1 0 8372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_102
timestamp 1649977179
transform 1 0 10488 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_114
timestamp 1649977179
transform 1 0 11592 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_124
timestamp 1649977179
transform 1 0 12512 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1649977179
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_151
timestamp 1649977179
transform 1 0 14996 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_173
timestamp 1649977179
transform 1 0 17020 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_181
timestamp 1649977179
transform 1 0 17756 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1649977179
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_213
timestamp 1649977179
transform 1 0 20700 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_226
timestamp 1649977179
transform 1 0 21896 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_238
timestamp 1649977179
transform 1 0 23000 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1649977179
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_263
timestamp 1649977179
transform 1 0 25300 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_275
timestamp 1649977179
transform 1 0 26404 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_287
timestamp 1649977179
transform 1 0 27508 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_295
timestamp 1649977179
transform 1 0 28244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_328
timestamp 1649977179
transform 1 0 31280 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_336
timestamp 1649977179
transform 1 0 32016 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_342
timestamp 1649977179
transform 1 0 32568 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_354
timestamp 1649977179
transform 1 0 33672 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_362
timestamp 1649977179
transform 1 0 34408 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1649977179
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_31
timestamp 1649977179
transform 1 0 3956 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_40
timestamp 1649977179
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1649977179
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_63
timestamp 1649977179
transform 1 0 6900 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_71
timestamp 1649977179
transform 1 0 7636 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_75
timestamp 1649977179
transform 1 0 8004 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_87
timestamp 1649977179
transform 1 0 9108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_99
timestamp 1649977179
transform 1 0 10212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_121
timestamp 1649977179
transform 1 0 12236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_128
timestamp 1649977179
transform 1 0 12880 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_148
timestamp 1649977179
transform 1 0 14720 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_156
timestamp 1649977179
transform 1 0 15456 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_177
timestamp 1649977179
transform 1 0 17388 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_185
timestamp 1649977179
transform 1 0 18124 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_192
timestamp 1649977179
transform 1 0 18768 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_198
timestamp 1649977179
transform 1 0 19320 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_204
timestamp 1649977179
transform 1 0 19872 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_216
timestamp 1649977179
transform 1 0 20976 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_251
timestamp 1649977179
transform 1 0 24196 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_255
timestamp 1649977179
transform 1 0 24564 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_264
timestamp 1649977179
transform 1 0 25392 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_270
timestamp 1649977179
transform 1 0 25944 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1649977179
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_299
timestamp 1649977179
transform 1 0 28612 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_307
timestamp 1649977179
transform 1 0 29348 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_310
timestamp 1649977179
transform 1 0 29624 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_318
timestamp 1649977179
transform 1 0 30360 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1649977179
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_350
timestamp 1649977179
transform 1 0 33304 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_359
timestamp 1649977179
transform 1 0 34132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_365
timestamp 1649977179
transform 1 0 34684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_382
timestamp 1649977179
transform 1 0 36248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1649977179
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_395
timestamp 1649977179
transform 1 0 37444 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_407
timestamp 1649977179
transform 1 0 38548 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_419
timestamp 1649977179
transform 1 0 39652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_431
timestamp 1649977179
transform 1 0 40756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_443
timestamp 1649977179
transform 1 0 41860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1649977179
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_9
timestamp 1649977179
transform 1 0 1932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_12
timestamp 1649977179
transform 1 0 2208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1649977179
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_37
timestamp 1649977179
transform 1 0 4508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_43
timestamp 1649977179
transform 1 0 5060 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_49
timestamp 1649977179
transform 1 0 5612 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_61
timestamp 1649977179
transform 1 0 6716 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_69
timestamp 1649977179
transform 1 0 7452 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_75
timestamp 1649977179
transform 1 0 8004 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_93
timestamp 1649977179
transform 1 0 9660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_105
timestamp 1649977179
transform 1 0 10764 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_110
timestamp 1649977179
transform 1 0 11224 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_122
timestamp 1649977179
transform 1 0 12328 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_134
timestamp 1649977179
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_151
timestamp 1649977179
transform 1 0 14996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_157
timestamp 1649977179
transform 1 0 15548 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_166
timestamp 1649977179
transform 1 0 16376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_175
timestamp 1649977179
transform 1 0 17204 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_181
timestamp 1649977179
transform 1 0 17756 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_184
timestamp 1649977179
transform 1 0 18032 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1649977179
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_201
timestamp 1649977179
transform 1 0 19596 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_210
timestamp 1649977179
transform 1 0 20424 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_216
timestamp 1649977179
transform 1 0 20976 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_228
timestamp 1649977179
transform 1 0 22080 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_240
timestamp 1649977179
transform 1 0 23184 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1649977179
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_261
timestamp 1649977179
transform 1 0 25116 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1649977179
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_280
timestamp 1649977179
transform 1 0 26864 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_292
timestamp 1649977179
transform 1 0 27968 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1649977179
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_313
timestamp 1649977179
transform 1 0 29900 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_325
timestamp 1649977179
transform 1 0 31004 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_334
timestamp 1649977179
transform 1 0 31832 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_348
timestamp 1649977179
transform 1 0 33120 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1649977179
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_381
timestamp 1649977179
transform 1 0 36156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_409
timestamp 1649977179
transform 1 0 38732 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_417
timestamp 1649977179
transform 1 0 39468 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_31
timestamp 1649977179
transform 1 0 3956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_40
timestamp 1649977179
transform 1 0 4784 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_46
timestamp 1649977179
transform 1 0 5336 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1649977179
transform 1 0 5612 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_63
timestamp 1649977179
transform 1 0 6900 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_72
timestamp 1649977179
transform 1 0 7728 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_78
timestamp 1649977179
transform 1 0 8280 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_90
timestamp 1649977179
transform 1 0 9384 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_98
timestamp 1649977179
transform 1 0 10120 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1649977179
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_115
timestamp 1649977179
transform 1 0 11684 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_128
timestamp 1649977179
transform 1 0 12880 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_140
timestamp 1649977179
transform 1 0 13984 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_152
timestamp 1649977179
transform 1 0 15088 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1649977179
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_171
timestamp 1649977179
transform 1 0 16836 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_175
timestamp 1649977179
transform 1 0 17204 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_189
timestamp 1649977179
transform 1 0 18492 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_200
timestamp 1649977179
transform 1 0 19504 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1649977179
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_241
timestamp 1649977179
transform 1 0 23276 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_247
timestamp 1649977179
transform 1 0 23828 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_250
timestamp 1649977179
transform 1 0 24104 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_262
timestamp 1649977179
transform 1 0 25208 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_271
timestamp 1649977179
transform 1 0 26036 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_283
timestamp 1649977179
transform 1 0 27140 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_289
timestamp 1649977179
transform 1 0 27692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_301
timestamp 1649977179
transform 1 0 28796 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_314
timestamp 1649977179
transform 1 0 29992 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_328
timestamp 1649977179
transform 1 0 31280 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_340
timestamp 1649977179
transform 1 0 32384 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_353
timestamp 1649977179
transform 1 0 33580 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_365
timestamp 1649977179
transform 1 0 34684 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_377
timestamp 1649977179
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1649977179
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_37
timestamp 1649977179
transform 1 0 4508 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_47
timestamp 1649977179
transform 1 0 5428 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_70
timestamp 1649977179
transform 1 0 7544 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_80
timestamp 1649977179
transform 1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_117
timestamp 1649977179
transform 1 0 11868 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1649977179
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_173
timestamp 1649977179
transform 1 0 17020 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_190
timestamp 1649977179
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_201
timestamp 1649977179
transform 1 0 19596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_207
timestamp 1649977179
transform 1 0 20148 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_215
timestamp 1649977179
transform 1 0 20884 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_219
timestamp 1649977179
transform 1 0 21252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_231
timestamp 1649977179
transform 1 0 22356 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_240
timestamp 1649977179
transform 1 0 23184 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1649977179
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_269
timestamp 1649977179
transform 1 0 25852 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_278
timestamp 1649977179
transform 1 0 26680 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_294
timestamp 1649977179
transform 1 0 28152 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_303
timestamp 1649977179
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_317
timestamp 1649977179
transform 1 0 30268 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_337
timestamp 1649977179
transform 1 0 32108 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_351
timestamp 1649977179
transform 1 0 33396 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_617
timestamp 1649977179
transform 1 0 57868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1649977179
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_45
timestamp 1649977179
transform 1 0 5244 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1649977179
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_85
timestamp 1649977179
transform 1 0 8924 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_91
timestamp 1649977179
transform 1 0 9476 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_102
timestamp 1649977179
transform 1 0 10488 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_108
timestamp 1649977179
transform 1 0 11040 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_118
timestamp 1649977179
transform 1 0 11960 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_127
timestamp 1649977179
transform 1 0 12788 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_135
timestamp 1649977179
transform 1 0 13524 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_141
timestamp 1649977179
transform 1 0 14076 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_147
timestamp 1649977179
transform 1 0 14628 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_159
timestamp 1649977179
transform 1 0 15732 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_180
timestamp 1649977179
transform 1 0 17664 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_186
timestamp 1649977179
transform 1 0 18216 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_198
timestamp 1649977179
transform 1 0 19320 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_210
timestamp 1649977179
transform 1 0 20424 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1649977179
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_231
timestamp 1649977179
transform 1 0 22356 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_239
timestamp 1649977179
transform 1 0 23092 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_245
timestamp 1649977179
transform 1 0 23644 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_267
timestamp 1649977179
transform 1 0 25668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_301
timestamp 1649977179
transform 1 0 28796 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_311
timestamp 1649977179
transform 1 0 29716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_323
timestamp 1649977179
transform 1 0 30820 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1649977179
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_347
timestamp 1649977179
transform 1 0 33028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_359
timestamp 1649977179
transform 1 0 34132 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_370
timestamp 1649977179
transform 1 0 35144 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_382
timestamp 1649977179
transform 1 0 36248 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1649977179
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_45
timestamp 1649977179
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_57
timestamp 1649977179
transform 1 0 6348 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_73
timestamp 1649977179
transform 1 0 7820 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_79
timestamp 1649977179
transform 1 0 8372 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_89
timestamp 1649977179
transform 1 0 9292 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_93
timestamp 1649977179
transform 1 0 9660 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_113
timestamp 1649977179
transform 1 0 11500 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_149
timestamp 1649977179
transform 1 0 14812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_155
timestamp 1649977179
transform 1 0 15364 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_163
timestamp 1649977179
transform 1 0 16100 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_166
timestamp 1649977179
transform 1 0 16376 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_178
timestamp 1649977179
transform 1 0 17480 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_190
timestamp 1649977179
transform 1 0 18584 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_234
timestamp 1649977179
transform 1 0 22632 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_238
timestamp 1649977179
transform 1 0 23000 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_241
timestamp 1649977179
transform 1 0 23276 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1649977179
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_255
timestamp 1649977179
transform 1 0 24564 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_267
timestamp 1649977179
transform 1 0 25668 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_279
timestamp 1649977179
transform 1 0 26772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_284
timestamp 1649977179
transform 1 0 27232 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_292
timestamp 1649977179
transform 1 0 27968 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1649977179
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_314
timestamp 1649977179
transform 1 0 29992 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_326
timestamp 1649977179
transform 1 0 31096 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_338
timestamp 1649977179
transform 1 0 32200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_341
timestamp 1649977179
transform 1 0 32476 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_349
timestamp 1649977179
transform 1 0 33212 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_356
timestamp 1649977179
transform 1 0 33856 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_373
timestamp 1649977179
transform 1 0 35420 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_385
timestamp 1649977179
transform 1 0 36524 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_397
timestamp 1649977179
transform 1 0 37628 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_409
timestamp 1649977179
transform 1 0 38732 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_417
timestamp 1649977179
transform 1 0 39468 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_617
timestamp 1649977179
transform 1 0 57868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1649977179
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_64
timestamp 1649977179
transform 1 0 6992 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_73
timestamp 1649977179
transform 1 0 7820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_85
timestamp 1649977179
transform 1 0 8924 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_106
timestamp 1649977179
transform 1 0 10856 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_123
timestamp 1649977179
transform 1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1649977179
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_151
timestamp 1649977179
transform 1 0 14996 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_155
timestamp 1649977179
transform 1 0 15364 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1649977179
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_174
timestamp 1649977179
transform 1 0 17112 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_185
timestamp 1649977179
transform 1 0 18124 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_197
timestamp 1649977179
transform 1 0 19228 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_231
timestamp 1649977179
transform 1 0 22356 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_242
timestamp 1649977179
transform 1 0 23368 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1649977179
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1649977179
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_289
timestamp 1649977179
transform 1 0 27692 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_294
timestamp 1649977179
transform 1 0 28152 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_306
timestamp 1649977179
transform 1 0 29256 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_318
timestamp 1649977179
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1649977179
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_367
timestamp 1649977179
transform 1 0 34868 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_371
timestamp 1649977179
transform 1 0 35236 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1649977179
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1649977179
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1649977179
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_31
timestamp 1649977179
transform 1 0 3956 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_43
timestamp 1649977179
transform 1 0 5060 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_51
timestamp 1649977179
transform 1 0 5796 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1649977179
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1649977179
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_112
timestamp 1649977179
transform 1 0 11408 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_136
timestamp 1649977179
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_149
timestamp 1649977179
transform 1 0 14812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_170
timestamp 1649977179
transform 1 0 16744 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_176
timestamp 1649977179
transform 1 0 17296 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1649977179
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_191
timestamp 1649977179
transform 1 0 18676 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_205
timestamp 1649977179
transform 1 0 19964 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_226
timestamp 1649977179
transform 1 0 21896 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_238
timestamp 1649977179
transform 1 0 23000 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1649977179
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_261
timestamp 1649977179
transform 1 0 25116 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_273
timestamp 1649977179
transform 1 0 26220 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_285
timestamp 1649977179
transform 1 0 27324 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_297
timestamp 1649977179
transform 1 0 28428 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1649977179
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_317
timestamp 1649977179
transform 1 0 30268 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_320
timestamp 1649977179
transform 1 0 30544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_334
timestamp 1649977179
transform 1 0 31832 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_342
timestamp 1649977179
transform 1 0 32568 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_348
timestamp 1649977179
transform 1 0 33120 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1649977179
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_381
timestamp 1649977179
transform 1 0 36156 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_393
timestamp 1649977179
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_405
timestamp 1649977179
transform 1 0 38364 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1649977179
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_25
timestamp 1649977179
transform 1 0 3404 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_34
timestamp 1649977179
transform 1 0 4232 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_43
timestamp 1649977179
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_67
timestamp 1649977179
transform 1 0 7268 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_79
timestamp 1649977179
transform 1 0 8372 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_91
timestamp 1649977179
transform 1 0 9476 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_103
timestamp 1649977179
transform 1 0 10580 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_120
timestamp 1649977179
transform 1 0 12144 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_132
timestamp 1649977179
transform 1 0 13248 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_145
timestamp 1649977179
transform 1 0 14444 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_157
timestamp 1649977179
transform 1 0 15548 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_165
timestamp 1649977179
transform 1 0 16284 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_201
timestamp 1649977179
transform 1 0 19596 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_213
timestamp 1649977179
transform 1 0 20700 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_219
timestamp 1649977179
transform 1 0 21252 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_267
timestamp 1649977179
transform 1 0 25668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1649977179
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_287
timestamp 1649977179
transform 1 0 27508 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_299
timestamp 1649977179
transform 1 0 28612 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_303
timestamp 1649977179
transform 1 0 28980 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_320
timestamp 1649977179
transform 1 0 30544 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_331
timestamp 1649977179
transform 1 0 31556 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_348
timestamp 1649977179
transform 1 0 33120 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_354
timestamp 1649977179
transform 1 0 33672 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_360
timestamp 1649977179
transform 1 0 34224 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_372
timestamp 1649977179
transform 1 0 35328 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_384
timestamp 1649977179
transform 1 0 36432 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_621
timestamp 1649977179
transform 1 0 58236 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_7
timestamp 1649977179
transform 1 0 1748 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1649977179
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_73
timestamp 1649977179
transform 1 0 7820 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_92
timestamp 1649977179
transform 1 0 9568 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_104
timestamp 1649977179
transform 1 0 10672 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_116
timestamp 1649977179
transform 1 0 11776 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_128
timestamp 1649977179
transform 1 0 12880 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_148
timestamp 1649977179
transform 1 0 14720 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_160
timestamp 1649977179
transform 1 0 15824 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_172
timestamp 1649977179
transform 1 0 16928 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_178
timestamp 1649977179
transform 1 0 17480 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_187
timestamp 1649977179
transform 1 0 18308 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_205
timestamp 1649977179
transform 1 0 19964 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_214
timestamp 1649977179
transform 1 0 20792 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_226
timestamp 1649977179
transform 1 0 21896 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_238
timestamp 1649977179
transform 1 0 23000 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1649977179
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_263
timestamp 1649977179
transform 1 0 25300 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_283
timestamp 1649977179
transform 1 0 27140 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_295
timestamp 1649977179
transform 1 0 28244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1649977179
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_315
timestamp 1649977179
transform 1 0 30084 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_332
timestamp 1649977179
transform 1 0 31648 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_340
timestamp 1649977179
transform 1 0 32384 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_359
timestamp 1649977179
transform 1 0 34132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_25
timestamp 1649977179
transform 1 0 3404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_31
timestamp 1649977179
transform 1 0 3956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_37
timestamp 1649977179
transform 1 0 4508 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_40
timestamp 1649977179
transform 1 0 4784 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 1649977179
transform 1 0 5888 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_62
timestamp 1649977179
transform 1 0 6808 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_68
timestamp 1649977179
transform 1 0 7360 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_79
timestamp 1649977179
transform 1 0 8372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_101
timestamp 1649977179
transform 1 0 10396 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_109
timestamp 1649977179
transform 1 0 11132 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_121
timestamp 1649977179
transform 1 0 12236 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_126
timestamp 1649977179
transform 1 0 12696 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_130
timestamp 1649977179
transform 1 0 13064 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_141
timestamp 1649977179
transform 1 0 14076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_153
timestamp 1649977179
transform 1 0 15180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_165
timestamp 1649977179
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_228
timestamp 1649977179
transform 1 0 22080 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_255
timestamp 1649977179
transform 1 0 24564 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_258
timestamp 1649977179
transform 1 0 24840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_270
timestamp 1649977179
transform 1 0 25944 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_276
timestamp 1649977179
transform 1 0 26496 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_291
timestamp 1649977179
transform 1 0 27876 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_315
timestamp 1649977179
transform 1 0 30084 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_327
timestamp 1649977179
transform 1 0 31188 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_342
timestamp 1649977179
transform 1 0 32568 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_354
timestamp 1649977179
transform 1 0 33672 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_366
timestamp 1649977179
transform 1 0 34776 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_378
timestamp 1649977179
transform 1 0 35880 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1649977179
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_621
timestamp 1649977179
transform 1 0 58236 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_35
timestamp 1649977179
transform 1 0 4324 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_52
timestamp 1649977179
transform 1 0 5888 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_66
timestamp 1649977179
transform 1 0 7176 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_72
timestamp 1649977179
transform 1 0 7728 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_103
timestamp 1649977179
transform 1 0 10580 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_126
timestamp 1649977179
transform 1 0 12696 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_138
timestamp 1649977179
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_172
timestamp 1649977179
transform 1 0 16928 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_184
timestamp 1649977179
transform 1 0 18032 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_213
timestamp 1649977179
transform 1 0 20700 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_219
timestamp 1649977179
transform 1 0 21252 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_228
timestamp 1649977179
transform 1 0 22080 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1649977179
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_299
timestamp 1649977179
transform 1 0 28612 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_313
timestamp 1649977179
transform 1 0 29900 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_319
timestamp 1649977179
transform 1 0 30452 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_341
timestamp 1649977179
transform 1 0 32476 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_353
timestamp 1649977179
transform 1 0 33580 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1649977179
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_31
timestamp 1649977179
transform 1 0 3956 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_40
timestamp 1649977179
transform 1 0 4784 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1649977179
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_62
timestamp 1649977179
transform 1 0 6808 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_82
timestamp 1649977179
transform 1 0 8648 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_102
timestamp 1649977179
transform 1 0 10488 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_108
timestamp 1649977179
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_129
timestamp 1649977179
transform 1 0 12972 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_141
timestamp 1649977179
transform 1 0 14076 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_147
timestamp 1649977179
transform 1 0 14628 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_164
timestamp 1649977179
transform 1 0 16192 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_179
timestamp 1649977179
transform 1 0 17572 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_203
timestamp 1649977179
transform 1 0 19780 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_209
timestamp 1649977179
transform 1 0 20332 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1649977179
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_231
timestamp 1649977179
transform 1 0 22356 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_240
timestamp 1649977179
transform 1 0 23184 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_260
timestamp 1649977179
transform 1 0 25024 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_272
timestamp 1649977179
transform 1 0 26128 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_289
timestamp 1649977179
transform 1 0 27692 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_297
timestamp 1649977179
transform 1 0 28428 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_309
timestamp 1649977179
transform 1 0 29532 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_313
timestamp 1649977179
transform 1 0 29900 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_316
timestamp 1649977179
transform 1 0 30176 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_328
timestamp 1649977179
transform 1 0 31280 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_37
timestamp 1649977179
transform 1 0 4508 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_43
timestamp 1649977179
transform 1 0 5060 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_47
timestamp 1649977179
transform 1 0 5428 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_50
timestamp 1649977179
transform 1 0 5704 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_70
timestamp 1649977179
transform 1 0 7544 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_82
timestamp 1649977179
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_101
timestamp 1649977179
transform 1 0 10396 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_110
timestamp 1649977179
transform 1 0 11224 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_118
timestamp 1649977179
transform 1 0 11960 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_135
timestamp 1649977179
transform 1 0 13524 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_145
timestamp 1649977179
transform 1 0 14444 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_151
timestamp 1649977179
transform 1 0 14996 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_171
timestamp 1649977179
transform 1 0 16836 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_179
timestamp 1649977179
transform 1 0 17572 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_183
timestamp 1649977179
transform 1 0 17940 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1649977179
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_205
timestamp 1649977179
transform 1 0 19964 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_229
timestamp 1649977179
transform 1 0 22172 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_241
timestamp 1649977179
transform 1 0 23276 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_247
timestamp 1649977179
transform 1 0 23828 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_283
timestamp 1649977179
transform 1 0 27140 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_300
timestamp 1649977179
transform 1 0 28704 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_617
timestamp 1649977179
transform 1 0 57868 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_621
timestamp 1649977179
transform 1 0 58236 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_102
timestamp 1649977179
transform 1 0 10488 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_108
timestamp 1649977179
transform 1 0 11040 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_121
timestamp 1649977179
transform 1 0 12236 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_130
timestamp 1649977179
transform 1 0 13064 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_136
timestamp 1649977179
transform 1 0 13616 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_156
timestamp 1649977179
transform 1 0 15456 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_162
timestamp 1649977179
transform 1 0 16008 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_203
timestamp 1649977179
transform 1 0 19780 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_212
timestamp 1649977179
transform 1 0 20608 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_238
timestamp 1649977179
transform 1 0 23000 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_244
timestamp 1649977179
transform 1 0 23552 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_256
timestamp 1649977179
transform 1 0 24656 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_268
timestamp 1649977179
transform 1 0 25760 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_95
timestamp 1649977179
transform 1 0 9844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_107
timestamp 1649977179
transform 1 0 10948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_118
timestamp 1649977179
transform 1 0 11960 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_130
timestamp 1649977179
transform 1 0 13064 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_136
timestamp 1649977179
transform 1 0 13616 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_148
timestamp 1649977179
transform 1 0 14720 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_160
timestamp 1649977179
transform 1 0 15824 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_169
timestamp 1649977179
transform 1 0 16652 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_175
timestamp 1649977179
transform 1 0 17204 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_187
timestamp 1649977179
transform 1 0 18308 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_192
timestamp 1649977179
transform 1 0 18768 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_205
timestamp 1649977179
transform 1 0 19964 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_211
timestamp 1649977179
transform 1 0 20516 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_223
timestamp 1649977179
transform 1 0 21620 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_235
timestamp 1649977179
transform 1 0 22724 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_247
timestamp 1649977179
transform 1 0 23828 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_617
timestamp 1649977179
transform 1 0 57868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1649977179
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_126
timestamp 1649977179
transform 1 0 12696 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_138
timestamp 1649977179
transform 1 0 13800 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_150
timestamp 1649977179
transform 1 0 14904 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_159
timestamp 1649977179
transform 1 0 15732 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_161
timestamp 1649977179
transform 1 0 15916 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_173
timestamp 1649977179
transform 1 0 17020 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_185
timestamp 1649977179
transform 1 0 18124 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_193
timestamp 1649977179
transform 1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_621
timestamp 1649977179
transform 1 0 58236 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_621
timestamp 1649977179
transform 1 0 58236 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_603
timestamp 1649977179
transform 1 0 56580 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_617
timestamp 1649977179
transform 1 0 57868 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_621
timestamp 1649977179
transform 1 0 58236 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_617
timestamp 1649977179
transform 1 0 57868 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_621
timestamp 1649977179
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_621
timestamp 1649977179
transform 1 0 58236 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_621
timestamp 1649977179
transform 1 0 58236 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_460
timestamp 1649977179
transform 1 0 43424 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_466
timestamp 1649977179
transform 1 0 43976 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_474
timestamp 1649977179
transform 1 0 44712 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_617
timestamp 1649977179
transform 1 0 57868 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_621
timestamp 1649977179
transform 1 0 58236 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_617
timestamp 1649977179
transform 1 0 57868 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_621
timestamp 1649977179
transform 1 0 58236 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_621
timestamp 1649977179
transform 1 0 58236 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_621
timestamp 1649977179
transform 1 0 58236 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_143
timestamp 1649977179
transform 1 0 14260 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_151
timestamp 1649977179
transform 1 0 14996 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_154
timestamp 1649977179
transform 1 0 15272 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_166
timestamp 1649977179
transform 1 0 16376 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_169
timestamp 1649977179
transform 1 0 16652 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_173
timestamp 1649977179
transform 1 0 17020 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_176
timestamp 1649977179
transform 1 0 17296 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_180
timestamp 1649977179
transform 1 0 17664 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_183
timestamp 1649977179
transform 1 0 17940 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_187
timestamp 1649977179
transform 1 0 18308 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_190
timestamp 1649977179
transform 1 0 18584 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_98_199
timestamp 1649977179
transform 1 0 19412 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_207
timestamp 1649977179
transform 1 0 20148 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_212
timestamp 1649977179
transform 1 0 20608 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_98_219
timestamp 1649977179
transform 1 0 21252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_225
timestamp 1649977179
transform 1 0 21804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_228
timestamp 1649977179
transform 1 0 22080 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_240
timestamp 1649977179
transform 1 0 23184 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_285
timestamp 1649977179
transform 1 0 27324 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_291
timestamp 1649977179
transform 1 0 27876 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_98_297
timestamp 1649977179
transform 1 0 28428 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_305
timestamp 1649977179
transform 1 0 29164 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_313
timestamp 1649977179
transform 1 0 29900 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_316
timestamp 1649977179
transform 1 0 30176 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_328
timestamp 1649977179
transform 1 0 31280 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_340
timestamp 1649977179
transform 1 0 32384 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_352
timestamp 1649977179
transform 1 0 33488 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_451
timestamp 1649977179
transform 1 0 42596 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_454
timestamp 1649977179
transform 1 0 42872 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_458
timestamp 1649977179
transform 1 0 43240 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_461
timestamp 1649977179
transform 1 0 43516 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_465
timestamp 1649977179
transform 1 0 43884 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_468
timestamp 1649977179
transform 1 0 44160 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_98_479
timestamp 1649977179
transform 1 0 45172 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_493
timestamp 1649977179
transform 1 0 46460 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_496
timestamp 1649977179
transform 1 0 46736 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_508
timestamp 1649977179
transform 1 0 47840 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_520
timestamp 1649977179
transform 1 0 48944 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_140
timestamp 1649977179
transform 1 0 13984 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_148
timestamp 1649977179
transform 1 0 14720 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_152
timestamp 1649977179
transform 1 0 15088 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_158
timestamp 1649977179
transform 1 0 15640 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_99_162
timestamp 1649977179
transform 1 0 16008 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_172
timestamp 1649977179
transform 1 0 16928 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_179
timestamp 1649977179
transform 1 0 17572 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_186
timestamp 1649977179
transform 1 0 18216 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_200
timestamp 1649977179
transform 1 0 19504 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_210
timestamp 1649977179
transform 1 0 20424 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_218
timestamp 1649977179
transform 1 0 21160 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_99_231
timestamp 1649977179
transform 1 0 22356 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_242
timestamp 1649977179
transform 1 0 23368 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_248
timestamp 1649977179
transform 1 0 23920 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_260
timestamp 1649977179
transform 1 0 25024 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_272
timestamp 1649977179
transform 1 0 26128 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_284
timestamp 1649977179
transform 1 0 27232 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_291
timestamp 1649977179
transform 1 0 27876 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_298
timestamp 1649977179
transform 1 0 28520 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_304
timestamp 1649977179
transform 1 0 29072 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_308
timestamp 1649977179
transform 1 0 29440 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_319
timestamp 1649977179
transform 1 0 30452 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_325
timestamp 1649977179
transform 1 0 31004 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_332
timestamp 1649977179
transform 1 0 31648 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_340
timestamp 1649977179
transform 1 0 32384 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_346
timestamp 1649977179
transform 1 0 32936 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_352
timestamp 1649977179
transform 1 0 33488 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_356
timestamp 1649977179
transform 1 0 33856 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_362
timestamp 1649977179
transform 1 0 34408 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_99_374
timestamp 1649977179
transform 1 0 35512 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_380
timestamp 1649977179
transform 1 0 36064 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_386
timestamp 1649977179
transform 1 0 36616 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_453
timestamp 1649977179
transform 1 0 42780 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_457
timestamp 1649977179
transform 1 0 43148 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_464
timestamp 1649977179
transform 1 0 43792 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_471
timestamp 1649977179
transform 1 0 44436 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_478
timestamp 1649977179
transform 1 0 45080 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_492
timestamp 1649977179
transform 1 0 46368 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_499
timestamp 1649977179
transform 1 0 47012 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_621
timestamp 1649977179
transform 1 0 58236 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_161
timestamp 1649977179
transform 1 0 15916 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_164
timestamp 1649977179
transform 1 0 16192 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_176
timestamp 1649977179
transform 1 0 17296 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_188
timestamp 1649977179
transform 1 0 18400 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1649977179
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1649977179
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1649977179
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_277
timestamp 1649977179
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_289
timestamp 1649977179
transform 1 0 27692 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_295
timestamp 1649977179
transform 1 0 28244 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_307
timestamp 1649977179
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_311
timestamp 1649977179
transform 1 0 29716 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_323
timestamp 1649977179
transform 1 0 30820 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_335
timestamp 1649977179
transform 1 0 31924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_347
timestamp 1649977179
transform 1 0 33028 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_359
timestamp 1649977179
transform 1 0 34132 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_429
timestamp 1649977179
transform 1 0 40572 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_450
timestamp 1649977179
transform 1 0 42504 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_462
timestamp 1649977179
transform 1 0 43608 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_474
timestamp 1649977179
transform 1 0 44712 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_482
timestamp 1649977179
transform 1 0 45448 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_494
timestamp 1649977179
transform 1 0 46552 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_506
timestamp 1649977179
transform 1 0 47656 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_518
timestamp 1649977179
transform 1 0 48760 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_530
timestamp 1649977179
transform 1 0 49864 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_609
timestamp 1649977179
transform 1 0 57132 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_614
timestamp 1649977179
transform 1 0 57592 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1649977179
transform 1 0 58236 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_7
timestamp 1649977179
transform 1 0 1748 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_11
timestamp 1649977179
transform 1 0 2116 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_23
timestamp 1649977179
transform 1 0 3220 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1649977179
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_32
timestamp 1649977179
transform 1 0 4048 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_40
timestamp 1649977179
transform 1 0 4784 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_45
timestamp 1649977179
transform 1 0 5244 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_53
timestamp 1649977179
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_62
timestamp 1649977179
transform 1 0 6808 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_74
timestamp 1649977179
transform 1 0 7912 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_79
timestamp 1649977179
transform 1 0 8372 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_83
timestamp 1649977179
transform 1 0 8740 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_96
timestamp 1649977179
transform 1 0 9936 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_108
timestamp 1649977179
transform 1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_116
timestamp 1649977179
transform 1 0 11776 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_124
timestamp 1649977179
transform 1 0 12512 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_131
timestamp 1649977179
transform 1 0 13156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_139
timestamp 1649977179
transform 1 0 13892 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_148
timestamp 1649977179
transform 1 0 14720 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_160
timestamp 1649977179
transform 1 0 15824 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_173
timestamp 1649977179
transform 1 0 17020 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_177
timestamp 1649977179
transform 1 0 17388 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_182
timestamp 1649977179
transform 1 0 17848 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_194
timestamp 1649977179
transform 1 0 18952 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_201
timestamp 1649977179
transform 1 0 19596 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_209
timestamp 1649977179
transform 1 0 20332 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_216
timestamp 1649977179
transform 1 0 20976 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_233
timestamp 1649977179
transform 1 0 22540 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_245
timestamp 1649977179
transform 1 0 23644 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_251
timestamp 1649977179
transform 1 0 24196 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_257
timestamp 1649977179
transform 1 0 24748 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_267
timestamp 1649977179
transform 1 0 25668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1649977179
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_285
timestamp 1649977179
transform 1 0 27324 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_301
timestamp 1649977179
transform 1 0 28796 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_307
timestamp 1649977179
transform 1 0 29348 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_313
timestamp 1649977179
transform 1 0 29900 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_318
timestamp 1649977179
transform 1 0 30360 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_330
timestamp 1649977179
transform 1 0 31464 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_341
timestamp 1649977179
transform 1 0 32476 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_347
timestamp 1649977179
transform 1 0 33028 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_352
timestamp 1649977179
transform 1 0 33488 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_369
timestamp 1649977179
transform 1 0 35052 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_381
timestamp 1649977179
transform 1 0 36156 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_386
timestamp 1649977179
transform 1 0 36616 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_403
timestamp 1649977179
transform 1 0 38180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_415
timestamp 1649977179
transform 1 0 39284 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_419
timestamp 1649977179
transform 1 0 39652 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_425
timestamp 1649977179
transform 1 0 40204 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_101_437
timestamp 1649977179
transform 1 0 41308 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1649977179
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_454
timestamp 1649977179
transform 1 0 42872 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_466
timestamp 1649977179
transform 1 0 43976 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_471
timestamp 1649977179
transform 1 0 44436 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_475
timestamp 1649977179
transform 1 0 44804 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_477
timestamp 1649977179
transform 1 0 44988 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_483
timestamp 1649977179
transform 1 0 45540 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_488
timestamp 1649977179
transform 1 0 46000 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_500
timestamp 1649977179
transform 1 0 47104 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_509
timestamp 1649977179
transform 1 0 47932 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_517
timestamp 1649977179
transform 1 0 48668 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_522
timestamp 1649977179
transform 1 0 49128 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_530
timestamp 1649977179
transform 1 0 49864 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1649977179
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_539
timestamp 1649977179
transform 1 0 50692 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_551
timestamp 1649977179
transform 1 0 51796 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_556
timestamp 1649977179
transform 1 0 52256 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_573
timestamp 1649977179
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_585
timestamp 1649977179
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_593
timestamp 1649977179
transform 1 0 55660 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_599
timestamp 1649977179
transform 1 0 56212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_607
timestamp 1649977179
transform 1 0 56948 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_615
timestamp 1649977179
transform 1 0 57684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1649977179
transform 1 0 58236 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0855_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0856_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6440 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0857_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0858_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1649977179
transform -1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0862_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0863_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0864_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0865_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0866_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0867_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0868_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4692 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0869_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0870_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0871_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1649977179
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0874_
timestamp 1649977179
transform -1 0 2576 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 1649977179
transform 1 0 3772 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 1649977179
transform 1 0 2944 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp 1649977179
transform 1 0 4048 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1649977179
transform -1 0 2944 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1649977179
transform 1 0 4232 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1649977179
transform 1 0 5152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0888_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1649977179
transform -1 0 4784 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0892_
timestamp 1649977179
transform -1 0 3128 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1649977179
transform 1 0 9568 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1649977179
transform 1 0 2392 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0897_
timestamp 1649977179
transform -1 0 2576 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1649977179
transform 1 0 2392 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1649977179
transform -1 0 2576 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0905_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1649977179
transform -1 0 7176 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1649977179
transform -1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0909_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6624 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0910_
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0911_
timestamp 1649977179
transform 1 0 18216 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_4  _0912_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11408 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0913_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12052 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1649977179
transform -1 0 11960 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0915_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0916_
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1649977179
transform -1 0 11960 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1649977179
transform 1 0 7912 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0919_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4784 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1649977179
transform 1 0 6256 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0921_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0922_
timestamp 1649977179
transform -1 0 6808 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1649977179
transform -1 0 5060 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0924_
timestamp 1649977179
transform 1 0 2668 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0925_
timestamp 1649977179
transform -1 0 7360 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 1649977179
transform -1 0 4232 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0927_
timestamp 1649977179
transform 1 0 2668 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0928_
timestamp 1649977179
transform -1 0 8280 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1649977179
transform -1 0 6808 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0930_
timestamp 1649977179
transform 1 0 5152 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0931_
timestamp 1649977179
transform -1 0 10580 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1649977179
transform -1 0 6808 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0933_
timestamp 1649977179
transform -1 0 5888 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0934_
timestamp 1649977179
transform 1 0 23460 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0935_
timestamp 1649977179
transform 1 0 13156 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1649977179
transform -1 0 12696 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1649977179
transform -1 0 11960 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0938_
timestamp 1649977179
transform -1 0 13524 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0939_
timestamp 1649977179
transform 1 0 12328 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1649977179
transform -1 0 23920 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1649977179
transform 1 0 16192 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0942_
timestamp 1649977179
transform -1 0 15732 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1649977179
transform -1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 1649977179
transform 1 0 14260 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1649977179
transform -1 0 15824 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1649977179
transform -1 0 25668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0947_
timestamp 1649977179
transform 1 0 14536 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0948_
timestamp 1649977179
transform -1 0 15456 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0949_
timestamp 1649977179
transform -1 0 25300 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1649977179
transform 1 0 12236 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1649977179
transform 1 0 12328 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1649977179
transform -1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0953_
timestamp 1649977179
transform 1 0 12696 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1649977179
transform 1 0 13156 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0955_
timestamp 1649977179
transform 1 0 13064 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1649977179
transform -1 0 13800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1649977179
transform 1 0 13524 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1649977179
transform 1 0 12880 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0959_
timestamp 1649977179
transform -1 0 11040 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1649977179
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0961_
timestamp 1649977179
transform -1 0 30360 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0962_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 31188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0963_
timestamp 1649977179
transform -1 0 31004 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0964_
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0965_
timestamp 1649977179
transform 1 0 29992 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1649977179
transform 1 0 29992 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1649977179
transform -1 0 29992 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0968_
timestamp 1649977179
transform -1 0 29072 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1649977179
transform -1 0 28980 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0970_
timestamp 1649977179
transform 1 0 27416 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0971_
timestamp 1649977179
transform -1 0 28244 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0972_
timestamp 1649977179
transform 1 0 27232 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1649977179
transform 1 0 29532 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0974_
timestamp 1649977179
transform 1 0 12420 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0975_
timestamp 1649977179
transform -1 0 31280 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0976_
timestamp 1649977179
transform -1 0 30820 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1649977179
transform 1 0 31372 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1649977179
transform 1 0 30268 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0979_
timestamp 1649977179
transform 1 0 35512 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1649977179
transform -1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0981_
timestamp 1649977179
transform 1 0 35052 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0982_
timestamp 1649977179
transform -1 0 36708 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0983_
timestamp 1649977179
transform 1 0 35144 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0984_
timestamp 1649977179
transform -1 0 36616 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0985_
timestamp 1649977179
transform 1 0 35512 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0986_
timestamp 1649977179
transform -1 0 36524 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1649977179
transform 1 0 36064 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0988_
timestamp 1649977179
transform 1 0 28704 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0989_
timestamp 1649977179
transform -1 0 37536 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0990_
timestamp 1649977179
transform 1 0 35236 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0991_
timestamp 1649977179
transform -1 0 36800 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0992_
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0993_
timestamp 1649977179
transform -1 0 34960 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1649977179
transform 1 0 32292 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0995_
timestamp 1649977179
transform -1 0 33120 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _0996_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0998_
timestamp 1649977179
transform -1 0 30820 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1649977179
transform -1 0 31096 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1000_
timestamp 1649977179
transform -1 0 30728 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1649977179
transform 1 0 31372 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1002_
timestamp 1649977179
transform 1 0 32476 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1649977179
transform -1 0 28244 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 1649977179
transform 1 0 28244 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1649977179
transform -1 0 28428 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1006_
timestamp 1649977179
transform -1 0 31832 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1007_
timestamp 1649977179
transform 1 0 27140 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1649977179
transform -1 0 29072 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1649977179
transform 1 0 27508 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1649977179
transform -1 0 32568 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1649977179
transform 1 0 30452 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1649977179
transform -1 0 31556 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1013_
timestamp 1649977179
transform -1 0 31280 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1014_
timestamp 1649977179
transform 1 0 32384 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1649977179
transform -1 0 32384 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1649977179
transform 1 0 32660 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1649977179
transform -1 0 33120 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1649977179
transform 1 0 33672 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1019_
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1020_
timestamp 1649977179
transform -1 0 34224 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1649977179
transform 1 0 33120 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1649977179
transform -1 0 34684 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1649977179
transform 1 0 34684 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1024_
timestamp 1649977179
transform -1 0 35420 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1649977179
transform 1 0 33396 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1026_
timestamp 1649977179
transform -1 0 34224 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1649977179
transform 1 0 32108 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1028_
timestamp 1649977179
transform -1 0 32936 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1029_
timestamp 1649977179
transform 1 0 33764 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1030_
timestamp 1649977179
transform 1 0 29992 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1649977179
transform -1 0 31556 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1032_
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1649977179
transform -1 0 10488 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1034_
timestamp 1649977179
transform -1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1035_
timestamp 1649977179
transform 1 0 9200 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1036_
timestamp 1649977179
transform -1 0 8464 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1037_
timestamp 1649977179
transform 1 0 12328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1038_
timestamp 1649977179
transform 1 0 16744 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1039_
timestamp 1649977179
transform -1 0 10856 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1040_
timestamp 1649977179
transform -1 0 5888 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1041_
timestamp 1649977179
transform -1 0 5704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1649977179
transform -1 0 4784 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1649977179
transform 1 0 2576 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1649977179
transform -1 0 4784 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1649977179
transform -1 0 7636 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1047_
timestamp 1649977179
transform 1 0 6164 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1649977179
transform 1 0 6992 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1049_
timestamp 1649977179
transform 1 0 11776 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1050_
timestamp 1649977179
transform 1 0 23368 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1649977179
transform 1 0 18400 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1052_
timestamp 1649977179
transform 1 0 6992 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1053_
timestamp 1649977179
transform 1 0 16744 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_
timestamp 1649977179
transform 1 0 17480 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 1649977179
transform -1 0 20792 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1056_
timestamp 1649977179
transform -1 0 20700 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1649977179
transform 1 0 18308 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1058_
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1649977179
transform -1 0 20608 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1649977179
transform 1 0 19688 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 1649977179
transform -1 0 20424 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1649977179
transform -1 0 18768 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1064_
timestamp 1649977179
transform -1 0 19136 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1649977179
transform -1 0 18768 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1649977179
transform -1 0 16100 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1649977179
transform 1 0 14720 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1649977179
transform 1 0 15456 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1069_
timestamp 1649977179
transform -1 0 16100 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 1649977179
transform -1 0 18584 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1649977179
transform -1 0 18400 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1649977179
transform -1 0 16192 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1073_
timestamp 1649977179
transform -1 0 15732 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1074_
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1649977179
transform -1 0 11040 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1077_
timestamp 1649977179
transform 1 0 9476 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1649977179
transform -1 0 11224 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1649977179
transform 1 0 9568 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1649977179
transform 1 0 11684 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1081_
timestamp 1649977179
transform 1 0 23276 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1649977179
transform 1 0 11776 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1649977179
transform -1 0 15640 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1649977179
transform -1 0 13616 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1649977179
transform -1 0 15180 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1649977179
transform -1 0 24288 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1649977179
transform -1 0 26036 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1090_
timestamp 1649977179
transform 1 0 24472 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1649977179
transform -1 0 26680 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1093_
timestamp 1649977179
transform -1 0 25116 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp 1649977179
transform -1 0 25300 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1649977179
transform 1 0 24104 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1097_
timestamp 1649977179
transform -1 0 25392 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1649977179
transform -1 0 26496 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1649977179
transform -1 0 25944 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1649977179
transform 1 0 23644 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1649977179
transform -1 0 25300 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1649977179
transform 1 0 23368 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1103_
timestamp 1649977179
transform -1 0 24932 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1104_
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1105_
timestamp 1649977179
transform 1 0 21712 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1107_
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1649977179
transform -1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1109_
timestamp 1649977179
transform -1 0 25392 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1649977179
transform -1 0 23828 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1113_
timestamp 1649977179
transform -1 0 23920 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1649977179
transform 1 0 24380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1115_
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1649977179
transform -1 0 24380 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1649977179
transform -1 0 25116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1649977179
transform -1 0 24840 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1120_
timestamp 1649977179
transform 1 0 23184 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1121_
timestamp 1649977179
transform 1 0 18584 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1649977179
transform -1 0 26312 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1649977179
transform -1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1649977179
transform -1 0 26128 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1126_
timestamp 1649977179
transform -1 0 25944 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1649977179
transform 1 0 28520 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1128_
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1649977179
transform -1 0 28796 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1649977179
transform -1 0 31280 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1131_
timestamp 1649977179
transform 1 0 33120 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1649977179
transform -1 0 32936 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1649977179
transform 1 0 30084 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1134_
timestamp 1649977179
transform 1 0 30544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1649977179
transform 1 0 32292 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1649977179
transform -1 0 33212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1137_
timestamp 1649977179
transform 1 0 29900 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1649977179
transform -1 0 32568 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1139_
timestamp 1649977179
transform -1 0 31832 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1649977179
transform 1 0 27324 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1649977179
transform 1 0 31280 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1649977179
transform -1 0 32844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1143_
timestamp 1649977179
transform 1 0 27324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1649977179
transform 1 0 29532 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1145_
timestamp 1649977179
transform -1 0 31556 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1146_
timestamp 1649977179
transform 1 0 19780 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1649977179
transform -1 0 22724 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1148_
timestamp 1649977179
transform -1 0 27784 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1649977179
transform 1 0 22080 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1150_
timestamp 1649977179
transform 1 0 20516 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1151_
timestamp 1649977179
transform 1 0 24380 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1152_
timestamp 1649977179
transform 1 0 24932 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1649977179
transform -1 0 19780 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1156_
timestamp 1649977179
transform -1 0 21068 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1157_
timestamp 1649977179
transform 1 0 16100 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1158_
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1649977179
transform 1 0 19872 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1649977179
transform -1 0 13616 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1649977179
transform 1 0 15916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1166_
timestamp 1649977179
transform 1 0 14444 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1168_
timestamp 1649977179
transform 1 0 28152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1169_
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1170_
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1171_
timestamp 1649977179
transform 1 0 18584 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1172_
timestamp 1649977179
transform 1 0 22908 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1649977179
transform 1 0 28612 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1175_
timestamp 1649977179
transform 1 0 29072 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1649977179
transform 1 0 29808 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1177_
timestamp 1649977179
transform -1 0 31004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1178_
timestamp 1649977179
transform 1 0 28612 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1179_
timestamp 1649977179
transform 1 0 30360 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1649977179
transform -1 0 28704 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1181_
timestamp 1649977179
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1649977179
transform 1 0 27876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1649977179
transform -1 0 27324 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1184_
timestamp 1649977179
transform 1 0 25760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1649977179
transform -1 0 20240 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1186_
timestamp 1649977179
transform 1 0 20608 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1649977179
transform -1 0 22264 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1188_
timestamp 1649977179
transform 1 0 21160 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1189_
timestamp 1649977179
transform 1 0 7820 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1649977179
transform -1 0 22540 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1191_
timestamp 1649977179
transform -1 0 35696 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1192_
timestamp 1649977179
transform 1 0 36524 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1193_
timestamp 1649977179
transform -1 0 39652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1649977179
transform 1 0 36064 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1195_
timestamp 1649977179
transform -1 0 38640 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1649977179
transform -1 0 36616 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1649977179
transform 1 0 35052 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1649977179
transform 1 0 38640 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1199_
timestamp 1649977179
transform 1 0 34408 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1200_
timestamp 1649977179
transform 1 0 38456 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1649977179
transform -1 0 36432 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1202_
timestamp 1649977179
transform -1 0 36524 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1203_
timestamp 1649977179
transform 1 0 38364 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1204_
timestamp 1649977179
transform 1 0 38548 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1206_
timestamp 1649977179
transform 1 0 38640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1649977179
transform -1 0 40204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1208_
timestamp 1649977179
transform -1 0 39192 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1649977179
transform -1 0 37720 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1210_
timestamp 1649977179
transform 1 0 37720 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1649977179
transform 1 0 41032 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1212_
timestamp 1649977179
transform 1 0 33304 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1213_
timestamp 1649977179
transform 1 0 40664 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1649977179
transform 1 0 40112 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1215_
timestamp 1649977179
transform 1 0 40204 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1216_
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1217_
timestamp 1649977179
transform 1 0 40572 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1218_
timestamp 1649977179
transform 1 0 40296 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1649977179
transform 1 0 40388 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 1649977179
transform 1 0 40664 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1649977179
transform -1 0 37720 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1224_
timestamp 1649977179
transform -1 0 36064 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1649977179
transform -1 0 36800 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1226_
timestamp 1649977179
transform -1 0 22172 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1227_
timestamp 1649977179
transform -1 0 35512 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1228_
timestamp 1649977179
transform 1 0 35880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1229_
timestamp 1649977179
transform -1 0 37996 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1230_
timestamp 1649977179
transform 1 0 35144 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1231_
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1649977179
transform -1 0 35788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1649977179
transform 1 0 34960 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1649977179
transform -1 0 35420 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1235_
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1236_
timestamp 1649977179
transform -1 0 37352 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1237_
timestamp 1649977179
transform 1 0 34868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1238_
timestamp 1649977179
transform 1 0 36708 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1649977179
transform -1 0 38180 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1241_
timestamp 1649977179
transform -1 0 40020 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1242_
timestamp 1649977179
transform -1 0 39284 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1243_
timestamp 1649977179
transform 1 0 37628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1244_
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1246_
timestamp 1649977179
transform 1 0 37536 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1247_
timestamp 1649977179
transform 1 0 38916 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1248_
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1249_
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1250_
timestamp 1649977179
transform -1 0 41676 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1251_
timestamp 1649977179
transform 1 0 38180 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1252_
timestamp 1649977179
transform 1 0 38456 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1253_
timestamp 1649977179
transform 1 0 39928 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1254_
timestamp 1649977179
transform 1 0 40204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1255_
timestamp 1649977179
transform -1 0 41308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1649977179
transform 1 0 37352 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1257_
timestamp 1649977179
transform -1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1649977179
transform -1 0 36524 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1649977179
transform 1 0 35696 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1260_
timestamp 1649977179
transform -1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1261_
timestamp 1649977179
transform 1 0 23460 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1262_
timestamp 1649977179
transform -1 0 26496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1263_
timestamp 1649977179
transform 1 0 29900 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1649977179
transform -1 0 27416 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1649977179
transform -1 0 29072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1649977179
transform 1 0 27324 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1267_
timestamp 1649977179
transform 1 0 27232 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1268_
timestamp 1649977179
transform -1 0 27324 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1269_
timestamp 1649977179
transform 1 0 27048 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1270_
timestamp 1649977179
transform 1 0 28612 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1271_
timestamp 1649977179
transform -1 0 33672 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1272_
timestamp 1649977179
transform -1 0 30176 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1649977179
transform 1 0 29992 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1649977179
transform 1 0 29992 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1649977179
transform -1 0 29624 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1278_
timestamp 1649977179
transform -1 0 31280 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1649977179
transform 1 0 32660 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1280_
timestamp 1649977179
transform 1 0 33488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1281_
timestamp 1649977179
transform 1 0 33488 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1282_
timestamp 1649977179
transform -1 0 34132 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1649977179
transform -1 0 33212 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1284_
timestamp 1649977179
transform 1 0 15548 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1649977179
transform 1 0 24288 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1286_
timestamp 1649977179
transform -1 0 33488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1287_
timestamp 1649977179
transform -1 0 33396 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1288_
timestamp 1649977179
transform -1 0 33304 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1649977179
transform 1 0 31924 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1290_
timestamp 1649977179
transform -1 0 33120 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1649977179
transform 1 0 26312 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1292_
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1649977179
transform -1 0 26220 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1294_
timestamp 1649977179
transform 1 0 25668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1295_
timestamp 1649977179
transform 1 0 5428 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1296_
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 1649977179
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1298_
timestamp 1649977179
transform -1 0 17112 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _1299_
timestamp 1649977179
transform -1 0 12052 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1300_
timestamp 1649977179
transform -1 0 7728 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1649977179
transform -1 0 15824 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1649977179
transform 1 0 8372 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1303_
timestamp 1649977179
transform -1 0 4692 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1304_
timestamp 1649977179
transform -1 0 7728 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1305_
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1306_
timestamp 1649977179
transform 1 0 5244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1307_
timestamp 1649977179
transform -1 0 2024 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1308_
timestamp 1649977179
transform 1 0 2300 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1309_
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1649977179
transform 1 0 2208 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1649977179
transform 1 0 2116 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1312_
timestamp 1649977179
transform 1 0 6900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1649977179
transform -1 0 7728 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1314_
timestamp 1649977179
transform -1 0 5888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1315_
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1649977179
transform 1 0 5428 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1317_
timestamp 1649977179
transform -1 0 6900 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1318_
timestamp 1649977179
transform 1 0 21896 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1319_
timestamp 1649977179
transform 1 0 20884 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1649977179
transform -1 0 21160 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1649977179
transform 1 0 20884 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1322_
timestamp 1649977179
transform -1 0 22448 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1649977179
transform 1 0 21344 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1324_
timestamp 1649977179
transform 1 0 25668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1649977179
transform 1 0 22540 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1326_
timestamp 1649977179
transform -1 0 23184 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1327_
timestamp 1649977179
transform -1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1649977179
transform 1 0 22448 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1329_
timestamp 1649977179
transform -1 0 23276 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1330_
timestamp 1649977179
transform 1 0 17020 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1649977179
transform 1 0 23000 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1332_
timestamp 1649977179
transform 1 0 21896 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1333_
timestamp 1649977179
transform 1 0 17020 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1649977179
transform -1 0 23184 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1335_
timestamp 1649977179
transform 1 0 21620 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1336_
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1649977179
transform 1 0 18308 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1649977179
transform 1 0 18492 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1339_
timestamp 1649977179
transform 1 0 18032 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1340_
timestamp 1649977179
transform 1 0 9384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1649977179
transform 1 0 19872 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1649977179
transform 1 0 19780 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_4  _1343_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1649977179
transform -1 0 22816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1345_
timestamp 1649977179
transform -1 0 23092 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1649977179
transform -1 0 21988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1347_
timestamp 1649977179
transform -1 0 21344 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1348_
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1349_
timestamp 1649977179
transform 1 0 21988 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1649977179
transform 1 0 22632 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1351_
timestamp 1649977179
transform -1 0 17848 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1352_
timestamp 1649977179
transform 1 0 16836 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1649977179
transform -1 0 19688 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1649977179
transform 1 0 18492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1649977179
transform -1 0 18400 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1356_
timestamp 1649977179
transform 1 0 16836 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp 1649977179
transform -1 0 18492 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1358_
timestamp 1649977179
transform 1 0 17664 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1359_
timestamp 1649977179
transform 1 0 17480 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1649977179
transform -1 0 22264 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1361_
timestamp 1649977179
transform -1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1649977179
transform -1 0 25300 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1649977179
transform -1 0 25116 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1365_
timestamp 1649977179
transform -1 0 25668 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1649977179
transform -1 0 26220 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1367_
timestamp 1649977179
transform -1 0 25300 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1649977179
transform 1 0 27508 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1369_
timestamp 1649977179
transform -1 0 26312 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1649977179
transform -1 0 26220 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1371_
timestamp 1649977179
transform 1 0 11868 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1372_
timestamp 1649977179
transform -1 0 11684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1373_
timestamp 1649977179
transform -1 0 25760 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1649977179
transform -1 0 27416 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1375_
timestamp 1649977179
transform -1 0 26220 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1649977179
transform -1 0 25024 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1377_
timestamp 1649977179
transform -1 0 23092 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 1649977179
transform -1 0 23920 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1379_
timestamp 1649977179
transform -1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1649977179
transform 1 0 10028 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1382_
timestamp 1649977179
transform -1 0 9200 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1383_
timestamp 1649977179
transform -1 0 7820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1384_
timestamp 1649977179
transform 1 0 10672 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1385_
timestamp 1649977179
transform -1 0 12512 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1386_
timestamp 1649977179
transform -1 0 10028 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1387_
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1388_
timestamp 1649977179
transform 1 0 7268 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1649977179
transform -1 0 4232 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1390_
timestamp 1649977179
transform -1 0 10948 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1391_
timestamp 1649977179
transform 1 0 2576 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1649977179
transform -1 0 3588 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1393_
timestamp 1649977179
transform 1 0 2576 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1649977179
transform 1 0 5428 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1395_
timestamp 1649977179
transform -1 0 6808 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1649977179
transform -1 0 9200 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1397_
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1398_
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1399_
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1649977179
transform 1 0 14352 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1649977179
transform -1 0 17112 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1403_
timestamp 1649977179
transform 1 0 12052 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1404_
timestamp 1649977179
transform 1 0 15456 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1649977179
transform 1 0 17664 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1406_
timestamp 1649977179
transform -1 0 18124 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1649977179
transform -1 0 17756 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1408_
timestamp 1649977179
transform 1 0 16928 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1649977179
transform -1 0 17204 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1410_
timestamp 1649977179
transform 1 0 15640 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1411_
timestamp 1649977179
transform -1 0 14168 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1412_
timestamp 1649977179
transform -1 0 13616 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1649977179
transform -1 0 11960 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1649977179
transform 1 0 10120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1415_
timestamp 1649977179
transform -1 0 10856 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1416_
timestamp 1649977179
transform -1 0 9936 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1417_
timestamp 1649977179
transform 1 0 9568 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1418_
timestamp 1649977179
transform -1 0 9568 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1419_
timestamp 1649977179
transform -1 0 8464 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1420_
timestamp 1649977179
transform -1 0 9384 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1421_
timestamp 1649977179
transform 1 0 8004 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1649977179
transform -1 0 4232 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1423_
timestamp 1649977179
transform 1 0 2760 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1424_
timestamp 1649977179
transform -1 0 3036 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1425_
timestamp 1649977179
transform 1 0 2208 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1649977179
transform -1 0 3680 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1427_
timestamp 1649977179
transform 1 0 2116 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1428_
timestamp 1649977179
transform 1 0 4784 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1429_
timestamp 1649977179
transform 1 0 4692 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1649977179
transform 1 0 7360 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1431_
timestamp 1649977179
transform -1 0 10856 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1433_
timestamp 1649977179
transform 1 0 9568 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1434_
timestamp 1649977179
transform -1 0 9660 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1435_
timestamp 1649977179
transform -1 0 9568 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1436_
timestamp 1649977179
transform 1 0 8924 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1649977179
transform -1 0 11224 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1438_
timestamp 1649977179
transform 1 0 9752 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1649977179
transform -1 0 10488 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1440_
timestamp 1649977179
transform 1 0 9660 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1441_
timestamp 1649977179
transform -1 0 11960 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1442_
timestamp 1649977179
transform -1 0 10028 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1443_
timestamp 1649977179
transform 1 0 12328 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1444_
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1445_
timestamp 1649977179
transform -1 0 11316 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1446_
timestamp 1649977179
transform 1 0 10304 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1649977179
transform 1 0 10396 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1448_
timestamp 1649977179
transform 1 0 9844 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1649977179
transform 1 0 8188 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1450_
timestamp 1649977179
transform 1 0 9016 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1451_
timestamp 1649977179
transform -1 0 14536 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1452_
timestamp 1649977179
transform 1 0 14444 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1453_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1454_
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1455_
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1456_
timestamp 1649977179
transform 1 0 15456 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 1649977179
transform -1 0 13064 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 1649977179
transform 1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1649977179
transform -1 0 11960 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1461_
timestamp 1649977179
transform 1 0 10396 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1649977179
transform -1 0 12788 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1463_
timestamp 1649977179
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1464_
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1465_
timestamp 1649977179
transform -1 0 14536 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1466_
timestamp 1649977179
transform -1 0 13616 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1467_
timestamp 1649977179
transform 1 0 12696 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1468_
timestamp 1649977179
transform 1 0 12420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1469_
timestamp 1649977179
transform -1 0 18124 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1649977179
transform -1 0 18768 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1471_
timestamp 1649977179
transform -1 0 19688 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1472_
timestamp 1649977179
transform -1 0 18676 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1473_
timestamp 1649977179
transform 1 0 18492 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1474_
timestamp 1649977179
transform -1 0 19964 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1475_
timestamp 1649977179
transform -1 0 21344 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1476_
timestamp 1649977179
transform -1 0 20884 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1477_
timestamp 1649977179
transform -1 0 21160 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1649977179
transform 1 0 22632 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1479_
timestamp 1649977179
transform -1 0 22264 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 1649977179
transform -1 0 19780 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1481_
timestamp 1649977179
transform 1 0 17296 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1649977179
transform -1 0 17572 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1483_
timestamp 1649977179
transform 1 0 16744 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1649977179
transform 1 0 17020 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1485_
timestamp 1649977179
transform -1 0 18584 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1486_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1487_
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1488_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1649977179
transform -1 0 21252 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1490_
timestamp 1649977179
transform 1 0 18032 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1649977179
transform 1 0 20884 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1649977179
transform 1 0 19320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1649977179
transform -1 0 17112 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1495_
timestamp 1649977179
transform 1 0 15364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1496_
timestamp 1649977179
transform -1 0 16284 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1497_
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 1649977179
transform -1 0 16192 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1499_
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1649977179
transform -1 0 19780 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1649977179
transform -1 0 18952 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1649977179
transform -1 0 19688 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1649977179
transform -1 0 18768 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1504_
timestamp 1649977179
transform 1 0 25760 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1505_
timestamp 1649977179
transform -1 0 27232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1649977179
transform -1 0 30820 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1507_
timestamp 1649977179
transform 1 0 25576 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1508_
timestamp 1649977179
transform -1 0 30452 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1649977179
transform -1 0 31280 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1510_
timestamp 1649977179
transform -1 0 30912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 1649977179
transform 1 0 31188 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1512_
timestamp 1649977179
transform -1 0 30820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1513_
timestamp 1649977179
transform -1 0 27784 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1514_
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1515_
timestamp 1649977179
transform -1 0 28520 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1516_
timestamp 1649977179
transform 1 0 27508 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1517_
timestamp 1649977179
transform -1 0 19688 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1518_
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1519_
timestamp 1649977179
transform 1 0 17296 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 1649977179
transform -1 0 19964 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1521_
timestamp 1649977179
transform -1 0 19136 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1522_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1523_
timestamp 1649977179
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1524_
timestamp 1649977179
transform -1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1525_
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1526_
timestamp 1649977179
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1527_
timestamp 1649977179
transform -1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1528_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_2  _1529_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1530_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1531_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35788 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1649977179
transform 1 0 23000 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1649977179
transform 1 0 22632 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1534_
timestamp 1649977179
transform -1 0 30544 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1535_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1536_
timestamp 1649977179
transform 1 0 4692 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1537_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1538_
timestamp 1649977179
transform 1 0 9844 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1539_
timestamp 1649977179
transform -1 0 11316 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1540_
timestamp 1649977179
transform -1 0 10212 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1541_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7360 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1542_
timestamp 1649977179
transform -1 0 35604 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1649977179
transform 1 0 23092 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 1649977179
transform -1 0 28336 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1546_
timestamp 1649977179
transform -1 0 24472 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1649977179
transform 1 0 4508 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1548_
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1549_
timestamp 1649977179
transform 1 0 9844 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1550_
timestamp 1649977179
transform -1 0 11040 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1649977179
transform 1 0 7084 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1552_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1553_
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1554_
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1555_
timestamp 1649977179
transform -1 0 36616 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1556_
timestamp 1649977179
transform 1 0 21988 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1557_
timestamp 1649977179
transform 1 0 22356 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1558_
timestamp 1649977179
transform -1 0 29348 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1559_
timestamp 1649977179
transform -1 0 23552 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1560_
timestamp 1649977179
transform 1 0 4324 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1561_
timestamp 1649977179
transform 1 0 4784 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1649977179
transform 1 0 11408 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1563_
timestamp 1649977179
transform 1 0 12420 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1564_
timestamp 1649977179
transform -1 0 8188 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1565_
timestamp 1649977179
transform -1 0 5888 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1566_
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1567_
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1568_
timestamp 1649977179
transform 1 0 35512 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1569_
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1570_
timestamp 1649977179
transform 1 0 35328 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1571_
timestamp 1649977179
transform 1 0 35972 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1649977179
transform -1 0 36524 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1573_
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1574_
timestamp 1649977179
transform 1 0 29808 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1649977179
transform 1 0 22724 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1576_
timestamp 1649977179
transform 1 0 29624 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1649977179
transform 1 0 29624 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1578_
timestamp 1649977179
transform 1 0 21896 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1649977179
transform 1 0 28244 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1580_
timestamp 1649977179
transform 1 0 21896 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1581_
timestamp 1649977179
transform 1 0 28152 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1649977179
transform 1 0 27140 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1583_
timestamp 1649977179
transform 1 0 31004 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1584_
timestamp 1649977179
transform -1 0 33856 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1585_
timestamp 1649977179
transform -1 0 31648 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1586_
timestamp 1649977179
transform -1 0 33764 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1587_
timestamp 1649977179
transform -1 0 31464 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1588_
timestamp 1649977179
transform -1 0 31188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1589_
timestamp 1649977179
transform 1 0 12052 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1590_
timestamp 1649977179
transform -1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1591_
timestamp 1649977179
transform 1 0 10856 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1592_
timestamp 1649977179
transform 1 0 12420 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1593_
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1594_
timestamp 1649977179
transform 1 0 6900 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1595_
timestamp 1649977179
transform 1 0 19688 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1596_
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1597_
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1598_
timestamp 1649977179
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1599_
timestamp 1649977179
transform -1 0 14812 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1600_
timestamp 1649977179
transform -1 0 14628 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1601_
timestamp 1649977179
transform -1 0 8464 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1602_
timestamp 1649977179
transform 1 0 4692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1603_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1604_
timestamp 1649977179
transform -1 0 7636 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1649977179
transform -1 0 36432 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1606_
timestamp 1649977179
transform 1 0 28612 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1649977179
transform 1 0 27600 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 1649977179
transform -1 0 31372 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1609_
timestamp 1649977179
transform -1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1610_
timestamp 1649977179
transform -1 0 15456 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1611_
timestamp 1649977179
transform -1 0 12880 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1612_
timestamp 1649977179
transform 1 0 7820 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1613_
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1614_
timestamp 1649977179
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1615_
timestamp 1649977179
transform -1 0 15916 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1616_
timestamp 1649977179
transform 1 0 14812 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1617_
timestamp 1649977179
transform 1 0 15272 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1618_
timestamp 1649977179
transform -1 0 9384 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1619_
timestamp 1649977179
transform 1 0 4968 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1620_
timestamp 1649977179
transform -1 0 8188 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1621_
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1622_
timestamp 1649977179
transform -1 0 36248 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1624_
timestamp 1649977179
transform 1 0 31004 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1649977179
transform -1 0 33580 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1626_
timestamp 1649977179
transform -1 0 33028 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1627_
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1628_
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1649977179
transform -1 0 22632 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1649977179
transform -1 0 21988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1631_
timestamp 1649977179
transform -1 0 21252 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1632_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1633_
timestamp 1649977179
transform -1 0 8372 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1634_
timestamp 1649977179
transform -1 0 35512 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1649977179
transform 1 0 32752 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp 1649977179
transform 1 0 32200 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1637_
timestamp 1649977179
transform -1 0 34040 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1638_
timestamp 1649977179
transform 1 0 33856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1639_
timestamp 1649977179
transform 1 0 13800 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp 1649977179
transform 1 0 17572 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1641_
timestamp 1649977179
transform -1 0 23092 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1642_
timestamp 1649977179
transform -1 0 22264 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1643_
timestamp 1649977179
transform -1 0 20240 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1644_
timestamp 1649977179
transform 1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1645_
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1646_
timestamp 1649977179
transform -1 0 10120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1647_
timestamp 1649977179
transform -1 0 36248 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 1649977179
transform 1 0 31004 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1649977179
transform 1 0 32108 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1650_
timestamp 1649977179
transform 1 0 32384 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1651_
timestamp 1649977179
transform 1 0 33396 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1652_
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1653_
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1649977179
transform -1 0 23368 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1655_
timestamp 1649977179
transform -1 0 23000 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1656_
timestamp 1649977179
transform -1 0 21252 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1657_
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1658_
timestamp 1649977179
transform -1 0 13340 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1659_
timestamp 1649977179
transform -1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1649977179
transform -1 0 37904 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1649977179
transform 1 0 29256 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1663_
timestamp 1649977179
transform -1 0 35328 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1664_
timestamp 1649977179
transform -1 0 30084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1665_
timestamp 1649977179
transform 1 0 12972 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1666_
timestamp 1649977179
transform 1 0 18768 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1667_
timestamp 1649977179
transform -1 0 22816 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1668_
timestamp 1649977179
transform 1 0 22356 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1669_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23184 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1670_
timestamp 1649977179
transform 1 0 10304 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1671_
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1649977179
transform -1 0 37904 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1673_
timestamp 1649977179
transform 1 0 28428 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1674_
timestamp 1649977179
transform 1 0 28336 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1649977179
transform -1 0 34592 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1676_
timestamp 1649977179
transform -1 0 30820 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 1649977179
transform 1 0 12236 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1678_
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1679_
timestamp 1649977179
transform -1 0 22816 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1680_
timestamp 1649977179
transform -1 0 19964 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1681_
timestamp 1649977179
transform -1 0 18400 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1682_
timestamp 1649977179
transform -1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1683_
timestamp 1649977179
transform -1 0 12880 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1684_
timestamp 1649977179
transform -1 0 37904 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1685_
timestamp 1649977179
transform 1 0 24564 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1686_
timestamp 1649977179
transform 1 0 23092 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1687_
timestamp 1649977179
transform -1 0 33948 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1688_
timestamp 1649977179
transform -1 0 26128 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1689_
timestamp 1649977179
transform 1 0 12052 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1690_
timestamp 1649977179
transform 1 0 14536 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1691_
timestamp 1649977179
transform 1 0 19688 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1692_
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1693_
timestamp 1649977179
transform -1 0 15732 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1694_
timestamp 1649977179
transform -1 0 4692 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1695_
timestamp 1649977179
transform -1 0 4600 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1696_
timestamp 1649977179
transform -1 0 37444 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1697_
timestamp 1649977179
transform 1 0 25208 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1698_
timestamp 1649977179
transform 1 0 25208 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1699_
timestamp 1649977179
transform -1 0 32936 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1700_
timestamp 1649977179
transform -1 0 27508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1701_
timestamp 1649977179
transform 1 0 12512 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1702_
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1703_
timestamp 1649977179
transform -1 0 21712 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1704_
timestamp 1649977179
transform -1 0 20608 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1705_
timestamp 1649977179
transform -1 0 15364 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1706_
timestamp 1649977179
transform 1 0 7728 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1707_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1708_
timestamp 1649977179
transform -1 0 4416 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1709_
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1710_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1649977179
transform 1 0 2668 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1649977179
transform 1 0 2576 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1649977179
transform 1 0 1932 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1649977179
transform 1 0 3404 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1649977179
transform 1 0 6440 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1649977179
transform 1 0 1840 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1649977179
transform 1 0 1840 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1649977179
transform 1 0 4416 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1649977179
transform 1 0 6072 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1649977179
transform -1 0 12696 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1649977179
transform 1 0 15364 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1649977179
transform -1 0 16928 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1649977179
transform -1 0 16192 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1649977179
transform -1 0 13340 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1649977179
transform 1 0 12144 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1649977179
transform 1 0 29072 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1649977179
transform 1 0 27324 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1649977179
transform 1 0 27140 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1649977179
transform -1 0 32108 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1649977179
transform 1 0 29808 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1649977179
transform 1 0 37444 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1649977179
transform 1 0 37996 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1649977179
transform 1 0 37904 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1649977179
transform -1 0 39560 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1649977179
transform -1 0 38732 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1649977179
transform -1 0 36156 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1649977179
transform -1 0 34224 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1649977179
transform 1 0 27232 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1649977179
transform 1 0 27140 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1649977179
transform 1 0 30176 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1649977179
transform 1 0 31004 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1649977179
transform 1 0 32660 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1649977179
transform -1 0 36156 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1649977179
transform -1 0 36248 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1649977179
transform -1 0 36800 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1649977179
transform -1 0 36156 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1649977179
transform -1 0 34040 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1649977179
transform 1 0 31924 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1649977179
transform 1 0 5336 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1649977179
transform 1 0 6072 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1649977179
transform -1 0 21896 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1649977179
transform -1 0 19780 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1649977179
transform -1 0 21344 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1649977179
transform 1 0 14720 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1649977179
transform -1 0 16652 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1649977179
transform 1 0 10948 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1649977179
transform 1 0 13156 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1649977179
transform 1 0 14168 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1649977179
transform 1 0 24196 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1649977179
transform -1 0 25668 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1649977179
transform -1 0 26404 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1649977179
transform 1 0 25668 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1649977179
transform -1 0 27140 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1649977179
transform -1 0 26680 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1649977179
transform -1 0 24012 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1649977179
transform -1 0 25852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1649977179
transform -1 0 23920 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1649977179
transform 1 0 25668 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1649977179
transform 1 0 25944 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1649977179
transform 1 0 30176 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1649977179
transform -1 0 34776 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1649977179
transform -1 0 33672 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1649977179
transform -1 0 33948 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1649977179
transform -1 0 31648 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1649977179
transform 1 0 21528 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1649977179
transform 1 0 24840 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1649977179
transform -1 0 15180 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1649977179
transform -1 0 18492 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1649977179
transform -1 0 18216 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1649977179
transform 1 0 28520 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1649977179
transform -1 0 32844 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1649977179
transform -1 0 31004 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1649977179
transform 1 0 27600 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1649977179
transform -1 0 26496 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1649977179
transform -1 0 21344 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1649977179
transform 1 0 21344 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1649977179
transform 1 0 34868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1649977179
transform 1 0 38272 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1649977179
transform -1 0 38732 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1649977179
transform 1 0 38732 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1649977179
transform -1 0 37352 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1649977179
transform -1 0 40204 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1649977179
transform -1 0 40204 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1649977179
transform 1 0 38732 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1649977179
transform 1 0 38824 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1649977179
transform 1 0 38824 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1649977179
transform 1 0 36800 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1649977179
transform 1 0 34960 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1649977179
transform 1 0 34592 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1649977179
transform 1 0 34684 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1649977179
transform 1 0 37904 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1649977179
transform 1 0 38640 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1649977179
transform -1 0 37168 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1649977179
transform -1 0 40020 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1649977179
transform -1 0 40020 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1649977179
transform -1 0 39008 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1649977179
transform 1 0 38732 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1649977179
transform 1 0 38824 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1649977179
transform 1 0 35328 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1649977179
transform 1 0 26956 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1649977179
transform -1 0 26588 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1649977179
transform -1 0 31004 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1649977179
transform -1 0 31464 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1649977179
transform -1 0 31004 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1649977179
transform -1 0 34224 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1649977179
transform -1 0 34408 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1649977179
transform -1 0 34224 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1649977179
transform -1 0 35144 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1649977179
transform -1 0 34132 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1649977179
transform -1 0 28060 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1649977179
transform 1 0 24472 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1649977179
transform 1 0 2392 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1649977179
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1649977179
transform 1 0 6532 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1649977179
transform 1 0 20700 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1649977179
transform -1 0 25024 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1649977179
transform -1 0 23920 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1649977179
transform 1 0 21528 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1649977179
transform 1 0 17940 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1649977179
transform 1 0 18032 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1649977179
transform 1 0 20792 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1649977179
transform 1 0 25668 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1649977179
transform -1 0 29624 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1649977179
transform 1 0 25852 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1649977179
transform 1 0 22724 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1649977179
transform 1 0 23000 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1649977179
transform -1 0 7820 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1649977179
transform 1 0 2576 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1649977179
transform 1 0 2576 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1649977179
transform 1 0 6348 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1649977179
transform 1 0 6900 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1649977179
transform 1 0 13524 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1649977179
transform 1 0 15272 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1649977179
transform 1 0 18124 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1649977179
transform 1 0 17112 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1649977179
transform 1 0 15548 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1649977179
transform 1 0 13248 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1649977179
transform 1 0 10488 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1649977179
transform 1 0 2576 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1649977179
transform 1 0 2392 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1649977179
transform 1 0 1840 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1649977179
transform 1 0 7176 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1649977179
transform 1 0 9108 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1649977179
transform 1 0 8924 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1649977179
transform 1 0 10396 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1649977179
transform 1 0 9568 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1649977179
transform 1 0 9568 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1649977179
transform 1 0 9200 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1649977179
transform 1 0 11684 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1649977179
transform 1 0 19044 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1649977179
transform -1 0 20516 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1649977179
transform 1 0 22172 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1649977179
transform 1 0 16652 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1649977179
transform 1 0 16376 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1649977179
transform 1 0 17940 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1649977179
transform 1 0 29992 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1649977179
transform 1 0 30912 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1649977179
transform 1 0 31004 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1649977179
transform -1 0 29072 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1649977179
transform -1 0 5244 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1649977179
transform -1 0 9200 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1649977179
transform -1 0 8372 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1649977179
transform 1 0 6624 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1649977179
transform -1 0 8464 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1649977179
transform -1 0 8464 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1649977179
transform 1 0 9476 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1649977179
transform 1 0 11316 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1649977179
transform -1 0 13156 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1649977179
transform 1 0 1840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1649977179
transform 1 0 2392 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2167_
timestamp 1649977179
transform -1 0 43148 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2168_
timestamp 1649977179
transform -1 0 45080 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2169_
timestamp 1649977179
transform -1 0 44436 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2170_
timestamp 1649977179
transform -1 0 22356 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2171_
timestamp 1649977179
transform 1 0 20792 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _2172_
timestamp 1649977179
transform -1 0 29440 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2173_
timestamp 1649977179
transform -1 0 43792 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2174_
timestamp 1649977179
transform -1 0 46368 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2175_
timestamp 1649977179
transform -1 0 45724 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2176_
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2177_
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2178_
timestamp 1649977179
transform -1 0 16008 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2179_
timestamp 1649977179
transform -1 0 16928 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2180_
timestamp 1649977179
transform -1 0 17572 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2181_
timestamp 1649977179
transform -1 0 18860 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2182_
timestamp 1649977179
transform -1 0 21252 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2183_
timestamp 1649977179
transform -1 0 23368 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2184_
timestamp 1649977179
transform -1 0 18216 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2185_
timestamp 1649977179
transform -1 0 19504 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2186_
timestamp 1649977179
transform -1 0 27876 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2187_
timestamp 1649977179
transform -1 0 28520 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2188_
timestamp 1649977179
transform -1 0 30452 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2189_
timestamp 1649977179
transform -1 0 32384 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2190_
timestamp 1649977179
transform -1 0 33856 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2191_
timestamp 1649977179
transform -1 0 31648 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2192_
timestamp 1649977179
transform -1 0 36064 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2193_
timestamp 1649977179
transform -1 0 27876 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2194_
timestamp 1649977179
transform -1 0 47012 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2195_
timestamp 1649977179
transform -1 0 43424 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2196_
timestamp 1649977179
transform -1 0 56580 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20976 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1649977179
transform -1 0 12236 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1649977179
transform 1 0 16008 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1649977179
transform 1 0 9292 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1649977179
transform -1 0 5980 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1649977179
transform 1 0 5244 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1649977179
transform 1 0 11776 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1649977179
transform 1 0 17940 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1649977179
transform 1 0 16928 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1649977179
transform -1 0 22908 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1649977179
transform -1 0 28888 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1649977179
transform 1 0 23736 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1649977179
transform 1 0 28244 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1649977179
transform -1 0 34316 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1649977179
transform 1 0 38732 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1649977179
transform -1 0 33856 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1649977179
transform -1 0 28612 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1649977179
transform 1 0 25668 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1649977179
transform -1 0 32936 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1649977179
transform 1 0 37536 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1649977179
transform 1 0 36156 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1649977179
transform 1 0 37536 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1649977179
transform 1 0 32384 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1649977179
transform -1 0 31188 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1649977179
transform -1 0 26496 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1649977179
transform 1 0 24748 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1649977179
transform 1 0 18216 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1649977179
transform 1 0 17020 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1649977179
transform 1 0 17020 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1649977179
transform 1 0 10120 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1649977179
transform -1 0 5060 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_32_wb_clk_i
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_33_wb_clk_i
timestamp 1649977179
transform 1 0 3772 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1649977179
transform -1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1649977179
transform -1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1649977179
transform -1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1649977179
transform -1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1649977179
transform -1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1649977179
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform 1 0 19504 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform -1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform -1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1649977179
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input14
timestamp 1649977179
transform -1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1649977179
transform 1 0 21712 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1649977179
transform -1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1649977179
transform 1 0 22080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1649977179
transform -1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1649977179
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1649977179
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform 1 0 23368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 4600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 13616 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 7360 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 7912 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1649977179
transform -1 0 9292 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1649977179
transform -1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform 1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input49
timestamp 1649977179
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input53
timestamp 1649977179
transform 1 0 7912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input54
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1649977179
transform 1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 6716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform -1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 53452 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 50324 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 55292 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 40940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 42504 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform 1 0 44068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 45632 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 48760 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 13156 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 14720 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 16652 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 17480 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 19228 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 20608 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 22172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 24380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 25300 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 28428 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 29992 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 33120 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 36248 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 37812 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 39836 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 51888 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 56580 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 10672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 5060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8372 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform -1 0 9936 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform -1 0 11776 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform -1 0 5244 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform -1 0 6808 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform -1 0 2116 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform -1 0 4048 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform 1 0 57960 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform 1 0 57960 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform 1 0 57316 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform 1 0 57960 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform -1 0 51428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform -1 0 52440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform -1 0 52072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform -1 0 53728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform -1 0 52992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform -1 0 52440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform -1 0 53084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform -1 0 54372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform -1 0 53636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform -1 0 53728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform -1 0 54280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform -1 0 54924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform -1 0 54372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform -1 0 55568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform -1 0 54004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform -1 0 54648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform -1 0 55568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform -1 0 56212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform -1 0 55292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform -1 0 56212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform 1 0 57960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform 1 0 57316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform 1 0 57960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform 1 0 57960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform 1 0 57960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform 1 0 57960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform 1 0 57960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform 1 0 57960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform 1 0 57960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform 1 0 57960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform 1 0 57960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform 1 0 57960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 57960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform 1 0 57960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform 1 0 57960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform 1 0 57960 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform 1 0 57960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 57960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform 1 0 57960 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform 1 0 57960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform 1 0 57960 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform 1 0 57960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform 1 0 57960 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 57960 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform 1 0 57960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform 1 0 57960 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform 1 0 57960 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform 1 0 57960 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 57960 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform 1 0 57960 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform 1 0 57960 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform 1 0 57960 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform 1 0 57960 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform 1 0 57960 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform 1 0 57960 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform 1 0 57960 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform 1 0 57960 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform 1 0 57960 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform -1 0 51796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform 1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform -1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform 1 0 15272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform 1 0 17572 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform -1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 25116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform -1 0 25944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform -1 0 27048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform -1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform 1 0 29348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform 1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform -1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform -1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform -1 0 33672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform -1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform -1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform -1 0 34960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform -1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform -1 0 35052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform -1 0 35696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform -1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform -1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform -1 0 36984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform -1 0 37812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform -1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_278
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_279
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_280
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_281
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_282
timestamp 1649977179
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_283
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_284
timestamp 1649977179
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_285
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_286
timestamp 1649977179
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_287
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_288
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_289
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_290
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_291
timestamp 1649977179
transform -1 0 42780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_292
timestamp 1649977179
transform -1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_293
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_294
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_295
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_296
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_297
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_298
timestamp 1649977179
transform -1 0 45264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_299
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_300
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_301
timestamp 1649977179
transform -1 0 45908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_302
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_303
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_304
timestamp 1649977179
transform -1 0 46552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_305
timestamp 1649977179
transform -1 0 47196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_306
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_307
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_308
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_309
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_310
timestamp 1649977179
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_311
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_312
timestamp 1649977179
transform -1 0 48668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_313
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_314
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_315
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_316
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_317
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_318
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_319
timestamp 1649977179
transform -1 0 50508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_320
timestamp 1649977179
transform -1 0 51152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_321
timestamp 1649977179
transform 1 0 57960 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_322
timestamp 1649977179
transform 1 0 57960 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_323
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_324
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_325
timestamp 1649977179
transform -1 0 10672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_326
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_327
timestamp 1649977179
transform -1 0 11316 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_328
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_329
timestamp 1649977179
transform -1 0 11960 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_330
timestamp 1649977179
transform -1 0 12236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_331
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_332
timestamp 1649977179
transform -1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_333
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_334
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_335
timestamp 1649977179
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_336
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_337
timestamp 1649977179
transform 1 0 13248 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_338
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_339
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_340
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_341
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_342
timestamp 1649977179
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
<< labels >>
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 CMP_out_c
port 0 nsew signal tristate
flabel metal2 s 50250 59200 50306 60000 0 FreeSans 224 90 0 0 OTA_out_c
port 1 nsew signal tristate
flabel metal2 s 54942 59200 54998 60000 0 FreeSans 224 90 0 0 OTA_sh_c
port 2 nsew signal tristate
flabel metal2 s 40866 59200 40922 60000 0 FreeSans 224 90 0 0 Pd10_a
port 3 nsew signal tristate
flabel metal2 s 42430 59200 42486 60000 0 FreeSans 224 90 0 0 Pd10_b
port 4 nsew signal tristate
flabel metal2 s 43994 59200 44050 60000 0 FreeSans 224 90 0 0 Pd11_a
port 5 nsew signal tristate
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 Pd11_b
port 6 nsew signal tristate
flabel metal2 s 47122 59200 47178 60000 0 FreeSans 224 90 0 0 Pd12_a
port 7 nsew signal tristate
flabel metal2 s 48686 59200 48742 60000 0 FreeSans 224 90 0 0 Pd12_b
port 8 nsew signal tristate
flabel metal2 s 12714 59200 12770 60000 0 FreeSans 224 90 0 0 Pd1_a
port 9 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 Pd1_b
port 10 nsew signal tristate
flabel metal2 s 15842 59200 15898 60000 0 FreeSans 224 90 0 0 Pd2_a
port 11 nsew signal tristate
flabel metal2 s 17406 59200 17462 60000 0 FreeSans 224 90 0 0 Pd2_b
port 12 nsew signal tristate
flabel metal2 s 18970 59200 19026 60000 0 FreeSans 224 90 0 0 Pd3_a
port 13 nsew signal tristate
flabel metal2 s 20534 59200 20590 60000 0 FreeSans 224 90 0 0 Pd3_b
port 14 nsew signal tristate
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 Pd4_a
port 15 nsew signal tristate
flabel metal2 s 23662 59200 23718 60000 0 FreeSans 224 90 0 0 Pd4_b
port 16 nsew signal tristate
flabel metal2 s 25226 59200 25282 60000 0 FreeSans 224 90 0 0 Pd5_a
port 17 nsew signal tristate
flabel metal2 s 26790 59200 26846 60000 0 FreeSans 224 90 0 0 Pd5_b
port 18 nsew signal tristate
flabel metal2 s 28354 59200 28410 60000 0 FreeSans 224 90 0 0 Pd6_a
port 19 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 Pd6_b
port 20 nsew signal tristate
flabel metal2 s 31482 59200 31538 60000 0 FreeSans 224 90 0 0 Pd7_a
port 21 nsew signal tristate
flabel metal2 s 33046 59200 33102 60000 0 FreeSans 224 90 0 0 Pd7_b
port 22 nsew signal tristate
flabel metal2 s 34610 59200 34666 60000 0 FreeSans 224 90 0 0 Pd8_a
port 23 nsew signal tristate
flabel metal2 s 36174 59200 36230 60000 0 FreeSans 224 90 0 0 Pd8_b
port 24 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 Pd9_a
port 25 nsew signal tristate
flabel metal2 s 39302 59200 39358 60000 0 FreeSans 224 90 0 0 Pd9_b
port 26 nsew signal tristate
flabel metal2 s 51814 59200 51870 60000 0 FreeSans 224 90 0 0 SH_out_c
port 27 nsew signal tristate
flabel metal2 s 8022 59200 8078 60000 0 FreeSans 224 90 0 0 Sh
port 28 nsew signal tristate
flabel metal2 s 9586 59200 9642 60000 0 FreeSans 224 90 0 0 Sh_cmp
port 29 nsew signal tristate
flabel metal2 s 11150 59200 11206 60000 0 FreeSans 224 90 0 0 Sh_rst
port 30 nsew signal tristate
flabel metal2 s 4894 59200 4950 60000 0 FreeSans 224 90 0 0 Sw1
port 31 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 Sw2
port 32 nsew signal tristate
flabel metal2 s 1766 59200 1822 60000 0 FreeSans 224 90 0 0 Vd1
port 33 nsew signal tristate
flabel metal2 s 3330 59200 3386 60000 0 FreeSans 224 90 0 0 Vd2
port 34 nsew signal tristate
flabel metal2 s 56506 59200 56562 60000 0 FreeSans 224 90 0 0 Vref_cmp_c
port 35 nsew signal tristate
flabel metal2 s 58070 59200 58126 60000 0 FreeSans 224 90 0 0 Vref_sel_c
port 36 nsew signal tristate
flabel metal3 s 59200 52368 60000 52488 0 FreeSans 480 0 0 0 clk_o
port 37 nsew signal tristate
flabel metal3 s 59200 59168 60000 59288 0 FreeSans 480 0 0 0 counter_rst
port 38 nsew signal tristate
flabel metal3 s 59200 57808 60000 57928 0 FreeSans 480 0 0 0 data_o
port 39 nsew signal tristate
flabel metal3 s 59200 55088 60000 55208 0 FreeSans 480 0 0 0 done_o
port 40 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 io_in[0]
port 41 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_in[10]
port 42 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[11]
port 43 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 io_in[12]
port 44 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 io_in[13]
port 45 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 io_in[14]
port 46 nsew signal input
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 io_in[15]
port 47 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_in[16]
port 48 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 io_in[17]
port 49 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 io_in[18]
port 50 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_in[19]
port 51 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_in[1]
port 52 nsew signal input
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 io_in[20]
port 53 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 io_in[21]
port 54 nsew signal input
flabel metal3 s 0 35096 800 35216 0 FreeSans 480 0 0 0 io_in[22]
port 55 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 io_in[23]
port 56 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_in[24]
port 57 nsew signal input
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 io_in[25]
port 58 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 io_in[26]
port 59 nsew signal input
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 io_in[27]
port 60 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 io_in[28]
port 61 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_in[29]
port 62 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_in[2]
port 63 nsew signal input
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 io_in[30]
port 64 nsew signal input
flabel metal3 s 0 48560 800 48680 0 FreeSans 480 0 0 0 io_in[31]
port 65 nsew signal input
flabel metal3 s 0 50056 800 50176 0 FreeSans 480 0 0 0 io_in[32]
port 66 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 io_in[33]
port 67 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 io_in[34]
port 68 nsew signal input
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 io_in[35]
port 69 nsew signal input
flabel metal3 s 0 56040 800 56160 0 FreeSans 480 0 0 0 io_in[36]
port 70 nsew signal input
flabel metal3 s 0 57536 800 57656 0 FreeSans 480 0 0 0 io_in[37]
port 71 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 io_in[3]
port 72 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_in[4]
port 73 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[5]
port 74 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_in[6]
port 75 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_in[7]
port 76 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_in[8]
port 77 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_in[9]
port 78 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 79 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 80 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 81 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 82 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 83 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 84 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 85 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 86 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 87 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 88 nsew signal tristate
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 89 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 90 nsew signal tristate
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 91 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 92 nsew signal tristate
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 93 nsew signal tristate
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 94 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 95 nsew signal tristate
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 96 nsew signal tristate
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 97 nsew signal tristate
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 98 nsew signal tristate
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 99 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 100 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 101 nsew signal tristate
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 102 nsew signal tristate
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 103 nsew signal tristate
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 104 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 105 nsew signal tristate
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 106 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 107 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 108 nsew signal tristate
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 109 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 110 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 111 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 112 nsew signal tristate
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 113 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 114 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 115 nsew signal tristate
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 116 nsew signal tristate
flabel metal3 s 59200 688 60000 808 0 FreeSans 480 0 0 0 io_out[0]
port 117 nsew signal tristate
flabel metal3 s 59200 14288 60000 14408 0 FreeSans 480 0 0 0 io_out[10]
port 118 nsew signal tristate
flabel metal3 s 59200 15648 60000 15768 0 FreeSans 480 0 0 0 io_out[11]
port 119 nsew signal tristate
flabel metal3 s 59200 17008 60000 17128 0 FreeSans 480 0 0 0 io_out[12]
port 120 nsew signal tristate
flabel metal3 s 59200 18368 60000 18488 0 FreeSans 480 0 0 0 io_out[13]
port 121 nsew signal tristate
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 io_out[14]
port 122 nsew signal tristate
flabel metal3 s 59200 21088 60000 21208 0 FreeSans 480 0 0 0 io_out[15]
port 123 nsew signal tristate
flabel metal3 s 59200 22448 60000 22568 0 FreeSans 480 0 0 0 io_out[16]
port 124 nsew signal tristate
flabel metal3 s 59200 23808 60000 23928 0 FreeSans 480 0 0 0 io_out[17]
port 125 nsew signal tristate
flabel metal3 s 59200 25168 60000 25288 0 FreeSans 480 0 0 0 io_out[18]
port 126 nsew signal tristate
flabel metal3 s 59200 26528 60000 26648 0 FreeSans 480 0 0 0 io_out[19]
port 127 nsew signal tristate
flabel metal3 s 59200 2048 60000 2168 0 FreeSans 480 0 0 0 io_out[1]
port 128 nsew signal tristate
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 io_out[20]
port 129 nsew signal tristate
flabel metal3 s 59200 29248 60000 29368 0 FreeSans 480 0 0 0 io_out[21]
port 130 nsew signal tristate
flabel metal3 s 59200 30608 60000 30728 0 FreeSans 480 0 0 0 io_out[22]
port 131 nsew signal tristate
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 io_out[23]
port 132 nsew signal tristate
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 io_out[24]
port 133 nsew signal tristate
flabel metal3 s 59200 34688 60000 34808 0 FreeSans 480 0 0 0 io_out[25]
port 134 nsew signal tristate
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 io_out[26]
port 135 nsew signal tristate
flabel metal3 s 59200 37408 60000 37528 0 FreeSans 480 0 0 0 io_out[27]
port 136 nsew signal tristate
flabel metal3 s 59200 38768 60000 38888 0 FreeSans 480 0 0 0 io_out[28]
port 137 nsew signal tristate
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 io_out[29]
port 138 nsew signal tristate
flabel metal3 s 59200 3408 60000 3528 0 FreeSans 480 0 0 0 io_out[2]
port 139 nsew signal tristate
flabel metal3 s 59200 41488 60000 41608 0 FreeSans 480 0 0 0 io_out[30]
port 140 nsew signal tristate
flabel metal3 s 59200 42848 60000 42968 0 FreeSans 480 0 0 0 io_out[31]
port 141 nsew signal tristate
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 io_out[32]
port 142 nsew signal tristate
flabel metal3 s 59200 45568 60000 45688 0 FreeSans 480 0 0 0 io_out[33]
port 143 nsew signal tristate
flabel metal3 s 59200 46928 60000 47048 0 FreeSans 480 0 0 0 io_out[34]
port 144 nsew signal tristate
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 io_out[35]
port 145 nsew signal tristate
flabel metal3 s 59200 49648 60000 49768 0 FreeSans 480 0 0 0 io_out[36]
port 146 nsew signal tristate
flabel metal3 s 59200 51008 60000 51128 0 FreeSans 480 0 0 0 io_out[37]
port 147 nsew signal tristate
flabel metal3 s 59200 4768 60000 4888 0 FreeSans 480 0 0 0 io_out[3]
port 148 nsew signal tristate
flabel metal3 s 59200 6128 60000 6248 0 FreeSans 480 0 0 0 io_out[4]
port 149 nsew signal tristate
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 150 nsew signal tristate
flabel metal3 s 59200 8848 60000 8968 0 FreeSans 480 0 0 0 io_out[6]
port 151 nsew signal tristate
flabel metal3 s 59200 10208 60000 10328 0 FreeSans 480 0 0 0 io_out[7]
port 152 nsew signal tristate
flabel metal3 s 59200 11568 60000 11688 0 FreeSans 480 0 0 0 io_out[8]
port 153 nsew signal tristate
flabel metal3 s 59200 12928 60000 13048 0 FreeSans 480 0 0 0 io_out[9]
port 154 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 irq[0]
port 155 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 irq[1]
port 156 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 irq[2]
port 157 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 158 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 159 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 160 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 161 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 162 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 163 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 164 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 165 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 166 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 167 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 168 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 169 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 170 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 171 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 172 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 173 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 174 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 175 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 176 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 177 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 178 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 179 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 180 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 181 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 182 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 183 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 184 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 185 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 186 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 187 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 188 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 189 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 190 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 191 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 192 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 193 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 194 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 195 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 196 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 197 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 198 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 199 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 200 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 201 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 202 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 203 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 204 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 205 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 206 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 207 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 208 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 209 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 210 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 211 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 212 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 213 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 214 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 215 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 216 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 217 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 218 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 219 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 220 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 221 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 222 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 223 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 224 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 225 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 226 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 227 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 228 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 229 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 230 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 231 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 232 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 233 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 234 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 235 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 236 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 237 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 238 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 239 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 240 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 241 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 242 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 243 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 244 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 245 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 246 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 247 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 248 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 249 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 250 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 251 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 252 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 253 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 254 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 255 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 256 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 257 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 258 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 259 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 260 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 261 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 262 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 263 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 264 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 265 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 266 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 267 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 268 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 269 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 270 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 271 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 272 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 273 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 274 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 275 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 276 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 277 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 278 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 279 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 280 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 281 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 282 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 283 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 284 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 285 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 286 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 287 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 288 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 289 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 290 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 291 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 292 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 293 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 294 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 295 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 296 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 297 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 298 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 299 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 300 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 301 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 302 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 303 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 304 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 305 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 306 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 307 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 308 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 309 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 310 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 311 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 312 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 313 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 314 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 315 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 316 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 317 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 318 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 319 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 320 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 321 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 322 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 323 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 324 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 325 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 326 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 327 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 328 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 329 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 330 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 331 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 332 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 333 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 334 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 335 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 336 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 337 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 338 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 339 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 340 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 341 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 342 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 343 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 344 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 345 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 346 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 347 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 348 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 349 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 350 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 351 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 352 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 353 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 354 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 355 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 356 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 357 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 358 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 359 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 360 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 361 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 362 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 363 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 364 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 365 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 366 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 367 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 368 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 369 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 370 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 371 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 372 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 373 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 374 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 375 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 376 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 377 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 378 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 379 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 380 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 381 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 382 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 383 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 384 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 385 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 386 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 387 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 388 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 389 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 390 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 391 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 392 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 393 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 394 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 395 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 396 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 397 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 398 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 399 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 400 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 401 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 402 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 403 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 404 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 405 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 406 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 407 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 408 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 409 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 410 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 411 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 412 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 413 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 414 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 415 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 416 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 417 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 418 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 419 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 420 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 421 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 422 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 423 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 424 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 425 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 426 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 427 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 428 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 429 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 430 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 431 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 432 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 433 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 434 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 435 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 436 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 437 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 438 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 439 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 440 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 441 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 442 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 443 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 444 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 445 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 446 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 447 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 448 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 449 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 450 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 451 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 452 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 453 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 454 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 455 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 456 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 457 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 458 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 459 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 460 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 461 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 462 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 463 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 464 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 465 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 466 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 467 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 468 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 469 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 470 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 471 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 472 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 473 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 474 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 475 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 476 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 477 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 478 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 479 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 480 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 481 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 482 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 483 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 484 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 485 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 486 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 487 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 488 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 489 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 490 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 491 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 492 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 493 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 494 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 495 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 496 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 497 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 498 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 499 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 500 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 501 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 502 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 503 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 504 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 505 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 506 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 507 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 508 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 509 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 510 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 511 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 512 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 513 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 514 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 515 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 516 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 517 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 518 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 519 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 520 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 521 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 522 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 523 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 524 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 525 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 526 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 527 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 528 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 529 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 530 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 531 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 532 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 533 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 534 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 535 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 536 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 537 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 538 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 539 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 540 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 541 nsew signal input
flabel metal3 s 59200 53728 60000 53848 0 FreeSans 480 0 0 0 rst_o
port 542 nsew signal tristate
flabel metal3 s 59200 56448 60000 56568 0 FreeSans 480 0 0 0 start_o
port 543 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 544 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 544 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 545 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 545 nsew ground bidirectional
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wb_clk_i
port 546 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wb_rst_i
port 547 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 548 nsew signal tristate
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 549 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 550 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 551 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 552 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 553 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 554 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 555 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 556 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 557 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 558 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 559 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 560 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 561 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 562 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 563 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 564 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 565 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 566 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 567 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 568 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 569 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 570 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 571 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 572 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 573 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 574 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 575 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 576 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 577 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 578 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 579 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 580 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 581 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 582 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 583 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 584 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 585 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 586 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 587 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 588 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 589 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 590 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 591 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 592 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 593 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 594 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 595 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 596 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 597 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 598 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 599 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 600 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 601 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 602 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 603 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 604 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 605 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 606 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 607 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 608 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 609 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 610 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 611 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 612 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 613 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 614 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 615 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 616 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 617 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 618 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 619 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 620 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 621 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 622 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 623 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 624 nsew signal tristate
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 625 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 626 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 627 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 628 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 629 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 630 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 631 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 632 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 633 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 634 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 635 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 636 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 637 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 638 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 639 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 640 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 641 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 642 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 643 nsew signal tristate
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 644 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 645 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 646 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 647 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 648 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 649 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 650 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_we_i
port 651 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
