VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN gpio_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2530.870 3517.600 2531.430 3524.800 ;
    END
  END gpio_analog[0]
  PIN gpio_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.290 -4.800 795.850 2.400 ;
    END
  END gpio_analog[10]
  PIN gpio_analog[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2087.340 2924.800 2088.540 ;
    END
  END gpio_analog[11]
  PIN gpio_analog[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2865.940 2.400 2867.140 ;
    END
  END gpio_analog[12]
  PIN gpio_analog[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2967.940 2924.800 2969.140 ;
    END
  END gpio_analog[13]
  PIN gpio_analog[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 -4.800 283.870 2.400 ;
    END
  END gpio_analog[14]
  PIN gpio_analog[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.730 3517.600 802.290 3524.800 ;
    END
  END gpio_analog[15]
  PIN gpio_analog[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1063.940 2924.800 1065.140 ;
    END
  END gpio_analog[16]
  PIN gpio_analog[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2505.540 2.400 2506.740 ;
    END
  END gpio_analog[17]
  PIN gpio_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.290 -4.800 1117.850 2.400 ;
    END
  END gpio_analog[1]
  PIN gpio_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1145.540 2924.800 1146.740 ;
    END
  END gpio_analog[2]
  PIN gpio_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1342.740 2.400 1343.940 ;
    END
  END gpio_analog[3]
  PIN gpio_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.470 -4.800 2145.030 2.400 ;
    END
  END gpio_analog[4]
  PIN gpio_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 621.940 2924.800 623.140 ;
    END
  END gpio_analog[5]
  PIN gpio_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2566.740 2924.800 2567.940 ;
    END
  END gpio_analog[6]
  PIN gpio_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.350 3517.600 1352.910 3524.800 ;
    END
  END gpio_analog[7]
  PIN gpio_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1645.340 2924.800 1646.540 ;
    END
  END gpio_analog[8]
  PIN gpio_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2028.550 -4.800 2029.110 2.400 ;
    END
  END gpio_analog[9]
  PIN gpio_noesd[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END gpio_noesd[0]
  PIN gpio_noesd[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 683.140 2924.800 684.340 ;
    END
  END gpio_noesd[10]
  PIN gpio_noesd[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END gpio_noesd[11]
  PIN gpio_noesd[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2202.430 -4.800 2202.990 2.400 ;
    END
  END gpio_noesd[12]
  PIN gpio_noesd[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1380.140 2.400 1381.340 ;
    END
  END gpio_noesd[13]
  PIN gpio_noesd[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2046.540 2924.800 2047.740 ;
    END
  END gpio_noesd[14]
  PIN gpio_noesd[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 604.940 2924.800 606.140 ;
    END
  END gpio_noesd[15]
  PIN gpio_noesd[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3328.340 2924.800 3329.540 ;
    END
  END gpio_noesd[16]
  PIN gpio_noesd[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.570 -4.800 1839.130 2.400 ;
    END
  END gpio_noesd[17]
  PIN gpio_noesd[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.830 -4.800 1462.390 2.400 ;
    END
  END gpio_noesd[1]
  PIN gpio_noesd[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1624.940 2924.800 1626.140 ;
    END
  END gpio_noesd[2]
  PIN gpio_noesd[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2107.740 2924.800 2108.940 ;
    END
  END gpio_noesd[3]
  PIN gpio_noesd[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2846.430 -4.800 2846.990 2.400 ;
    END
  END gpio_noesd[4]
  PIN gpio_noesd[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.730 3517.600 1124.290 3524.800 ;
    END
  END gpio_noesd[5]
  PIN gpio_noesd[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3345.340 2.400 3346.540 ;
    END
  END gpio_noesd[6]
  PIN gpio_noesd[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 3517.600 1864.890 3524.800 ;
    END
  END gpio_noesd[7]
  PIN gpio_noesd[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.190 -4.800 2067.750 2.400 ;
    END
  END gpio_noesd[8]
  PIN gpio_noesd[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3168.540 2924.800 3169.740 ;
    END
  END gpio_noesd[9]
  PIN io_analog[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 740.940 2.400 742.140 ;
    END
  END io_analog[0]
  PIN io_analog[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.570 -4.800 1195.130 2.400 ;
    END
  END io_analog[10]
  PIN io_analog[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.390 3517.600 650.950 3524.800 ;
    END
  END io_analog[1]
  PIN io_analog[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 159.540 2.400 160.740 ;
    END
  END io_analog[2]
  PIN io_analog[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1019.740 2.400 1020.940 ;
    END
  END io_analog[3]
  PIN io_analog[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 -4.800 303.190 2.400 ;
    END
  END io_analog[4]
  PIN io_analog[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.370 3517.600 1484.930 3524.800 ;
    END
  END io_analog[5]
  PIN io_analog[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3467.740 2.400 3468.940 ;
    END
  END io_analog[6]
  PIN io_analog[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2808.140 2924.800 2809.340 ;
    END
  END io_analog[7]
  PIN io_analog[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3365.740 2.400 3366.940 ;
    END
  END io_analog[8]
  PIN io_analog[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.610 3517.600 1942.170 3524.800 ;
    END
  END io_analog[9]
  PIN io_clamp_high[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.750 3517.600 934.310 3524.800 ;
    END
  END io_clamp_high[0]
  PIN io_clamp_high[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2124.740 2.400 2125.940 ;
    END
  END io_clamp_high[1]
  PIN io_clamp_high[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 -4.800 113.210 2.400 ;
    END
  END io_clamp_high[2]
  PIN io_clamp_low[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3090.340 2924.800 3091.540 ;
    END
  END io_clamp_low[0]
  PIN io_clamp_low[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 802.140 2924.800 803.340 ;
    END
  END io_clamp_low[1]
  PIN io_clamp_low[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 278.540 2.400 279.740 ;
    END
  END io_clamp_low[2]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2689.140 2924.800 2690.340 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1784.740 2924.800 1785.940 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 462.140 2924.800 463.340 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.670 -4.800 567.230 2.400 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 3517.600 174.390 3524.800 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2205.650 3517.600 2206.210 3524.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1084.340 2924.800 1085.540 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.470 -4.800 2467.030 2.400 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1907.140 2924.800 1908.340 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.330 -4.800 737.890 2.400 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2665.340 2.400 2666.540 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.730 3517.600 480.290 3524.800 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.590 3517.600 1810.150 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.490 3517.600 345.050 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.510 -4.800 2087.070 2.400 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.590 -4.800 683.150 2.400 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1199.940 2.400 1201.140 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.710 3517.600 670.270 3524.800 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2427.340 2924.800 2428.540 ;
    END
  END io_in[26]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.610 -4.800 493.170 2.400 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.330 -4.800 415.890 2.400 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2828.540 2924.800 2829.740 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.510 -4.800 1443.070 2.400 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3086.940 2.400 3088.140 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1703.140 2.400 1704.340 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 343.140 2924.800 344.340 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 961.940 2.400 963.140 ;
    END
  END io_in[9]
  PIN io_in_3v3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.670 3517.600 1694.230 3524.800 ;
    END
  END io_in_3v3[0]
  PIN io_in_3v3[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1961.540 2.400 1962.740 ;
    END
  END io_in_3v3[10]
  PIN io_in_3v3[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.650 -4.800 435.210 2.400 ;
    END
  END io_in_3v3[11]
  PIN io_in_3v3[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.390 3517.600 1294.950 3524.800 ;
    END
  END io_in_3v3[12]
  PIN io_in_3v3[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.750 3517.600 612.310 3524.800 ;
    END
  END io_in_3v3[13]
  PIN io_in_3v3[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1560.340 2.400 1561.540 ;
    END
  END io_in_3v3[14]
  PIN io_in_3v3[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 744.340 2924.800 745.540 ;
    END
  END io_in_3v3[15]
  PIN io_in_3v3[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 880.340 2.400 881.540 ;
    END
  END io_in_3v3[16]
  PIN io_in_3v3[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.690 -4.800 55.250 2.400 ;
    END
  END io_in_3v3[17]
  PIN io_in_3v3[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3246.740 2.400 3247.940 ;
    END
  END io_in_3v3[18]
  PIN io_in_3v3[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.630 3517.600 2074.190 3524.800 ;
    END
  END io_in_3v3[19]
  PIN io_in_3v3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2889.740 2924.800 2890.940 ;
    END
  END io_in_3v3[1]
  PIN io_in_3v3[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2104.340 2.400 2105.540 ;
    END
  END io_in_3v3[20]
  PIN io_in_3v3[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.090 3517.600 1085.650 3524.800 ;
    END
  END io_in_3v3[21]
  PIN io_in_3v3[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.170 -4.800 2257.730 2.400 ;
    END
  END io_in_3v3[22]
  PIN io_in_3v3[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 322.740 2924.800 323.940 ;
    END
  END io_in_3v3[23]
  PIN io_in_3v3[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3144.740 2.400 3145.940 ;
    END
  END io_in_3v3[24]
  PIN io_in_3v3[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1985.340 2924.800 1986.540 ;
    END
  END io_in_3v3[25]
  PIN io_in_3v3[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1068.990 3517.600 1069.550 3524.800 ;
    END
  END io_in_3v3[26]
  PIN io_in_3v3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3250.140 2924.800 3251.340 ;
    END
  END io_in_3v3[2]
  PIN io_in_3v3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2825.140 2.400 2826.340 ;
    END
  END io_in_3v3[3]
  PIN io_in_3v3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.070 3517.600 631.630 3524.800 ;
    END
  END io_in_3v3[4]
  PIN io_in_3v3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.230 -4.800 1365.790 2.400 ;
    END
  END io_in_3v3[5]
  PIN io_in_3v3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2910.140 2924.800 2911.340 ;
    END
  END io_in_3v3[6]
  PIN io_in_3v3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.310 3517.600 1732.870 3524.800 ;
    END
  END io_in_3v3[7]
  PIN io_in_3v3[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 319.340 2.400 320.540 ;
    END
  END io_in_3v3[8]
  PIN io_in_3v3[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2617.810 -4.800 2618.370 2.400 ;
    END
  END io_in_3v3[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3029.140 2924.800 3030.340 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1485.540 2924.800 1486.740 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.730 3517.600 1446.290 3524.800 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.550 -4.800 1063.110 2.400 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1023.140 2924.800 1024.340 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1981.940 2.400 1983.140 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 863.340 2924.800 864.540 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 842.940 2924.800 844.140 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 598.140 2.400 599.340 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1822.140 2.400 1823.340 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 421.340 2924.800 422.540 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.250 3517.600 1980.810 3524.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1359.740 2.400 1360.940 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 438.340 2.400 439.540 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1264.540 2924.800 1265.740 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.930 -4.800 834.490 2.400 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2944.140 2.400 2945.340 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2002.340 2.400 2003.540 ;
    END
  END io_oeb[26]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1601.140 2.400 1602.340 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.770 3517.600 744.330 3524.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.710 3517.600 1636.270 3524.800 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 383.940 2924.800 385.140 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 581.140 2.400 582.340 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.450 3517.600 725.010 3524.800 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2736.950 3517.600 2737.510 3524.800 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.950 -4.800 644.510 2.400 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 118.740 2.400 119.940 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2083.940 2.400 2085.140 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.070 -4.800 2563.630 2.400 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3491.540 2924.800 3492.740 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.950 3517.600 2415.510 3524.800 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.430 3517.600 914.990 3524.800 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3369.140 2924.800 3370.340 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1482.140 2.400 1483.340 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.150 3517.600 193.710 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2852.870 3517.600 2853.430 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.890 3517.600 2341.450 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3290.940 2924.800 3292.140 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.630 3517.600 1430.190 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3185.540 2.400 3186.740 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 3517.600 2225.530 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3229.740 2924.800 3230.940 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 16.740 2.400 17.940 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 302.340 2924.800 303.540 ;
    END
  END io_out[26]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2522.540 2.400 2523.740 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1686.140 2924.800 1687.340 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3505.140 2.400 3506.340 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3447.340 2.400 3448.540 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2264.140 2.400 2265.340 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.570 -4.800 873.130 2.400 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 -4.800 225.910 2.400 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2598.490 -4.800 2599.050 2.400 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.090 3517.600 119.650 3524.800 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2988.340 2924.800 2989.540 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2804.740 2.400 2805.940 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1903.740 2.400 1904.940 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.650 3517.600 1884.210 3524.800 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.910 -4.800 1346.470 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1125.140 2924.800 1126.340 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 40.540 2924.800 41.740 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3124.340 2.400 3125.540 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2604.140 2.400 2605.340 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.830 -4.800 2428.390 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 237.740 2.400 238.940 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2648.340 2924.800 2649.540 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 122.140 2924.800 123.340 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3406.540 2.400 3407.740 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 921.140 2.400 922.340 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.530 -4.800 1575.090 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1947.940 2924.800 1949.140 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 900.740 2.400 901.940 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2563.340 2.400 2564.540 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.850 -4.800 2238.410 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2675.770 -4.800 2676.330 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1505.940 2924.800 1507.140 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.990 3517.600 1713.550 3524.800 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2423.940 2.400 2425.140 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2468.140 2924.800 2469.340 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 3517.600 1220.890 3524.800 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.610 -4.800 815.170 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3107.340 2.400 3108.540 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1346.140 2924.800 1347.340 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2223.340 2.400 2224.540 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.150 -4.800 2447.710 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2947.540 2924.800 2948.740 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3131.140 2924.800 3132.340 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2128.140 2924.800 2129.340 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.270 -4.800 1307.830 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2767.340 2924.800 2768.540 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2723.140 2.400 2724.340 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.190 -4.800 2389.750 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 819.140 2.400 820.340 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 543.740 2924.800 544.940 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1723.540 2.400 1724.740 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.570 -4.800 1517.130 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 3517.600 2586.170 3524.800 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 944.940 2924.800 946.140 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.130 -4.800 2315.690 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3488.140 2.400 3489.340 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.570 3517.600 2644.130 3524.800 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3025.740 2.400 3026.940 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1522.940 2.400 1524.140 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.930 -4.800 1478.490 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2284.540 2.400 2285.740 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.690 -4.800 377.250 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.010 3517.600 879.570 3524.800 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.010 3517.600 1523.570 3524.800 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1662.340 2.400 1663.540 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3287.540 2.400 3288.740 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2607.540 2924.800 2608.740 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2267.540 2924.800 2268.740 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 798.740 2.400 799.940 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.730 -4.800 2734.290 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2701.530 3517.600 2702.090 3524.800 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 261.540 2924.800 262.740 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1825.540 2924.800 1826.740 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 380.540 2.400 381.740 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 37.140 2.400 38.340 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1023.910 -4.800 1024.470 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 720.540 2.400 721.740 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 203.740 2924.800 204.940 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.650 -4.800 757.210 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.270 -4.800 985.830 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1567.140 2924.800 1568.340 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.390 -4.800 2904.950 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.030 3517.600 1333.590 3524.800 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2141.740 2.400 2142.940 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 618.540 2.400 619.740 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.710 3517.600 1314.270 3524.800 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2549.740 2924.800 2550.940 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2743.540 2.400 2744.740 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.950 -4.800 1288.510 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 -4.800 16.610 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2206.340 2924.800 2207.540 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 162.940 2924.800 164.140 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.750 3517.600 290.310 3524.800 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2508.940 2924.800 2510.140 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 479.140 2.400 480.340 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2444.340 2.400 2445.540 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2644.940 2.400 2646.140 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3386.140 2.400 3387.340 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 281.940 2924.800 283.140 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2244.290 3517.600 2244.850 3524.800 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 904.140 2924.800 905.340 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2930.540 2924.800 2931.740 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1706.540 2924.800 1707.740 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.010 -4.800 396.570 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2869.340 2924.800 2870.540 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1543.340 2.400 1544.540 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.430 3517.600 592.990 3524.800 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2746.940 2924.800 2748.140 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1960.930 3517.600 1961.490 3524.800 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2604.930 3517.600 2605.490 3524.800 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1441.340 2.400 1442.540 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1665.740 2924.800 1666.940 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3389.540 2924.800 3390.740 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.390 3517.600 972.950 3524.800 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.910 3517.600 2473.470 3524.800 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.370 3517.600 1162.930 3524.800 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2403.540 2.400 2404.740 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 360.140 2.400 361.340 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2453.590 3517.600 2454.150 3524.800 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1641.940 2.400 1643.140 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1747.340 2924.800 1748.540 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 458.740 2.400 459.940 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3.140 2924.800 4.340 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1420.940 2.400 1422.140 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 519.940 2.400 521.140 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.290 -4.800 473.850 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 978.940 2.400 980.140 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.850 -4.800 1272.410 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.550 -4.800 1385.110 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.110 3517.600 251.670 3524.800 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2769.150 -4.800 2769.710 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2775.590 3517.600 2776.150 3524.800 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1162.540 2.400 1163.740 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1604.540 2924.800 1605.740 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 946.630 -4.800 947.190 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2542.940 2.400 2544.140 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3046.140 2.400 3047.340 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.190 -4.800 1423.750 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 985.740 2924.800 986.940 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2066.940 2924.800 2068.140 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3426.940 2.400 3428.140 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3226.340 2.400 3227.540 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.930 -4.800 1156.490 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.050 3517.600 821.610 3524.800 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1305.340 2924.800 1306.540 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.410 3517.600 782.970 3524.800 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.770 3517.600 422.330 3524.800 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.970 -4.800 776.530 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1964.940 2924.800 1966.140 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2325.340 2.400 2326.540 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.550 3517.600 2512.110 3524.800 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1924.140 2.400 1925.340 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1060.540 2.400 1061.740 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2833.550 3517.600 2834.110 3524.800 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2485.140 2.400 2486.340 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.590 -4.800 1005.150 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2814.230 3517.600 2814.790 3524.800 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 339.740 2.400 340.940 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3270.540 2924.800 3271.740 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2005.740 2924.800 2006.940 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 142.540 2924.800 143.740 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 941.540 2.400 942.740 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.330 -4.800 93.890 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 3517.600 895.670 3524.800 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 3517.600 535.030 3524.800 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2376.310 3517.600 2376.870 3524.800 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 703.540 2924.800 704.740 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2447.740 2924.800 2448.940 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 139.140 2.400 140.340 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1424.340 2924.800 1425.540 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.610 -4.800 1137.170 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 220.740 2924.800 221.940 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1973.810 -4.800 1974.370 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.090 3517.600 441.650 3524.800 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.350 3517.600 1674.910 3524.800 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.370 3517.600 840.930 3524.800 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.570 -4.800 551.130 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2349.140 2924.800 2350.340 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2243.740 2.400 2244.940 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2524.430 -4.800 2524.990 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1165.940 2924.800 1167.140 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 3517.600 2911.390 3524.800 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2202.940 2.400 2204.140 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 81.340 2924.800 82.540 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2360.210 3517.600 2360.770 3524.800 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2386.540 2924.800 2387.740 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1886.740 2924.800 1887.940 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.210 -4.800 1555.770 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1535.890 -4.800 1536.450 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2063.540 2.400 2064.740 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2165.540 2924.800 2166.740 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1179.540 2.400 1180.740 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1584.140 2924.800 1585.340 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1043.540 2924.800 1044.740 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 638.940 2.400 640.140 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 785.140 2924.800 786.340 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2624.250 3517.600 2624.810 3524.800 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 60.940 2924.800 62.140 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 363.540 2924.800 364.740 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 662.740 2924.800 663.940 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.970 3517.600 1259.530 3524.800 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1767.740 2924.800 1768.940 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.170 -4.800 1613.730 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.010 3517.600 1201.570 3524.800 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3165.140 2.400 3166.340 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.770 -4.800 2354.330 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1896.530 -4.800 1897.090 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.450 3517.600 403.010 3524.800 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.070 3517.600 309.630 3524.800 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2583.740 2.400 2584.940 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.350 3517.600 708.910 3524.800 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1142.140 2.400 1143.340 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1760.940 2.400 1762.140 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 417.940 2.400 419.140 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.230 3517.600 2170.790 3524.800 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.130 -4.800 1993.690 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 999.340 2.400 1000.540 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.670 3517.600 1372.230 3524.800 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2247.140 2924.800 2248.340 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 642.340 2924.800 643.540 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2148.540 2924.800 2149.740 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.830 -4.800 1784.390 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3205.940 2.400 3207.140 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.610 3517.600 2264.170 3524.800 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2150.910 3517.600 2151.470 3524.800 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2342.340 2.400 2343.540 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2685.740 2.400 2686.940 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.070 3517.600 953.630 3524.800 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1223.740 2924.800 1224.940 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 924.540 2924.800 925.740 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.850 -4.800 1594.410 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.090 -4.800 2373.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.210 -4.800 1233.770 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2186.330 3517.600 2186.890 3524.800 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1803.150 -4.800 1803.710 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.170 3517.600 3.730 3524.800 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2304.940 2.400 2306.140 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3324.940 2.400 3326.140 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2406.940 2924.800 2408.140 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 764.740 2924.800 765.940 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 241.140 2924.800 242.340 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1186.340 2924.800 1187.540 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2845.540 2.400 2846.740 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.530 -4.800 1253.090 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 298.940 2.400 300.140 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.450 -4.800 2335.010 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.290 3517.600 2566.850 3524.800 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.790 3517.600 554.350 3524.800 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1400.540 2.400 1401.740 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 560.740 2.400 561.940 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 404.340 2924.800 405.540 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.470 3517.600 213.030 3524.800 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.410 3517.600 1104.970 3524.800 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.150 -4.800 2125.710 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1842.540 2.400 1843.740 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 2.400 1041.340 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.790 -4.800 2486.350 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2807.790 -4.800 2808.350 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.490 3517.600 23.050 3524.800 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.130 3517.600 383.690 3524.800 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2756.270 3517.600 2756.830 3524.800 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.170 -4.800 2579.730 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.130 3517.600 61.690 3524.800 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.270 3517.600 2112.830 3524.800 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.670 3517.600 2016.230 3524.800 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2383.140 2.400 2384.340 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.250 -4.800 1497.810 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.510 -4.800 1765.070 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.890 3517.600 2663.450 3524.800 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 822.540 2924.800 823.740 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.950 3517.600 2093.510 3524.800 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.250 -4.800 853.810 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2366.140 2924.800 2367.340 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 3517.600 860.250 3524.800 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 3517.600 2550.750 3524.800 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.730 3517.600 158.290 3524.800 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1902.970 3517.600 1903.530 3524.800 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1621.540 2.400 1622.740 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3008.740 2924.800 3009.940 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2185.940 2924.800 2187.140 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.630 -4.800 625.190 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 397.540 2.400 398.740 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2162.140 2.400 2163.340 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.550 -4.800 1707.110 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2794.910 3517.600 2795.470 3524.800 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1883.340 2.400 1884.540 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1682.740 2.400 1683.940 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.810 3517.600 42.370 3524.800 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 3517.600 232.350 3524.800 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.250 -4.800 1175.810 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.310 3517.600 1410.870 3524.800 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3209.340 2924.800 3210.540 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1526.340 2924.800 1527.540 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1580.740 2.400 1581.940 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1244.140 2924.800 1245.340 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2729.940 2924.800 2731.140 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.990 3517.600 1391.550 3524.800 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 761.340 2.400 762.540 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.310 -4.800 927.870 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 965.340 2924.800 966.540 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 -4.800 206.590 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 883.740 2924.800 884.940 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2891.510 3517.600 2892.070 3524.800 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1805.140 2924.800 1806.340 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1080.940 2.400 1082.140 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 77.940 2.400 79.140 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1220.340 2.400 1221.540 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2105.830 -4.800 2106.390 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2226.740 2924.800 2227.940 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.210 3517.600 2682.770 3524.800 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2984.940 2.400 2986.140 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 3517.600 1504.250 3524.800 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.850 3517.600 2721.410 3524.800 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.810 3517.600 364.370 3524.800 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1502.540 2.400 1503.740 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 584.540 2924.800 585.740 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1465.140 2924.800 1466.340 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2328.740 2924.800 2329.940 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1049.670 3517.600 1050.230 3524.800 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.110 -4.800 2505.670 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3267.140 2.400 3268.340 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 499.540 2.400 500.740 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.270 3517.600 2434.830 3524.800 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3409.940 2924.800 3411.140 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 101.740 2924.800 102.940 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 57.540 2.400 58.740 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2885.070 -4.800 2885.630 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 564.140 2924.800 565.340 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.990 -4.800 586.550 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.890 -4.800 892.450 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 183.340 2924.800 184.540 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1366.540 2924.800 1367.740 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3110.740 2924.800 3111.940 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.050 3517.600 1143.610 3524.800 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.030 3517.600 1011.590 3524.800 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 3517.600 499.610 3524.800 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1101.190 -4.800 1101.750 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3450.740 2924.800 3451.940 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 778.340 2.400 779.540 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.390 3517.600 328.950 3524.800 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 258.140 2.400 259.340 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3049.540 2924.800 3050.740 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.630 3517.600 1752.190 3524.800 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.650 3517.600 1562.210 3524.800 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.590 3517.600 2132.150 3524.800 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.250 3517.600 2302.810 3524.800 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.570 3517.600 2322.130 3524.800 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1261.140 2.400 1262.340 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.650 3517.600 1240.210 3524.800 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1121.740 2.400 1122.940 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.370 -4.800 35.930 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2865.750 -4.800 2866.310 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1002.740 2924.800 1003.940 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 3517.600 1581.530 3524.800 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1325.740 2924.800 1326.940 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2906.740 2.400 2907.940 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1301.940 2.400 1303.140 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 859.940 2.400 861.140 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.690 3517.600 1182.250 3524.800 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 23.540 2924.800 24.740 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.870 -4.800 1404.430 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2464.740 2.400 2465.940 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2668.740 2924.800 2669.940 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3348.740 2924.800 3349.940 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2827.110 -4.800 2827.670 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2923.740 2.400 2924.940 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 659.340 2.400 660.540 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3188.940 2924.800 3190.140 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.090 3517.600 763.650 3524.800 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 196.940 2.400 198.140 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2753.050 -4.800 2753.610 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.330 3517.600 1542.890 3524.800 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1104.740 2924.800 1105.940 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.370 3517.600 518.930 3524.800 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1862.940 2.400 1864.140 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2784.340 2.400 2785.540 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.970 -4.800 454.530 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2587.140 2924.800 2588.340 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_oenb[9]
  PIN pxl_done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1101.340 2.400 1102.540 ;
    END
  END pxl_done
  PIN pxl_start_in_path
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.210 -4.800 911.770 2.400 ;
    END
  END pxl_start_in_path
  PIN pxl_start_out_path
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1461.740 2.400 1462.940 ;
    END
  END pxl_start_out_path
  PIN serial_data_rlbp_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3066.540 2.400 3067.740 ;
    END
  END serial_data_rlbp_out
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.290 3517.600 1600.850 3524.800 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3511.940 2924.800 3513.140 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3304.540 2.400 3305.740 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -38.270 12.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -38.270 192.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -38.270 372.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -38.270 552.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -38.270 732.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 710.000 732.070 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1310.000 732.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -38.270 912.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 710.000 912.070 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 1310.000 912.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -38.270 1092.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -38.270 1272.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -38.270 1452.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -38.270 1632.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -38.270 1812.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -38.270 1992.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -38.270 2172.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -38.270 2352.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -38.270 2532.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -38.270 2712.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -38.270 2892.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 14.330 2963.250 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 194.330 2963.250 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 374.330 2963.250 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 554.330 2963.250 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 734.330 2963.250 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 914.330 2963.250 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1094.330 2963.250 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1274.330 2963.250 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1454.330 2963.250 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1634.330 2963.250 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1814.330 2963.250 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1994.330 2963.250 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2174.330 2963.250 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2354.330 2963.250 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2534.330 2963.250 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2714.330 2963.250 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2894.330 2963.250 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3074.330 2963.250 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3254.330 2963.250 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3434.330 2963.250 3437.430 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.970 -38.270 57.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.970 -38.270 237.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.970 -38.270 417.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 -38.270 597.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 710.000 597.070 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 1310.000 597.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 -38.270 777.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 710.000 777.070 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 1310.000 777.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.970 -38.270 957.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.970 710.000 957.070 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.970 1310.000 957.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1133.970 -38.270 1137.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1313.970 -38.270 1317.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.970 -38.270 1497.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1673.970 -38.270 1677.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1853.970 -38.270 1857.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2033.970 -38.270 2037.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2213.970 -38.270 2217.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.970 -38.270 2397.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2573.970 -38.270 2577.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2753.970 -38.270 2757.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 59.330 2963.250 62.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 239.330 2963.250 242.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 419.330 2963.250 422.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 599.330 2963.250 602.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 779.330 2963.250 782.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 959.330 2963.250 962.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1139.330 2963.250 1142.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1319.330 2963.250 1322.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1499.330 2963.250 1502.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1679.330 2963.250 1682.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1859.330 2963.250 1862.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2039.330 2963.250 2042.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2219.330 2963.250 2222.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2399.330 2963.250 2402.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2579.330 2963.250 2582.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2759.330 2963.250 2762.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2939.330 2963.250 2942.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3119.330 2963.250 3122.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3299.330 2963.250 3302.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3479.330 2963.250 3482.430 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 -38.270 102.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 -38.270 282.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -38.270 462.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -38.270 642.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1310.000 642.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 -38.270 822.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 1310.000 822.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 -38.270 1002.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 -38.270 1182.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -38.270 1362.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 -38.270 1542.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 -38.270 1722.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -38.270 1902.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 -38.270 2082.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -38.270 2262.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 -38.270 2442.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 -38.270 2622.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 -38.270 2802.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 104.330 2963.250 107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 284.330 2963.250 287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 464.330 2963.250 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 644.330 2963.250 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 824.330 2963.250 827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1004.330 2963.250 1007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1184.330 2963.250 1187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1364.330 2963.250 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1544.330 2963.250 1547.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1724.330 2963.250 1727.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1904.330 2963.250 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2084.330 2963.250 2087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2264.330 2963.250 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2444.330 2963.250 2447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2624.330 2963.250 2627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2804.330 2963.250 2807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2984.330 2963.250 2987.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3164.330 2963.250 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3344.330 2963.250 3347.430 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.970 -38.270 147.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 -38.270 327.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.970 -38.270 507.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 -38.270 687.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 1310.000 687.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 -38.270 867.070 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 1310.000 867.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1043.970 -38.270 1047.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.970 -38.270 1227.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.970 -38.270 1407.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1583.970 -38.270 1587.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.970 -38.270 1767.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.970 -38.270 1947.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 -38.270 2127.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2303.970 -38.270 2307.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2483.970 -38.270 2487.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2663.970 -38.270 2667.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2843.970 -38.270 2847.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 149.330 2963.250 152.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 329.330 2963.250 332.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 509.330 2963.250 512.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 689.330 2963.250 692.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 869.330 2963.250 872.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1049.330 2963.250 1052.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1229.330 2963.250 1232.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1409.330 2963.250 1412.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1589.330 2963.250 1592.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1769.330 2963.250 1772.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1949.330 2963.250 1952.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2129.330 2963.250 2132.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2309.330 2963.250 2312.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2489.330 2963.250 2492.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2669.330 2963.250 2672.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2849.330 2963.250 2852.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3029.330 2963.250 3032.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3209.330 2963.250 3212.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3389.330 2963.250 3392.430 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.470 -38.270 124.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.470 -38.270 304.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.470 -38.270 484.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 -38.270 664.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 1310.000 664.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 841.470 -38.270 844.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 841.470 1310.000 844.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.470 -38.270 1024.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1201.470 -38.270 1204.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1381.470 -38.270 1384.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1561.470 -38.270 1564.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1741.470 -38.270 1744.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.470 -38.270 1924.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2101.470 -38.270 2104.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 -38.270 2284.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2461.470 -38.270 2464.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2641.470 -38.270 2644.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2821.470 -38.270 2824.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 126.830 2963.250 129.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 306.830 2963.250 309.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 486.830 2963.250 489.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 666.830 2963.250 669.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 846.830 2963.250 849.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1026.830 2963.250 1029.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1206.830 2963.250 1209.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1386.830 2963.250 1389.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1566.830 2963.250 1569.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1746.830 2963.250 1749.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1926.830 2963.250 1929.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2106.830 2963.250 2109.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2286.830 2963.250 2289.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2466.830 2963.250 2469.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2646.830 2963.250 2649.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2826.830 2963.250 2829.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3006.830 2963.250 3009.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3186.830 2963.250 3189.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3366.830 2963.250 3369.930 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.470 -38.270 169.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 -38.270 349.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.470 -38.270 529.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 -38.270 709.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 710.000 709.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 1310.000 709.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 -38.270 889.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 710.000 889.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 1310.000 889.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1066.470 -38.270 1069.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.470 -38.270 1249.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1426.470 -38.270 1429.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1606.470 -38.270 1609.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.470 -38.270 1789.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.470 -38.270 1969.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.470 -38.270 2149.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2326.470 -38.270 2329.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2506.470 -38.270 2509.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2686.470 -38.270 2689.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2866.470 -38.270 2869.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 171.830 2963.250 174.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 351.830 2963.250 354.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 531.830 2963.250 534.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 711.830 2963.250 714.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 891.830 2963.250 894.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1071.830 2963.250 1074.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1251.830 2963.250 1254.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1431.830 2963.250 1434.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1611.830 2963.250 1614.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1791.830 2963.250 1794.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1971.830 2963.250 1974.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2151.830 2963.250 2154.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2331.830 2963.250 2334.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2511.830 2963.250 2514.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2691.830 2963.250 2694.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2871.830 2963.250 2874.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3051.830 2963.250 3054.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3231.830 2963.250 3234.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3411.830 2963.250 3414.930 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.470 -38.270 34.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 -38.270 214.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 -38.270 394.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 -38.270 574.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 -38.270 754.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 710.000 754.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 1310.000 754.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.470 -38.270 934.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.470 710.000 934.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.470 1310.000 934.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1111.470 -38.270 1114.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1291.470 -38.270 1294.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.470 -38.270 1474.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.470 -38.270 1654.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 -38.270 1834.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 -38.270 2014.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.470 -38.270 2194.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.470 -38.270 2374.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2551.470 -38.270 2554.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.470 -38.270 2734.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2911.470 -38.270 2914.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 36.830 2963.250 39.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 216.830 2963.250 219.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 396.830 2963.250 399.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 576.830 2963.250 579.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 756.830 2963.250 759.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 936.830 2963.250 939.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1116.830 2963.250 1119.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1296.830 2963.250 1299.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1476.830 2963.250 1479.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1656.830 2963.250 1659.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1836.830 2963.250 1839.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2016.830 2963.250 2019.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2196.830 2963.250 2199.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2376.830 2963.250 2379.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2556.830 2963.250 2559.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2736.830 2963.250 2739.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2916.830 2963.250 2919.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3096.830 2963.250 3099.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3276.830 2963.250 3279.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3456.830 2963.250 3459.930 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.470 -38.270 79.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.470 -38.270 259.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.470 -38.270 439.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 -38.270 619.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 710.000 619.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 1310.000 619.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 -38.270 799.570 390.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 710.000 799.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 1310.000 799.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 976.470 -38.270 979.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.470 -38.270 1159.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1336.470 -38.270 1339.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.470 -38.270 1519.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.470 -38.270 1699.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1876.470 -38.270 1879.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.470 -38.270 2059.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.470 -38.270 2239.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2416.470 -38.270 2419.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2596.470 -38.270 2599.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2776.470 -38.270 2779.570 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 81.830 2963.250 84.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 261.830 2963.250 264.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 441.830 2963.250 444.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 621.830 2963.250 624.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 801.830 2963.250 804.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 981.830 2963.250 984.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1161.830 2963.250 1164.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1341.830 2963.250 1344.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1521.830 2963.250 1524.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1701.830 2963.250 1704.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1881.830 2963.250 1884.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2061.830 2963.250 2064.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2241.830 2963.250 2244.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2421.830 2963.250 2424.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2601.830 2963.250 2604.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2781.830 2963.250 2784.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2961.830 2963.250 2964.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3141.830 2963.250 3144.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3321.830 2963.250 3324.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3501.830 2963.250 3504.930 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1284.940 2924.800 1286.140 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1743.940 2.400 1745.140 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1927.540 2924.800 1928.740 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.710 3517.600 992.270 3524.800 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.430 3517.600 270.990 3524.800 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2362.740 2.400 2363.940 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.950 -4.800 322.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1801.740 2.400 1802.940 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3311.340 2924.800 3312.540 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3069.940 2924.800 3071.140 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.530 -4.800 2219.090 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2787.740 2924.800 2788.940 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1726.940 2924.800 1728.140 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 441.740 2924.800 442.940 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.350 3517.600 1030.910 3524.800 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.990 3517.600 2035.550 3524.800 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1954.490 -4.800 1955.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2788.470 -4.800 2789.030 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1383.540 2924.800 1384.740 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2763.940 2.400 2765.140 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.210 -4.800 1877.770 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.590 -4.800 361.150 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 98.340 2.400 99.540 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2627.940 2924.800 2629.140 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2492.230 3517.600 2492.790 3524.800 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.030 3517.600 1655.590 3524.800 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2026.140 2924.800 2027.340 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.610 3517.600 1620.170 3524.800 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 540.340 2.400 541.540 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.870 -4.800 1082.430 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 -4.800 171.170 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 482.540 2924.800 483.740 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1444.740 2924.800 1445.940 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 3517.600 138.970 3524.800 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2872.190 3517.600 2872.750 3524.800 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1781.340 2.400 1782.540 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2043.140 2.400 2044.340 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1941.140 2.400 1942.340 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 -4.800 132.530 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.230 -4.800 721.790 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2287.940 2924.800 2289.140 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 217.340 2.400 218.540 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.050 3517.600 1465.610 3524.800 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.930 3517.600 2283.490 3524.800 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2886.340 2.400 2887.540 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.930 -4.800 512.490 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2529.340 2924.800 2530.540 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.630 3517.600 2396.190 3524.800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1322.340 2.400 1323.540 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3148.140 2924.800 3149.340 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1546.740 2924.800 1547.940 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.310 3517.600 2054.870 3524.800 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.770 3517.600 100.330 3524.800 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2488.540 2924.800 2489.740 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2695.090 -4.800 2695.650 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1403.940 2924.800 1405.140 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1240.740 2.400 1241.940 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 502.940 2924.800 504.140 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.250 -4.800 531.810 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.490 -4.800 1633.050 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1866.340 2924.800 1867.540 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1999.570 3517.600 2000.130 3524.800 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3430.340 2924.800 3431.540 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 523.340 2924.800 524.540 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2308.340 2924.800 2309.540 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3471.140 2924.800 3472.340 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.290 3517.600 1922.850 3524.800 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 723.940 2924.800 725.140 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.690 3517.600 1826.250 3524.800 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.110 -4.800 2183.670 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 679.740 2.400 680.940 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.790 -4.800 2164.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 -4.800 0.510 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2543.750 -4.800 2544.310 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1281.540 2.400 1282.740 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2624.540 2.400 2625.740 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.410 3517.600 460.970 3524.800 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 839.540 2.400 840.740 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.270 -4.800 663.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.070 3517.600 1275.630 3524.800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.110 3517.600 573.670 3524.800 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.870 -4.800 1726.430 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.010 3517.600 1845.570 3524.800 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1203.340 2924.800 1204.540 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2022.740 2.400 2023.940 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2848.940 2924.800 2850.140 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.910 -4.800 702.470 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.890 -4.800 1214.450 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 179.940 2.400 181.140 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2709.540 2924.800 2710.740 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.850 -4.800 1916.410 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.270 3517.600 1790.830 3524.800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.950 3517.600 1771.510 3524.800 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3005.340 2.400 3006.540 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 3517.600 81.010 3524.800 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.490 -4.800 2277.050 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 700.140 2.400 701.340 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2706.140 2.400 2707.340 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1845.940 2924.800 1847.140 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 605.520 410.795 944.080 1288.405 ;
      LAYER met1 ;
        RECT 0.070 14.320 2913.570 3515.220 ;
      LAYER met2 ;
        RECT 0.100 3517.320 2.890 3518.050 ;
        RECT 4.010 3517.320 22.210 3518.050 ;
        RECT 23.330 3517.320 41.530 3518.050 ;
        RECT 42.650 3517.320 60.850 3518.050 ;
        RECT 61.970 3517.320 80.170 3518.050 ;
        RECT 81.290 3517.320 99.490 3518.050 ;
        RECT 100.610 3517.320 118.810 3518.050 ;
        RECT 119.930 3517.320 138.130 3518.050 ;
        RECT 139.250 3517.320 157.450 3518.050 ;
        RECT 158.570 3517.320 173.550 3518.050 ;
        RECT 174.670 3517.320 192.870 3518.050 ;
        RECT 193.990 3517.320 212.190 3518.050 ;
        RECT 213.310 3517.320 231.510 3518.050 ;
        RECT 232.630 3517.320 250.830 3518.050 ;
        RECT 251.950 3517.320 270.150 3518.050 ;
        RECT 271.270 3517.320 289.470 3518.050 ;
        RECT 290.590 3517.320 308.790 3518.050 ;
        RECT 309.910 3517.320 328.110 3518.050 ;
        RECT 329.230 3517.320 344.210 3518.050 ;
        RECT 345.330 3517.320 363.530 3518.050 ;
        RECT 364.650 3517.320 382.850 3518.050 ;
        RECT 383.970 3517.320 402.170 3518.050 ;
        RECT 403.290 3517.320 421.490 3518.050 ;
        RECT 422.610 3517.320 440.810 3518.050 ;
        RECT 441.930 3517.320 460.130 3518.050 ;
        RECT 461.250 3517.320 479.450 3518.050 ;
        RECT 480.570 3517.320 498.770 3518.050 ;
        RECT 499.890 3517.320 518.090 3518.050 ;
        RECT 519.210 3517.320 534.190 3518.050 ;
        RECT 535.310 3517.320 553.510 3518.050 ;
        RECT 554.630 3517.320 572.830 3518.050 ;
        RECT 573.950 3517.320 592.150 3518.050 ;
        RECT 593.270 3517.320 611.470 3518.050 ;
        RECT 612.590 3517.320 630.790 3518.050 ;
        RECT 631.910 3517.320 650.110 3518.050 ;
        RECT 651.230 3517.320 669.430 3518.050 ;
        RECT 670.550 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 708.070 3518.050 ;
        RECT 709.190 3517.320 724.170 3518.050 ;
        RECT 725.290 3517.320 743.490 3518.050 ;
        RECT 744.610 3517.320 762.810 3518.050 ;
        RECT 763.930 3517.320 782.130 3518.050 ;
        RECT 783.250 3517.320 801.450 3518.050 ;
        RECT 802.570 3517.320 820.770 3518.050 ;
        RECT 821.890 3517.320 840.090 3518.050 ;
        RECT 841.210 3517.320 859.410 3518.050 ;
        RECT 860.530 3517.320 878.730 3518.050 ;
        RECT 879.850 3517.320 894.830 3518.050 ;
        RECT 895.950 3517.320 914.150 3518.050 ;
        RECT 915.270 3517.320 933.470 3518.050 ;
        RECT 934.590 3517.320 952.790 3518.050 ;
        RECT 953.910 3517.320 972.110 3518.050 ;
        RECT 973.230 3517.320 991.430 3518.050 ;
        RECT 992.550 3517.320 1010.750 3518.050 ;
        RECT 1011.870 3517.320 1030.070 3518.050 ;
        RECT 1031.190 3517.320 1049.390 3518.050 ;
        RECT 1050.510 3517.320 1068.710 3518.050 ;
        RECT 1069.830 3517.320 1084.810 3518.050 ;
        RECT 1085.930 3517.320 1104.130 3518.050 ;
        RECT 1105.250 3517.320 1123.450 3518.050 ;
        RECT 1124.570 3517.320 1142.770 3518.050 ;
        RECT 1143.890 3517.320 1162.090 3518.050 ;
        RECT 1163.210 3517.320 1181.410 3518.050 ;
        RECT 1182.530 3517.320 1200.730 3518.050 ;
        RECT 1201.850 3517.320 1220.050 3518.050 ;
        RECT 1221.170 3517.320 1239.370 3518.050 ;
        RECT 1240.490 3517.320 1258.690 3518.050 ;
        RECT 1259.810 3517.320 1274.790 3518.050 ;
        RECT 1275.910 3517.320 1294.110 3518.050 ;
        RECT 1295.230 3517.320 1313.430 3518.050 ;
        RECT 1314.550 3517.320 1332.750 3518.050 ;
        RECT 1333.870 3517.320 1352.070 3518.050 ;
        RECT 1353.190 3517.320 1371.390 3518.050 ;
        RECT 1372.510 3517.320 1390.710 3518.050 ;
        RECT 1391.830 3517.320 1410.030 3518.050 ;
        RECT 1411.150 3517.320 1429.350 3518.050 ;
        RECT 1430.470 3517.320 1445.450 3518.050 ;
        RECT 1446.570 3517.320 1464.770 3518.050 ;
        RECT 1465.890 3517.320 1484.090 3518.050 ;
        RECT 1485.210 3517.320 1503.410 3518.050 ;
        RECT 1504.530 3517.320 1522.730 3518.050 ;
        RECT 1523.850 3517.320 1542.050 3518.050 ;
        RECT 1543.170 3517.320 1561.370 3518.050 ;
        RECT 1562.490 3517.320 1580.690 3518.050 ;
        RECT 1581.810 3517.320 1600.010 3518.050 ;
        RECT 1601.130 3517.320 1619.330 3518.050 ;
        RECT 1620.450 3517.320 1635.430 3518.050 ;
        RECT 1636.550 3517.320 1654.750 3518.050 ;
        RECT 1655.870 3517.320 1674.070 3518.050 ;
        RECT 1675.190 3517.320 1693.390 3518.050 ;
        RECT 1694.510 3517.320 1712.710 3518.050 ;
        RECT 1713.830 3517.320 1732.030 3518.050 ;
        RECT 1733.150 3517.320 1751.350 3518.050 ;
        RECT 1752.470 3517.320 1770.670 3518.050 ;
        RECT 1771.790 3517.320 1789.990 3518.050 ;
        RECT 1791.110 3517.320 1809.310 3518.050 ;
        RECT 1810.430 3517.320 1825.410 3518.050 ;
        RECT 1826.530 3517.320 1844.730 3518.050 ;
        RECT 1845.850 3517.320 1864.050 3518.050 ;
        RECT 1865.170 3517.320 1883.370 3518.050 ;
        RECT 1884.490 3517.320 1902.690 3518.050 ;
        RECT 1903.810 3517.320 1922.010 3518.050 ;
        RECT 1923.130 3517.320 1941.330 3518.050 ;
        RECT 1942.450 3517.320 1960.650 3518.050 ;
        RECT 1961.770 3517.320 1979.970 3518.050 ;
        RECT 1981.090 3517.320 1999.290 3518.050 ;
        RECT 2000.410 3517.320 2015.390 3518.050 ;
        RECT 2016.510 3517.320 2034.710 3518.050 ;
        RECT 2035.830 3517.320 2054.030 3518.050 ;
        RECT 2055.150 3517.320 2073.350 3518.050 ;
        RECT 2074.470 3517.320 2092.670 3518.050 ;
        RECT 2093.790 3517.320 2111.990 3518.050 ;
        RECT 2113.110 3517.320 2131.310 3518.050 ;
        RECT 2132.430 3517.320 2150.630 3518.050 ;
        RECT 2151.750 3517.320 2169.950 3518.050 ;
        RECT 2171.070 3517.320 2186.050 3518.050 ;
        RECT 2187.170 3517.320 2205.370 3518.050 ;
        RECT 2206.490 3517.320 2224.690 3518.050 ;
        RECT 2225.810 3517.320 2244.010 3518.050 ;
        RECT 2245.130 3517.320 2263.330 3518.050 ;
        RECT 2264.450 3517.320 2282.650 3518.050 ;
        RECT 2283.770 3517.320 2301.970 3518.050 ;
        RECT 2303.090 3517.320 2321.290 3518.050 ;
        RECT 2322.410 3517.320 2340.610 3518.050 ;
        RECT 2341.730 3517.320 2359.930 3518.050 ;
        RECT 2361.050 3517.320 2376.030 3518.050 ;
        RECT 2377.150 3517.320 2395.350 3518.050 ;
        RECT 2396.470 3517.320 2414.670 3518.050 ;
        RECT 2415.790 3517.320 2433.990 3518.050 ;
        RECT 2435.110 3517.320 2453.310 3518.050 ;
        RECT 2454.430 3517.320 2472.630 3518.050 ;
        RECT 2473.750 3517.320 2491.950 3518.050 ;
        RECT 2493.070 3517.320 2511.270 3518.050 ;
        RECT 2512.390 3517.320 2530.590 3518.050 ;
        RECT 2531.710 3517.320 2549.910 3518.050 ;
        RECT 2551.030 3517.320 2566.010 3518.050 ;
        RECT 2567.130 3517.320 2585.330 3518.050 ;
        RECT 2586.450 3517.320 2604.650 3518.050 ;
        RECT 2605.770 3517.320 2623.970 3518.050 ;
        RECT 2625.090 3517.320 2643.290 3518.050 ;
        RECT 2644.410 3517.320 2662.610 3518.050 ;
        RECT 2663.730 3517.320 2681.930 3518.050 ;
        RECT 2683.050 3517.320 2701.250 3518.050 ;
        RECT 2702.370 3517.320 2720.570 3518.050 ;
        RECT 2721.690 3517.320 2736.670 3518.050 ;
        RECT 2737.790 3517.320 2755.990 3518.050 ;
        RECT 2757.110 3517.320 2775.310 3518.050 ;
        RECT 2776.430 3517.320 2794.630 3518.050 ;
        RECT 2795.750 3517.320 2813.950 3518.050 ;
        RECT 2815.070 3517.320 2833.270 3518.050 ;
        RECT 2834.390 3517.320 2852.590 3518.050 ;
        RECT 2853.710 3517.320 2871.910 3518.050 ;
        RECT 2873.030 3517.320 2891.230 3518.050 ;
        RECT 2892.350 3517.320 2910.550 3518.050 ;
        RECT 2911.670 3517.320 2914.470 3518.050 ;
        RECT 0.100 2.680 2914.470 3517.320 ;
        RECT 0.790 1.630 15.770 2.680 ;
        RECT 16.890 1.630 35.090 2.680 ;
        RECT 36.210 1.630 54.410 2.680 ;
        RECT 55.530 1.630 73.730 2.680 ;
        RECT 74.850 1.630 93.050 2.680 ;
        RECT 94.170 1.630 112.370 2.680 ;
        RECT 113.490 1.630 131.690 2.680 ;
        RECT 132.810 1.630 151.010 2.680 ;
        RECT 152.130 1.630 170.330 2.680 ;
        RECT 171.450 1.630 186.430 2.680 ;
        RECT 187.550 1.630 205.750 2.680 ;
        RECT 206.870 1.630 225.070 2.680 ;
        RECT 226.190 1.630 244.390 2.680 ;
        RECT 245.510 1.630 263.710 2.680 ;
        RECT 264.830 1.630 283.030 2.680 ;
        RECT 284.150 1.630 302.350 2.680 ;
        RECT 303.470 1.630 321.670 2.680 ;
        RECT 322.790 1.630 340.990 2.680 ;
        RECT 342.110 1.630 360.310 2.680 ;
        RECT 361.430 1.630 376.410 2.680 ;
        RECT 377.530 1.630 395.730 2.680 ;
        RECT 396.850 1.630 415.050 2.680 ;
        RECT 416.170 1.630 434.370 2.680 ;
        RECT 435.490 1.630 453.690 2.680 ;
        RECT 454.810 1.630 473.010 2.680 ;
        RECT 474.130 1.630 492.330 2.680 ;
        RECT 493.450 1.630 511.650 2.680 ;
        RECT 512.770 1.630 530.970 2.680 ;
        RECT 532.090 1.630 550.290 2.680 ;
        RECT 551.410 1.630 566.390 2.680 ;
        RECT 567.510 1.630 585.710 2.680 ;
        RECT 586.830 1.630 605.030 2.680 ;
        RECT 606.150 1.630 624.350 2.680 ;
        RECT 625.470 1.630 643.670 2.680 ;
        RECT 644.790 1.630 662.990 2.680 ;
        RECT 664.110 1.630 682.310 2.680 ;
        RECT 683.430 1.630 701.630 2.680 ;
        RECT 702.750 1.630 720.950 2.680 ;
        RECT 722.070 1.630 737.050 2.680 ;
        RECT 738.170 1.630 756.370 2.680 ;
        RECT 757.490 1.630 775.690 2.680 ;
        RECT 776.810 1.630 795.010 2.680 ;
        RECT 796.130 1.630 814.330 2.680 ;
        RECT 815.450 1.630 833.650 2.680 ;
        RECT 834.770 1.630 852.970 2.680 ;
        RECT 854.090 1.630 872.290 2.680 ;
        RECT 873.410 1.630 891.610 2.680 ;
        RECT 892.730 1.630 910.930 2.680 ;
        RECT 912.050 1.630 927.030 2.680 ;
        RECT 928.150 1.630 946.350 2.680 ;
        RECT 947.470 1.630 965.670 2.680 ;
        RECT 966.790 1.630 984.990 2.680 ;
        RECT 986.110 1.630 1004.310 2.680 ;
        RECT 1005.430 1.630 1023.630 2.680 ;
        RECT 1024.750 1.630 1042.950 2.680 ;
        RECT 1044.070 1.630 1062.270 2.680 ;
        RECT 1063.390 1.630 1081.590 2.680 ;
        RECT 1082.710 1.630 1100.910 2.680 ;
        RECT 1102.030 1.630 1117.010 2.680 ;
        RECT 1118.130 1.630 1136.330 2.680 ;
        RECT 1137.450 1.630 1155.650 2.680 ;
        RECT 1156.770 1.630 1174.970 2.680 ;
        RECT 1176.090 1.630 1194.290 2.680 ;
        RECT 1195.410 1.630 1213.610 2.680 ;
        RECT 1214.730 1.630 1232.930 2.680 ;
        RECT 1234.050 1.630 1252.250 2.680 ;
        RECT 1253.370 1.630 1271.570 2.680 ;
        RECT 1272.690 1.630 1287.670 2.680 ;
        RECT 1288.790 1.630 1306.990 2.680 ;
        RECT 1308.110 1.630 1326.310 2.680 ;
        RECT 1327.430 1.630 1345.630 2.680 ;
        RECT 1346.750 1.630 1364.950 2.680 ;
        RECT 1366.070 1.630 1384.270 2.680 ;
        RECT 1385.390 1.630 1403.590 2.680 ;
        RECT 1404.710 1.630 1422.910 2.680 ;
        RECT 1424.030 1.630 1442.230 2.680 ;
        RECT 1443.350 1.630 1461.550 2.680 ;
        RECT 1462.670 1.630 1477.650 2.680 ;
        RECT 1478.770 1.630 1496.970 2.680 ;
        RECT 1498.090 1.630 1516.290 2.680 ;
        RECT 1517.410 1.630 1535.610 2.680 ;
        RECT 1536.730 1.630 1554.930 2.680 ;
        RECT 1556.050 1.630 1574.250 2.680 ;
        RECT 1575.370 1.630 1593.570 2.680 ;
        RECT 1594.690 1.630 1612.890 2.680 ;
        RECT 1614.010 1.630 1632.210 2.680 ;
        RECT 1633.330 1.630 1651.530 2.680 ;
        RECT 1652.650 1.630 1667.630 2.680 ;
        RECT 1668.750 1.630 1686.950 2.680 ;
        RECT 1688.070 1.630 1706.270 2.680 ;
        RECT 1707.390 1.630 1725.590 2.680 ;
        RECT 1726.710 1.630 1744.910 2.680 ;
        RECT 1746.030 1.630 1764.230 2.680 ;
        RECT 1765.350 1.630 1783.550 2.680 ;
        RECT 1784.670 1.630 1802.870 2.680 ;
        RECT 1803.990 1.630 1822.190 2.680 ;
        RECT 1823.310 1.630 1838.290 2.680 ;
        RECT 1839.410 1.630 1857.610 2.680 ;
        RECT 1858.730 1.630 1876.930 2.680 ;
        RECT 1878.050 1.630 1896.250 2.680 ;
        RECT 1897.370 1.630 1915.570 2.680 ;
        RECT 1916.690 1.630 1934.890 2.680 ;
        RECT 1936.010 1.630 1954.210 2.680 ;
        RECT 1955.330 1.630 1973.530 2.680 ;
        RECT 1974.650 1.630 1992.850 2.680 ;
        RECT 1993.970 1.630 2012.170 2.680 ;
        RECT 2013.290 1.630 2028.270 2.680 ;
        RECT 2029.390 1.630 2047.590 2.680 ;
        RECT 2048.710 1.630 2066.910 2.680 ;
        RECT 2068.030 1.630 2086.230 2.680 ;
        RECT 2087.350 1.630 2105.550 2.680 ;
        RECT 2106.670 1.630 2124.870 2.680 ;
        RECT 2125.990 1.630 2144.190 2.680 ;
        RECT 2145.310 1.630 2163.510 2.680 ;
        RECT 2164.630 1.630 2182.830 2.680 ;
        RECT 2183.950 1.630 2202.150 2.680 ;
        RECT 2203.270 1.630 2218.250 2.680 ;
        RECT 2219.370 1.630 2237.570 2.680 ;
        RECT 2238.690 1.630 2256.890 2.680 ;
        RECT 2258.010 1.630 2276.210 2.680 ;
        RECT 2277.330 1.630 2295.530 2.680 ;
        RECT 2296.650 1.630 2314.850 2.680 ;
        RECT 2315.970 1.630 2334.170 2.680 ;
        RECT 2335.290 1.630 2353.490 2.680 ;
        RECT 2354.610 1.630 2372.810 2.680 ;
        RECT 2373.930 1.630 2388.910 2.680 ;
        RECT 2390.030 1.630 2408.230 2.680 ;
        RECT 2409.350 1.630 2427.550 2.680 ;
        RECT 2428.670 1.630 2446.870 2.680 ;
        RECT 2447.990 1.630 2466.190 2.680 ;
        RECT 2467.310 1.630 2485.510 2.680 ;
        RECT 2486.630 1.630 2504.830 2.680 ;
        RECT 2505.950 1.630 2524.150 2.680 ;
        RECT 2525.270 1.630 2543.470 2.680 ;
        RECT 2544.590 1.630 2562.790 2.680 ;
        RECT 2563.910 1.630 2578.890 2.680 ;
        RECT 2580.010 1.630 2598.210 2.680 ;
        RECT 2599.330 1.630 2617.530 2.680 ;
        RECT 2618.650 1.630 2636.850 2.680 ;
        RECT 2637.970 1.630 2656.170 2.680 ;
        RECT 2657.290 1.630 2675.490 2.680 ;
        RECT 2676.610 1.630 2694.810 2.680 ;
        RECT 2695.930 1.630 2714.130 2.680 ;
        RECT 2715.250 1.630 2733.450 2.680 ;
        RECT 2734.570 1.630 2752.770 2.680 ;
        RECT 2753.890 1.630 2768.870 2.680 ;
        RECT 2769.990 1.630 2788.190 2.680 ;
        RECT 2789.310 1.630 2807.510 2.680 ;
        RECT 2808.630 1.630 2826.830 2.680 ;
        RECT 2827.950 1.630 2846.150 2.680 ;
        RECT 2847.270 1.630 2865.470 2.680 ;
        RECT 2866.590 1.630 2884.790 2.680 ;
        RECT 2885.910 1.630 2904.110 2.680 ;
        RECT 2905.230 1.630 2914.470 2.680 ;
      LAYER met3 ;
        RECT 1.230 3511.540 2917.200 3512.705 ;
        RECT 1.230 3506.740 2917.930 3511.540 ;
        RECT 2.800 3504.740 2917.930 3506.740 ;
        RECT 1.230 3493.140 2917.930 3504.740 ;
        RECT 1.230 3491.140 2917.200 3493.140 ;
        RECT 1.230 3489.740 2917.930 3491.140 ;
        RECT 2.800 3487.740 2917.930 3489.740 ;
        RECT 1.230 3472.740 2917.930 3487.740 ;
        RECT 1.230 3470.740 2917.200 3472.740 ;
        RECT 1.230 3469.340 2917.930 3470.740 ;
        RECT 2.800 3467.340 2917.930 3469.340 ;
        RECT 1.230 3452.340 2917.930 3467.340 ;
        RECT 1.230 3450.340 2917.200 3452.340 ;
        RECT 1.230 3448.940 2917.930 3450.340 ;
        RECT 2.800 3446.940 2917.930 3448.940 ;
        RECT 1.230 3431.940 2917.930 3446.940 ;
        RECT 1.230 3429.940 2917.200 3431.940 ;
        RECT 1.230 3428.540 2917.930 3429.940 ;
        RECT 2.800 3426.540 2917.930 3428.540 ;
        RECT 1.230 3411.540 2917.930 3426.540 ;
        RECT 1.230 3409.540 2917.200 3411.540 ;
        RECT 1.230 3408.140 2917.930 3409.540 ;
        RECT 2.800 3406.140 2917.930 3408.140 ;
        RECT 1.230 3391.140 2917.930 3406.140 ;
        RECT 1.230 3389.140 2917.200 3391.140 ;
        RECT 1.230 3387.740 2917.930 3389.140 ;
        RECT 2.800 3385.740 2917.930 3387.740 ;
        RECT 1.230 3370.740 2917.930 3385.740 ;
        RECT 1.230 3368.740 2917.200 3370.740 ;
        RECT 1.230 3367.340 2917.930 3368.740 ;
        RECT 2.800 3365.340 2917.930 3367.340 ;
        RECT 1.230 3350.340 2917.930 3365.340 ;
        RECT 1.230 3348.340 2917.200 3350.340 ;
        RECT 1.230 3346.940 2917.930 3348.340 ;
        RECT 2.800 3344.940 2917.930 3346.940 ;
        RECT 1.230 3329.940 2917.930 3344.940 ;
        RECT 1.230 3327.940 2917.200 3329.940 ;
        RECT 1.230 3326.540 2917.930 3327.940 ;
        RECT 2.800 3324.540 2917.930 3326.540 ;
        RECT 1.230 3312.940 2917.930 3324.540 ;
        RECT 1.230 3310.940 2917.200 3312.940 ;
        RECT 1.230 3306.140 2917.930 3310.940 ;
        RECT 2.800 3304.140 2917.930 3306.140 ;
        RECT 1.230 3292.540 2917.930 3304.140 ;
        RECT 1.230 3290.540 2917.200 3292.540 ;
        RECT 1.230 3289.140 2917.930 3290.540 ;
        RECT 2.800 3287.140 2917.930 3289.140 ;
        RECT 1.230 3272.140 2917.930 3287.140 ;
        RECT 1.230 3270.140 2917.200 3272.140 ;
        RECT 1.230 3268.740 2917.930 3270.140 ;
        RECT 2.800 3266.740 2917.930 3268.740 ;
        RECT 1.230 3251.740 2917.930 3266.740 ;
        RECT 1.230 3249.740 2917.200 3251.740 ;
        RECT 1.230 3248.340 2917.930 3249.740 ;
        RECT 2.800 3246.340 2917.930 3248.340 ;
        RECT 1.230 3231.340 2917.930 3246.340 ;
        RECT 1.230 3229.340 2917.200 3231.340 ;
        RECT 1.230 3227.940 2917.930 3229.340 ;
        RECT 2.800 3225.940 2917.930 3227.940 ;
        RECT 1.230 3210.940 2917.930 3225.940 ;
        RECT 1.230 3208.940 2917.200 3210.940 ;
        RECT 1.230 3207.540 2917.930 3208.940 ;
        RECT 2.800 3205.540 2917.930 3207.540 ;
        RECT 1.230 3190.540 2917.930 3205.540 ;
        RECT 1.230 3188.540 2917.200 3190.540 ;
        RECT 1.230 3187.140 2917.930 3188.540 ;
        RECT 2.800 3185.140 2917.930 3187.140 ;
        RECT 1.230 3170.140 2917.930 3185.140 ;
        RECT 1.230 3168.140 2917.200 3170.140 ;
        RECT 1.230 3166.740 2917.930 3168.140 ;
        RECT 2.800 3164.740 2917.930 3166.740 ;
        RECT 1.230 3149.740 2917.930 3164.740 ;
        RECT 1.230 3147.740 2917.200 3149.740 ;
        RECT 1.230 3146.340 2917.930 3147.740 ;
        RECT 2.800 3144.340 2917.930 3146.340 ;
        RECT 1.230 3132.740 2917.930 3144.340 ;
        RECT 1.230 3130.740 2917.200 3132.740 ;
        RECT 1.230 3125.940 2917.930 3130.740 ;
        RECT 2.800 3123.940 2917.930 3125.940 ;
        RECT 1.230 3112.340 2917.930 3123.940 ;
        RECT 1.230 3110.340 2917.200 3112.340 ;
        RECT 1.230 3108.940 2917.930 3110.340 ;
        RECT 2.800 3106.940 2917.930 3108.940 ;
        RECT 1.230 3091.940 2917.930 3106.940 ;
        RECT 1.230 3089.940 2917.200 3091.940 ;
        RECT 1.230 3088.540 2917.930 3089.940 ;
        RECT 2.800 3086.540 2917.930 3088.540 ;
        RECT 1.230 3071.540 2917.930 3086.540 ;
        RECT 1.230 3069.540 2917.200 3071.540 ;
        RECT 1.230 3068.140 2917.930 3069.540 ;
        RECT 2.800 3066.140 2917.930 3068.140 ;
        RECT 1.230 3051.140 2917.930 3066.140 ;
        RECT 1.230 3049.140 2917.200 3051.140 ;
        RECT 1.230 3047.740 2917.930 3049.140 ;
        RECT 2.800 3045.740 2917.930 3047.740 ;
        RECT 1.230 3030.740 2917.930 3045.740 ;
        RECT 1.230 3028.740 2917.200 3030.740 ;
        RECT 1.230 3027.340 2917.930 3028.740 ;
        RECT 2.800 3025.340 2917.930 3027.340 ;
        RECT 1.230 3010.340 2917.930 3025.340 ;
        RECT 1.230 3008.340 2917.200 3010.340 ;
        RECT 1.230 3006.940 2917.930 3008.340 ;
        RECT 2.800 3004.940 2917.930 3006.940 ;
        RECT 1.230 2989.940 2917.930 3004.940 ;
        RECT 1.230 2987.940 2917.200 2989.940 ;
        RECT 1.230 2986.540 2917.930 2987.940 ;
        RECT 2.800 2984.540 2917.930 2986.540 ;
        RECT 1.230 2969.540 2917.930 2984.540 ;
        RECT 1.230 2967.540 2917.200 2969.540 ;
        RECT 1.230 2966.140 2917.930 2967.540 ;
        RECT 2.800 2964.140 2917.930 2966.140 ;
        RECT 1.230 2949.140 2917.930 2964.140 ;
        RECT 1.230 2947.140 2917.200 2949.140 ;
        RECT 1.230 2945.740 2917.930 2947.140 ;
        RECT 2.800 2943.740 2917.930 2945.740 ;
        RECT 1.230 2932.140 2917.930 2943.740 ;
        RECT 1.230 2930.140 2917.200 2932.140 ;
        RECT 1.230 2925.340 2917.930 2930.140 ;
        RECT 2.800 2923.340 2917.930 2925.340 ;
        RECT 1.230 2911.740 2917.930 2923.340 ;
        RECT 1.230 2909.740 2917.200 2911.740 ;
        RECT 1.230 2908.340 2917.930 2909.740 ;
        RECT 2.800 2906.340 2917.930 2908.340 ;
        RECT 1.230 2891.340 2917.930 2906.340 ;
        RECT 1.230 2889.340 2917.200 2891.340 ;
        RECT 1.230 2887.940 2917.930 2889.340 ;
        RECT 2.800 2885.940 2917.930 2887.940 ;
        RECT 1.230 2870.940 2917.930 2885.940 ;
        RECT 1.230 2868.940 2917.200 2870.940 ;
        RECT 1.230 2867.540 2917.930 2868.940 ;
        RECT 2.800 2865.540 2917.930 2867.540 ;
        RECT 1.230 2850.540 2917.930 2865.540 ;
        RECT 1.230 2848.540 2917.200 2850.540 ;
        RECT 1.230 2847.140 2917.930 2848.540 ;
        RECT 2.800 2845.140 2917.930 2847.140 ;
        RECT 1.230 2830.140 2917.930 2845.140 ;
        RECT 1.230 2828.140 2917.200 2830.140 ;
        RECT 1.230 2826.740 2917.930 2828.140 ;
        RECT 2.800 2824.740 2917.930 2826.740 ;
        RECT 1.230 2809.740 2917.930 2824.740 ;
        RECT 1.230 2807.740 2917.200 2809.740 ;
        RECT 1.230 2806.340 2917.930 2807.740 ;
        RECT 2.800 2804.340 2917.930 2806.340 ;
        RECT 1.230 2789.340 2917.930 2804.340 ;
        RECT 1.230 2787.340 2917.200 2789.340 ;
        RECT 1.230 2785.940 2917.930 2787.340 ;
        RECT 2.800 2783.940 2917.930 2785.940 ;
        RECT 1.230 2768.940 2917.930 2783.940 ;
        RECT 1.230 2766.940 2917.200 2768.940 ;
        RECT 1.230 2765.540 2917.930 2766.940 ;
        RECT 2.800 2763.540 2917.930 2765.540 ;
        RECT 1.230 2748.540 2917.930 2763.540 ;
        RECT 1.230 2746.540 2917.200 2748.540 ;
        RECT 1.230 2745.140 2917.930 2746.540 ;
        RECT 2.800 2743.140 2917.930 2745.140 ;
        RECT 1.230 2731.540 2917.930 2743.140 ;
        RECT 1.230 2729.540 2917.200 2731.540 ;
        RECT 1.230 2724.740 2917.930 2729.540 ;
        RECT 2.800 2722.740 2917.930 2724.740 ;
        RECT 1.230 2711.140 2917.930 2722.740 ;
        RECT 1.230 2709.140 2917.200 2711.140 ;
        RECT 1.230 2707.740 2917.930 2709.140 ;
        RECT 2.800 2705.740 2917.930 2707.740 ;
        RECT 1.230 2690.740 2917.930 2705.740 ;
        RECT 1.230 2688.740 2917.200 2690.740 ;
        RECT 1.230 2687.340 2917.930 2688.740 ;
        RECT 2.800 2685.340 2917.930 2687.340 ;
        RECT 1.230 2670.340 2917.930 2685.340 ;
        RECT 1.230 2668.340 2917.200 2670.340 ;
        RECT 1.230 2666.940 2917.930 2668.340 ;
        RECT 2.800 2664.940 2917.930 2666.940 ;
        RECT 1.230 2649.940 2917.930 2664.940 ;
        RECT 1.230 2647.940 2917.200 2649.940 ;
        RECT 1.230 2646.540 2917.930 2647.940 ;
        RECT 2.800 2644.540 2917.930 2646.540 ;
        RECT 1.230 2629.540 2917.930 2644.540 ;
        RECT 1.230 2627.540 2917.200 2629.540 ;
        RECT 1.230 2626.140 2917.930 2627.540 ;
        RECT 2.800 2624.140 2917.930 2626.140 ;
        RECT 1.230 2609.140 2917.930 2624.140 ;
        RECT 1.230 2607.140 2917.200 2609.140 ;
        RECT 1.230 2605.740 2917.930 2607.140 ;
        RECT 2.800 2603.740 2917.930 2605.740 ;
        RECT 1.230 2588.740 2917.930 2603.740 ;
        RECT 1.230 2586.740 2917.200 2588.740 ;
        RECT 1.230 2585.340 2917.930 2586.740 ;
        RECT 2.800 2583.340 2917.930 2585.340 ;
        RECT 1.230 2568.340 2917.930 2583.340 ;
        RECT 1.230 2566.340 2917.200 2568.340 ;
        RECT 1.230 2564.940 2917.930 2566.340 ;
        RECT 2.800 2562.940 2917.930 2564.940 ;
        RECT 1.230 2551.340 2917.930 2562.940 ;
        RECT 1.230 2549.340 2917.200 2551.340 ;
        RECT 1.230 2544.540 2917.930 2549.340 ;
        RECT 2.800 2542.540 2917.930 2544.540 ;
        RECT 1.230 2530.940 2917.930 2542.540 ;
        RECT 1.230 2528.940 2917.200 2530.940 ;
        RECT 1.230 2524.140 2917.930 2528.940 ;
        RECT 2.800 2522.140 2917.930 2524.140 ;
        RECT 1.230 2510.540 2917.930 2522.140 ;
        RECT 1.230 2508.540 2917.200 2510.540 ;
        RECT 1.230 2507.140 2917.930 2508.540 ;
        RECT 2.800 2505.140 2917.930 2507.140 ;
        RECT 1.230 2490.140 2917.930 2505.140 ;
        RECT 1.230 2488.140 2917.200 2490.140 ;
        RECT 1.230 2486.740 2917.930 2488.140 ;
        RECT 2.800 2484.740 2917.930 2486.740 ;
        RECT 1.230 2469.740 2917.930 2484.740 ;
        RECT 1.230 2467.740 2917.200 2469.740 ;
        RECT 1.230 2466.340 2917.930 2467.740 ;
        RECT 2.800 2464.340 2917.930 2466.340 ;
        RECT 1.230 2449.340 2917.930 2464.340 ;
        RECT 1.230 2447.340 2917.200 2449.340 ;
        RECT 1.230 2445.940 2917.930 2447.340 ;
        RECT 2.800 2443.940 2917.930 2445.940 ;
        RECT 1.230 2428.940 2917.930 2443.940 ;
        RECT 1.230 2426.940 2917.200 2428.940 ;
        RECT 1.230 2425.540 2917.930 2426.940 ;
        RECT 2.800 2423.540 2917.930 2425.540 ;
        RECT 1.230 2408.540 2917.930 2423.540 ;
        RECT 1.230 2406.540 2917.200 2408.540 ;
        RECT 1.230 2405.140 2917.930 2406.540 ;
        RECT 2.800 2403.140 2917.930 2405.140 ;
        RECT 1.230 2388.140 2917.930 2403.140 ;
        RECT 1.230 2386.140 2917.200 2388.140 ;
        RECT 1.230 2384.740 2917.930 2386.140 ;
        RECT 2.800 2382.740 2917.930 2384.740 ;
        RECT 1.230 2367.740 2917.930 2382.740 ;
        RECT 1.230 2365.740 2917.200 2367.740 ;
        RECT 1.230 2364.340 2917.930 2365.740 ;
        RECT 2.800 2362.340 2917.930 2364.340 ;
        RECT 1.230 2350.740 2917.930 2362.340 ;
        RECT 1.230 2348.740 2917.200 2350.740 ;
        RECT 1.230 2343.940 2917.930 2348.740 ;
        RECT 2.800 2341.940 2917.930 2343.940 ;
        RECT 1.230 2330.340 2917.930 2341.940 ;
        RECT 1.230 2328.340 2917.200 2330.340 ;
        RECT 1.230 2326.940 2917.930 2328.340 ;
        RECT 2.800 2324.940 2917.930 2326.940 ;
        RECT 1.230 2309.940 2917.930 2324.940 ;
        RECT 1.230 2307.940 2917.200 2309.940 ;
        RECT 1.230 2306.540 2917.930 2307.940 ;
        RECT 2.800 2304.540 2917.930 2306.540 ;
        RECT 1.230 2289.540 2917.930 2304.540 ;
        RECT 1.230 2287.540 2917.200 2289.540 ;
        RECT 1.230 2286.140 2917.930 2287.540 ;
        RECT 2.800 2284.140 2917.930 2286.140 ;
        RECT 1.230 2269.140 2917.930 2284.140 ;
        RECT 1.230 2267.140 2917.200 2269.140 ;
        RECT 1.230 2265.740 2917.930 2267.140 ;
        RECT 2.800 2263.740 2917.930 2265.740 ;
        RECT 1.230 2248.740 2917.930 2263.740 ;
        RECT 1.230 2246.740 2917.200 2248.740 ;
        RECT 1.230 2245.340 2917.930 2246.740 ;
        RECT 2.800 2243.340 2917.930 2245.340 ;
        RECT 1.230 2228.340 2917.930 2243.340 ;
        RECT 1.230 2226.340 2917.200 2228.340 ;
        RECT 1.230 2224.940 2917.930 2226.340 ;
        RECT 2.800 2222.940 2917.930 2224.940 ;
        RECT 1.230 2207.940 2917.930 2222.940 ;
        RECT 1.230 2205.940 2917.200 2207.940 ;
        RECT 1.230 2204.540 2917.930 2205.940 ;
        RECT 2.800 2202.540 2917.930 2204.540 ;
        RECT 1.230 2187.540 2917.930 2202.540 ;
        RECT 1.230 2185.540 2917.200 2187.540 ;
        RECT 1.230 2184.140 2917.930 2185.540 ;
        RECT 2.800 2182.140 2917.930 2184.140 ;
        RECT 1.230 2167.140 2917.930 2182.140 ;
        RECT 1.230 2165.140 2917.200 2167.140 ;
        RECT 1.230 2163.740 2917.930 2165.140 ;
        RECT 2.800 2161.740 2917.930 2163.740 ;
        RECT 1.230 2150.140 2917.930 2161.740 ;
        RECT 1.230 2148.140 2917.200 2150.140 ;
        RECT 1.230 2143.340 2917.930 2148.140 ;
        RECT 2.800 2141.340 2917.930 2143.340 ;
        RECT 1.230 2129.740 2917.930 2141.340 ;
        RECT 1.230 2127.740 2917.200 2129.740 ;
        RECT 1.230 2126.340 2917.930 2127.740 ;
        RECT 2.800 2124.340 2917.930 2126.340 ;
        RECT 1.230 2109.340 2917.930 2124.340 ;
        RECT 1.230 2107.340 2917.200 2109.340 ;
        RECT 1.230 2105.940 2917.930 2107.340 ;
        RECT 2.800 2103.940 2917.930 2105.940 ;
        RECT 1.230 2088.940 2917.930 2103.940 ;
        RECT 1.230 2086.940 2917.200 2088.940 ;
        RECT 1.230 2085.540 2917.930 2086.940 ;
        RECT 2.800 2083.540 2917.930 2085.540 ;
        RECT 1.230 2068.540 2917.930 2083.540 ;
        RECT 1.230 2066.540 2917.200 2068.540 ;
        RECT 1.230 2065.140 2917.930 2066.540 ;
        RECT 2.800 2063.140 2917.930 2065.140 ;
        RECT 1.230 2048.140 2917.930 2063.140 ;
        RECT 1.230 2046.140 2917.200 2048.140 ;
        RECT 1.230 2044.740 2917.930 2046.140 ;
        RECT 2.800 2042.740 2917.930 2044.740 ;
        RECT 1.230 2027.740 2917.930 2042.740 ;
        RECT 1.230 2025.740 2917.200 2027.740 ;
        RECT 1.230 2024.340 2917.930 2025.740 ;
        RECT 2.800 2022.340 2917.930 2024.340 ;
        RECT 1.230 2007.340 2917.930 2022.340 ;
        RECT 1.230 2005.340 2917.200 2007.340 ;
        RECT 1.230 2003.940 2917.930 2005.340 ;
        RECT 2.800 2001.940 2917.930 2003.940 ;
        RECT 1.230 1986.940 2917.930 2001.940 ;
        RECT 1.230 1984.940 2917.200 1986.940 ;
        RECT 1.230 1983.540 2917.930 1984.940 ;
        RECT 2.800 1981.540 2917.930 1983.540 ;
        RECT 1.230 1966.540 2917.930 1981.540 ;
        RECT 1.230 1964.540 2917.200 1966.540 ;
        RECT 1.230 1963.140 2917.930 1964.540 ;
        RECT 2.800 1961.140 2917.930 1963.140 ;
        RECT 1.230 1949.540 2917.930 1961.140 ;
        RECT 1.230 1947.540 2917.200 1949.540 ;
        RECT 1.230 1942.740 2917.930 1947.540 ;
        RECT 2.800 1940.740 2917.930 1942.740 ;
        RECT 1.230 1929.140 2917.930 1940.740 ;
        RECT 1.230 1927.140 2917.200 1929.140 ;
        RECT 1.230 1925.740 2917.930 1927.140 ;
        RECT 2.800 1923.740 2917.930 1925.740 ;
        RECT 1.230 1908.740 2917.930 1923.740 ;
        RECT 1.230 1906.740 2917.200 1908.740 ;
        RECT 1.230 1905.340 2917.930 1906.740 ;
        RECT 2.800 1903.340 2917.930 1905.340 ;
        RECT 1.230 1888.340 2917.930 1903.340 ;
        RECT 1.230 1886.340 2917.200 1888.340 ;
        RECT 1.230 1884.940 2917.930 1886.340 ;
        RECT 2.800 1882.940 2917.930 1884.940 ;
        RECT 1.230 1867.940 2917.930 1882.940 ;
        RECT 1.230 1865.940 2917.200 1867.940 ;
        RECT 1.230 1864.540 2917.930 1865.940 ;
        RECT 2.800 1862.540 2917.930 1864.540 ;
        RECT 1.230 1847.540 2917.930 1862.540 ;
        RECT 1.230 1845.540 2917.200 1847.540 ;
        RECT 1.230 1844.140 2917.930 1845.540 ;
        RECT 2.800 1842.140 2917.930 1844.140 ;
        RECT 1.230 1827.140 2917.930 1842.140 ;
        RECT 1.230 1825.140 2917.200 1827.140 ;
        RECT 1.230 1823.740 2917.930 1825.140 ;
        RECT 2.800 1821.740 2917.930 1823.740 ;
        RECT 1.230 1806.740 2917.930 1821.740 ;
        RECT 1.230 1804.740 2917.200 1806.740 ;
        RECT 1.230 1803.340 2917.930 1804.740 ;
        RECT 2.800 1801.340 2917.930 1803.340 ;
        RECT 1.230 1786.340 2917.930 1801.340 ;
        RECT 1.230 1784.340 2917.200 1786.340 ;
        RECT 1.230 1782.940 2917.930 1784.340 ;
        RECT 2.800 1780.940 2917.930 1782.940 ;
        RECT 1.230 1769.340 2917.930 1780.940 ;
        RECT 1.230 1767.340 2917.200 1769.340 ;
        RECT 1.230 1762.540 2917.930 1767.340 ;
        RECT 2.800 1760.540 2917.930 1762.540 ;
        RECT 1.230 1748.940 2917.930 1760.540 ;
        RECT 1.230 1746.940 2917.200 1748.940 ;
        RECT 1.230 1745.540 2917.930 1746.940 ;
        RECT 2.800 1743.540 2917.930 1745.540 ;
        RECT 1.230 1728.540 2917.930 1743.540 ;
        RECT 1.230 1726.540 2917.200 1728.540 ;
        RECT 1.230 1725.140 2917.930 1726.540 ;
        RECT 2.800 1723.140 2917.930 1725.140 ;
        RECT 1.230 1708.140 2917.930 1723.140 ;
        RECT 1.230 1706.140 2917.200 1708.140 ;
        RECT 1.230 1704.740 2917.930 1706.140 ;
        RECT 2.800 1702.740 2917.930 1704.740 ;
        RECT 1.230 1687.740 2917.930 1702.740 ;
        RECT 1.230 1685.740 2917.200 1687.740 ;
        RECT 1.230 1684.340 2917.930 1685.740 ;
        RECT 2.800 1682.340 2917.930 1684.340 ;
        RECT 1.230 1667.340 2917.930 1682.340 ;
        RECT 1.230 1665.340 2917.200 1667.340 ;
        RECT 1.230 1663.940 2917.930 1665.340 ;
        RECT 2.800 1661.940 2917.930 1663.940 ;
        RECT 1.230 1646.940 2917.930 1661.940 ;
        RECT 1.230 1644.940 2917.200 1646.940 ;
        RECT 1.230 1643.540 2917.930 1644.940 ;
        RECT 2.800 1641.540 2917.930 1643.540 ;
        RECT 1.230 1626.540 2917.930 1641.540 ;
        RECT 1.230 1624.540 2917.200 1626.540 ;
        RECT 1.230 1623.140 2917.930 1624.540 ;
        RECT 2.800 1621.140 2917.930 1623.140 ;
        RECT 1.230 1606.140 2917.930 1621.140 ;
        RECT 1.230 1604.140 2917.200 1606.140 ;
        RECT 1.230 1602.740 2917.930 1604.140 ;
        RECT 2.800 1600.740 2917.930 1602.740 ;
        RECT 1.230 1585.740 2917.930 1600.740 ;
        RECT 1.230 1583.740 2917.200 1585.740 ;
        RECT 1.230 1582.340 2917.930 1583.740 ;
        RECT 2.800 1580.340 2917.930 1582.340 ;
        RECT 1.230 1568.740 2917.930 1580.340 ;
        RECT 1.230 1566.740 2917.200 1568.740 ;
        RECT 1.230 1561.940 2917.930 1566.740 ;
        RECT 2.800 1559.940 2917.930 1561.940 ;
        RECT 1.230 1548.340 2917.930 1559.940 ;
        RECT 1.230 1546.340 2917.200 1548.340 ;
        RECT 1.230 1544.940 2917.930 1546.340 ;
        RECT 2.800 1542.940 2917.930 1544.940 ;
        RECT 1.230 1527.940 2917.930 1542.940 ;
        RECT 1.230 1525.940 2917.200 1527.940 ;
        RECT 1.230 1524.540 2917.930 1525.940 ;
        RECT 2.800 1522.540 2917.930 1524.540 ;
        RECT 1.230 1507.540 2917.930 1522.540 ;
        RECT 1.230 1505.540 2917.200 1507.540 ;
        RECT 1.230 1504.140 2917.930 1505.540 ;
        RECT 2.800 1502.140 2917.930 1504.140 ;
        RECT 1.230 1487.140 2917.930 1502.140 ;
        RECT 1.230 1485.140 2917.200 1487.140 ;
        RECT 1.230 1483.740 2917.930 1485.140 ;
        RECT 2.800 1481.740 2917.930 1483.740 ;
        RECT 1.230 1466.740 2917.930 1481.740 ;
        RECT 1.230 1464.740 2917.200 1466.740 ;
        RECT 1.230 1463.340 2917.930 1464.740 ;
        RECT 2.800 1461.340 2917.930 1463.340 ;
        RECT 1.230 1446.340 2917.930 1461.340 ;
        RECT 1.230 1444.340 2917.200 1446.340 ;
        RECT 1.230 1442.940 2917.930 1444.340 ;
        RECT 2.800 1440.940 2917.930 1442.940 ;
        RECT 1.230 1425.940 2917.930 1440.940 ;
        RECT 1.230 1423.940 2917.200 1425.940 ;
        RECT 1.230 1422.540 2917.930 1423.940 ;
        RECT 2.800 1420.540 2917.930 1422.540 ;
        RECT 1.230 1405.540 2917.930 1420.540 ;
        RECT 1.230 1403.540 2917.200 1405.540 ;
        RECT 1.230 1402.140 2917.930 1403.540 ;
        RECT 2.800 1400.140 2917.930 1402.140 ;
        RECT 1.230 1385.140 2917.930 1400.140 ;
        RECT 1.230 1383.140 2917.200 1385.140 ;
        RECT 1.230 1381.740 2917.930 1383.140 ;
        RECT 2.800 1379.740 2917.930 1381.740 ;
        RECT 1.230 1368.140 2917.930 1379.740 ;
        RECT 1.230 1366.140 2917.200 1368.140 ;
        RECT 1.230 1361.340 2917.930 1366.140 ;
        RECT 2.800 1359.340 2917.930 1361.340 ;
        RECT 1.230 1347.740 2917.930 1359.340 ;
        RECT 1.230 1345.740 2917.200 1347.740 ;
        RECT 1.230 1344.340 2917.930 1345.740 ;
        RECT 2.800 1342.340 2917.930 1344.340 ;
        RECT 1.230 1327.340 2917.930 1342.340 ;
        RECT 1.230 1325.340 2917.200 1327.340 ;
        RECT 1.230 1323.940 2917.930 1325.340 ;
        RECT 2.800 1321.940 2917.930 1323.940 ;
        RECT 1.230 1306.940 2917.930 1321.940 ;
        RECT 1.230 1304.940 2917.200 1306.940 ;
        RECT 1.230 1303.540 2917.930 1304.940 ;
        RECT 2.800 1301.540 2917.930 1303.540 ;
        RECT 1.230 1286.540 2917.930 1301.540 ;
        RECT 1.230 1284.540 2917.200 1286.540 ;
        RECT 1.230 1283.140 2917.930 1284.540 ;
        RECT 2.800 1281.140 2917.930 1283.140 ;
        RECT 1.230 1266.140 2917.930 1281.140 ;
        RECT 1.230 1264.140 2917.200 1266.140 ;
        RECT 1.230 1262.740 2917.930 1264.140 ;
        RECT 2.800 1260.740 2917.930 1262.740 ;
        RECT 1.230 1245.740 2917.930 1260.740 ;
        RECT 1.230 1243.740 2917.200 1245.740 ;
        RECT 1.230 1242.340 2917.930 1243.740 ;
        RECT 2.800 1240.340 2917.930 1242.340 ;
        RECT 1.230 1225.340 2917.930 1240.340 ;
        RECT 1.230 1223.340 2917.200 1225.340 ;
        RECT 1.230 1221.940 2917.930 1223.340 ;
        RECT 2.800 1219.940 2917.930 1221.940 ;
        RECT 1.230 1204.940 2917.930 1219.940 ;
        RECT 1.230 1202.940 2917.200 1204.940 ;
        RECT 1.230 1201.540 2917.930 1202.940 ;
        RECT 2.800 1199.540 2917.930 1201.540 ;
        RECT 1.230 1187.940 2917.930 1199.540 ;
        RECT 1.230 1185.940 2917.200 1187.940 ;
        RECT 1.230 1181.140 2917.930 1185.940 ;
        RECT 2.800 1179.140 2917.930 1181.140 ;
        RECT 1.230 1167.540 2917.930 1179.140 ;
        RECT 1.230 1165.540 2917.200 1167.540 ;
        RECT 1.230 1164.140 2917.930 1165.540 ;
        RECT 2.800 1162.140 2917.930 1164.140 ;
        RECT 1.230 1147.140 2917.930 1162.140 ;
        RECT 1.230 1145.140 2917.200 1147.140 ;
        RECT 1.230 1143.740 2917.930 1145.140 ;
        RECT 2.800 1141.740 2917.930 1143.740 ;
        RECT 1.230 1126.740 2917.930 1141.740 ;
        RECT 1.230 1124.740 2917.200 1126.740 ;
        RECT 1.230 1123.340 2917.930 1124.740 ;
        RECT 2.800 1121.340 2917.930 1123.340 ;
        RECT 1.230 1106.340 2917.930 1121.340 ;
        RECT 1.230 1104.340 2917.200 1106.340 ;
        RECT 1.230 1102.940 2917.930 1104.340 ;
        RECT 2.800 1100.940 2917.930 1102.940 ;
        RECT 1.230 1085.940 2917.930 1100.940 ;
        RECT 1.230 1083.940 2917.200 1085.940 ;
        RECT 1.230 1082.540 2917.930 1083.940 ;
        RECT 2.800 1080.540 2917.930 1082.540 ;
        RECT 1.230 1065.540 2917.930 1080.540 ;
        RECT 1.230 1063.540 2917.200 1065.540 ;
        RECT 1.230 1062.140 2917.930 1063.540 ;
        RECT 2.800 1060.140 2917.930 1062.140 ;
        RECT 1.230 1045.140 2917.930 1060.140 ;
        RECT 1.230 1043.140 2917.200 1045.140 ;
        RECT 1.230 1041.740 2917.930 1043.140 ;
        RECT 2.800 1039.740 2917.930 1041.740 ;
        RECT 1.230 1024.740 2917.930 1039.740 ;
        RECT 1.230 1022.740 2917.200 1024.740 ;
        RECT 1.230 1021.340 2917.930 1022.740 ;
        RECT 2.800 1019.340 2917.930 1021.340 ;
        RECT 1.230 1004.340 2917.930 1019.340 ;
        RECT 1.230 1002.340 2917.200 1004.340 ;
        RECT 1.230 1000.940 2917.930 1002.340 ;
        RECT 2.800 998.940 2917.930 1000.940 ;
        RECT 1.230 987.340 2917.930 998.940 ;
        RECT 1.230 985.340 2917.200 987.340 ;
        RECT 1.230 980.540 2917.930 985.340 ;
        RECT 2.800 978.540 2917.930 980.540 ;
        RECT 1.230 966.940 2917.930 978.540 ;
        RECT 1.230 964.940 2917.200 966.940 ;
        RECT 1.230 963.540 2917.930 964.940 ;
        RECT 2.800 961.540 2917.930 963.540 ;
        RECT 1.230 946.540 2917.930 961.540 ;
        RECT 1.230 944.540 2917.200 946.540 ;
        RECT 1.230 943.140 2917.930 944.540 ;
        RECT 2.800 941.140 2917.930 943.140 ;
        RECT 1.230 926.140 2917.930 941.140 ;
        RECT 1.230 924.140 2917.200 926.140 ;
        RECT 1.230 922.740 2917.930 924.140 ;
        RECT 2.800 920.740 2917.930 922.740 ;
        RECT 1.230 905.740 2917.930 920.740 ;
        RECT 1.230 903.740 2917.200 905.740 ;
        RECT 1.230 902.340 2917.930 903.740 ;
        RECT 2.800 900.340 2917.930 902.340 ;
        RECT 1.230 885.340 2917.930 900.340 ;
        RECT 1.230 883.340 2917.200 885.340 ;
        RECT 1.230 881.940 2917.930 883.340 ;
        RECT 2.800 879.940 2917.930 881.940 ;
        RECT 1.230 864.940 2917.930 879.940 ;
        RECT 1.230 862.940 2917.200 864.940 ;
        RECT 1.230 861.540 2917.930 862.940 ;
        RECT 2.800 859.540 2917.930 861.540 ;
        RECT 1.230 844.540 2917.930 859.540 ;
        RECT 1.230 842.540 2917.200 844.540 ;
        RECT 1.230 841.140 2917.930 842.540 ;
        RECT 2.800 839.140 2917.930 841.140 ;
        RECT 1.230 824.140 2917.930 839.140 ;
        RECT 1.230 822.140 2917.200 824.140 ;
        RECT 1.230 820.740 2917.930 822.140 ;
        RECT 2.800 818.740 2917.930 820.740 ;
        RECT 1.230 803.740 2917.930 818.740 ;
        RECT 1.230 801.740 2917.200 803.740 ;
        RECT 1.230 800.340 2917.930 801.740 ;
        RECT 2.800 798.340 2917.930 800.340 ;
        RECT 1.230 786.740 2917.930 798.340 ;
        RECT 1.230 784.740 2917.200 786.740 ;
        RECT 1.230 779.940 2917.930 784.740 ;
        RECT 2.800 777.940 2917.930 779.940 ;
        RECT 1.230 766.340 2917.930 777.940 ;
        RECT 1.230 764.340 2917.200 766.340 ;
        RECT 1.230 762.940 2917.930 764.340 ;
        RECT 2.800 760.940 2917.930 762.940 ;
        RECT 1.230 745.940 2917.930 760.940 ;
        RECT 1.230 743.940 2917.200 745.940 ;
        RECT 1.230 742.540 2917.930 743.940 ;
        RECT 2.800 740.540 2917.930 742.540 ;
        RECT 1.230 725.540 2917.930 740.540 ;
        RECT 1.230 723.540 2917.200 725.540 ;
        RECT 1.230 722.140 2917.930 723.540 ;
        RECT 2.800 720.140 2917.930 722.140 ;
        RECT 1.230 705.140 2917.930 720.140 ;
        RECT 1.230 703.140 2917.200 705.140 ;
        RECT 1.230 701.740 2917.930 703.140 ;
        RECT 2.800 699.740 2917.930 701.740 ;
        RECT 1.230 684.740 2917.930 699.740 ;
        RECT 1.230 682.740 2917.200 684.740 ;
        RECT 1.230 681.340 2917.930 682.740 ;
        RECT 2.800 679.340 2917.930 681.340 ;
        RECT 1.230 664.340 2917.930 679.340 ;
        RECT 1.230 662.340 2917.200 664.340 ;
        RECT 1.230 660.940 2917.930 662.340 ;
        RECT 2.800 658.940 2917.930 660.940 ;
        RECT 1.230 643.940 2917.930 658.940 ;
        RECT 1.230 641.940 2917.200 643.940 ;
        RECT 1.230 640.540 2917.930 641.940 ;
        RECT 2.800 638.540 2917.930 640.540 ;
        RECT 1.230 623.540 2917.930 638.540 ;
        RECT 1.230 621.540 2917.200 623.540 ;
        RECT 1.230 620.140 2917.930 621.540 ;
        RECT 2.800 618.140 2917.930 620.140 ;
        RECT 1.230 606.540 2917.930 618.140 ;
        RECT 1.230 604.540 2917.200 606.540 ;
        RECT 1.230 599.740 2917.930 604.540 ;
        RECT 2.800 597.740 2917.930 599.740 ;
        RECT 1.230 586.140 2917.930 597.740 ;
        RECT 1.230 584.140 2917.200 586.140 ;
        RECT 1.230 582.740 2917.930 584.140 ;
        RECT 2.800 580.740 2917.930 582.740 ;
        RECT 1.230 565.740 2917.930 580.740 ;
        RECT 1.230 563.740 2917.200 565.740 ;
        RECT 1.230 562.340 2917.930 563.740 ;
        RECT 2.800 560.340 2917.930 562.340 ;
        RECT 1.230 545.340 2917.930 560.340 ;
        RECT 1.230 543.340 2917.200 545.340 ;
        RECT 1.230 541.940 2917.930 543.340 ;
        RECT 2.800 539.940 2917.930 541.940 ;
        RECT 1.230 524.940 2917.930 539.940 ;
        RECT 1.230 522.940 2917.200 524.940 ;
        RECT 1.230 521.540 2917.930 522.940 ;
        RECT 2.800 519.540 2917.930 521.540 ;
        RECT 1.230 504.540 2917.930 519.540 ;
        RECT 1.230 502.540 2917.200 504.540 ;
        RECT 1.230 501.140 2917.930 502.540 ;
        RECT 2.800 499.140 2917.930 501.140 ;
        RECT 1.230 484.140 2917.930 499.140 ;
        RECT 1.230 482.140 2917.200 484.140 ;
        RECT 1.230 480.740 2917.930 482.140 ;
        RECT 2.800 478.740 2917.930 480.740 ;
        RECT 1.230 463.740 2917.930 478.740 ;
        RECT 1.230 461.740 2917.200 463.740 ;
        RECT 1.230 460.340 2917.930 461.740 ;
        RECT 2.800 458.340 2917.930 460.340 ;
        RECT 1.230 443.340 2917.930 458.340 ;
        RECT 1.230 441.340 2917.200 443.340 ;
        RECT 1.230 439.940 2917.930 441.340 ;
        RECT 2.800 437.940 2917.930 439.940 ;
        RECT 1.230 422.940 2917.930 437.940 ;
        RECT 1.230 420.940 2917.200 422.940 ;
        RECT 1.230 419.540 2917.930 420.940 ;
        RECT 2.800 417.540 2917.930 419.540 ;
        RECT 1.230 405.940 2917.930 417.540 ;
        RECT 1.230 403.940 2917.200 405.940 ;
        RECT 1.230 399.140 2917.930 403.940 ;
        RECT 2.800 397.140 2917.930 399.140 ;
        RECT 1.230 385.540 2917.930 397.140 ;
        RECT 1.230 383.540 2917.200 385.540 ;
        RECT 1.230 382.140 2917.930 383.540 ;
        RECT 2.800 380.140 2917.930 382.140 ;
        RECT 1.230 365.140 2917.930 380.140 ;
        RECT 1.230 363.140 2917.200 365.140 ;
        RECT 1.230 361.740 2917.930 363.140 ;
        RECT 2.800 359.740 2917.930 361.740 ;
        RECT 1.230 344.740 2917.930 359.740 ;
        RECT 1.230 342.740 2917.200 344.740 ;
        RECT 1.230 341.340 2917.930 342.740 ;
        RECT 2.800 339.340 2917.930 341.340 ;
        RECT 1.230 324.340 2917.930 339.340 ;
        RECT 1.230 322.340 2917.200 324.340 ;
        RECT 1.230 320.940 2917.930 322.340 ;
        RECT 2.800 318.940 2917.930 320.940 ;
        RECT 1.230 303.940 2917.930 318.940 ;
        RECT 1.230 301.940 2917.200 303.940 ;
        RECT 1.230 300.540 2917.930 301.940 ;
        RECT 2.800 298.540 2917.930 300.540 ;
        RECT 1.230 283.540 2917.930 298.540 ;
        RECT 1.230 281.540 2917.200 283.540 ;
        RECT 1.230 280.140 2917.930 281.540 ;
        RECT 2.800 278.140 2917.930 280.140 ;
        RECT 1.230 263.140 2917.930 278.140 ;
        RECT 1.230 261.140 2917.200 263.140 ;
        RECT 1.230 259.740 2917.930 261.140 ;
        RECT 2.800 257.740 2917.930 259.740 ;
        RECT 1.230 242.740 2917.930 257.740 ;
        RECT 1.230 240.740 2917.200 242.740 ;
        RECT 1.230 239.340 2917.930 240.740 ;
        RECT 2.800 237.340 2917.930 239.340 ;
        RECT 1.230 222.340 2917.930 237.340 ;
        RECT 1.230 220.340 2917.200 222.340 ;
        RECT 1.230 218.940 2917.930 220.340 ;
        RECT 2.800 216.940 2917.930 218.940 ;
        RECT 1.230 205.340 2917.930 216.940 ;
        RECT 1.230 203.340 2917.200 205.340 ;
        RECT 1.230 198.540 2917.930 203.340 ;
        RECT 2.800 196.540 2917.930 198.540 ;
        RECT 1.230 184.940 2917.930 196.540 ;
        RECT 1.230 182.940 2917.200 184.940 ;
        RECT 1.230 181.540 2917.930 182.940 ;
        RECT 2.800 179.540 2917.930 181.540 ;
        RECT 1.230 164.540 2917.930 179.540 ;
        RECT 1.230 162.540 2917.200 164.540 ;
        RECT 1.230 161.140 2917.930 162.540 ;
        RECT 2.800 159.140 2917.930 161.140 ;
        RECT 1.230 144.140 2917.930 159.140 ;
        RECT 1.230 142.140 2917.200 144.140 ;
        RECT 1.230 140.740 2917.930 142.140 ;
        RECT 2.800 138.740 2917.930 140.740 ;
        RECT 1.230 123.740 2917.930 138.740 ;
        RECT 1.230 121.740 2917.200 123.740 ;
        RECT 1.230 120.340 2917.930 121.740 ;
        RECT 2.800 118.340 2917.930 120.340 ;
        RECT 1.230 103.340 2917.930 118.340 ;
        RECT 1.230 101.340 2917.200 103.340 ;
        RECT 1.230 99.940 2917.930 101.340 ;
        RECT 2.800 97.940 2917.930 99.940 ;
        RECT 1.230 82.940 2917.930 97.940 ;
        RECT 1.230 80.940 2917.200 82.940 ;
        RECT 1.230 79.540 2917.930 80.940 ;
        RECT 2.800 77.540 2917.930 79.540 ;
        RECT 1.230 62.540 2917.930 77.540 ;
        RECT 1.230 60.540 2917.200 62.540 ;
        RECT 1.230 59.140 2917.930 60.540 ;
        RECT 2.800 57.140 2917.930 59.140 ;
        RECT 1.230 42.140 2917.930 57.140 ;
        RECT 1.230 40.140 2917.200 42.140 ;
        RECT 1.230 38.740 2917.930 40.140 ;
        RECT 2.800 36.740 2917.930 38.740 ;
        RECT 1.230 25.140 2917.930 36.740 ;
        RECT 1.230 23.140 2917.200 25.140 ;
        RECT 1.230 18.340 2917.930 23.140 ;
        RECT 2.800 16.340 2917.930 18.340 ;
        RECT 1.230 4.740 2917.930 16.340 ;
        RECT 1.230 3.575 2917.200 4.740 ;
      LAYER met4 ;
        RECT 478.695 172.215 481.070 3284.905 ;
        RECT 484.970 172.215 503.570 3284.905 ;
        RECT 507.470 172.215 526.070 3284.905 ;
        RECT 529.970 172.215 548.570 3284.905 ;
        RECT 552.470 172.215 571.070 3284.905 ;
        RECT 574.970 1309.600 593.570 3284.905 ;
        RECT 597.470 1309.600 616.070 3284.905 ;
        RECT 619.970 1309.600 638.570 3284.905 ;
        RECT 642.470 1309.600 661.070 3284.905 ;
        RECT 664.970 1309.600 683.570 3284.905 ;
        RECT 687.470 1309.600 706.070 3284.905 ;
        RECT 709.970 1309.600 728.570 3284.905 ;
        RECT 732.470 1309.600 751.070 3284.905 ;
        RECT 754.970 1309.600 773.570 3284.905 ;
        RECT 777.470 1309.600 796.070 3284.905 ;
        RECT 799.970 1309.600 818.570 3284.905 ;
        RECT 822.470 1309.600 841.070 3284.905 ;
        RECT 844.970 1309.600 863.570 3284.905 ;
        RECT 867.470 1309.600 886.070 3284.905 ;
        RECT 889.970 1309.600 908.570 3284.905 ;
        RECT 912.470 1309.600 931.070 3284.905 ;
        RECT 934.970 1309.600 953.570 3284.905 ;
        RECT 957.470 1309.600 976.070 3284.905 ;
        RECT 574.970 990.400 976.070 1309.600 ;
        RECT 574.970 709.600 593.570 990.400 ;
        RECT 597.470 709.600 616.070 990.400 ;
        RECT 619.970 709.600 706.070 990.400 ;
        RECT 709.970 709.600 728.570 990.400 ;
        RECT 732.470 709.600 751.070 990.400 ;
        RECT 754.970 709.600 773.570 990.400 ;
        RECT 777.470 709.600 796.070 990.400 ;
        RECT 799.970 709.600 886.070 990.400 ;
        RECT 889.970 709.600 908.570 990.400 ;
        RECT 912.470 709.600 931.070 990.400 ;
        RECT 934.970 709.600 953.570 990.400 ;
        RECT 957.470 709.600 976.070 990.400 ;
        RECT 574.970 390.400 976.070 709.600 ;
        RECT 574.970 172.215 593.570 390.400 ;
        RECT 597.470 172.215 616.070 390.400 ;
        RECT 619.970 172.215 638.570 390.400 ;
        RECT 642.470 172.215 661.070 390.400 ;
        RECT 664.970 172.215 683.570 390.400 ;
        RECT 687.470 172.215 706.070 390.400 ;
        RECT 709.970 172.215 728.570 390.400 ;
        RECT 732.470 172.215 751.070 390.400 ;
        RECT 754.970 172.215 773.570 390.400 ;
        RECT 777.470 172.215 796.070 390.400 ;
        RECT 799.970 172.215 818.570 390.400 ;
        RECT 822.470 172.215 841.070 390.400 ;
        RECT 844.970 172.215 863.570 390.400 ;
        RECT 867.470 172.215 886.070 390.400 ;
        RECT 889.970 172.215 908.570 390.400 ;
        RECT 912.470 172.215 931.070 390.400 ;
        RECT 934.970 172.215 953.570 390.400 ;
        RECT 957.470 172.215 976.070 390.400 ;
        RECT 979.970 172.215 998.570 3284.905 ;
        RECT 1002.470 172.215 1021.070 3284.905 ;
        RECT 1024.970 172.215 1043.570 3284.905 ;
        RECT 1047.470 172.215 1055.865 3284.905 ;
  END
END user_project_wrapper
END LIBRARY

